module fake_jpeg_1123_n_691 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_691);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_691;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_612;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_19),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_19),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_61),
.B(n_62),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_18),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g156 ( 
.A(n_63),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_39),
.B(n_16),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_64),
.B(n_75),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_26),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_68),
.Y(n_207)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_70),
.B(n_84),
.Y(n_138)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_73),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_74),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_48),
.B(n_57),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_76),
.Y(n_200)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_77),
.Y(n_193)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_78),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_35),
.B(n_16),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_79),
.B(n_94),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_80),
.Y(n_194)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_81),
.Y(n_204)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_82),
.Y(n_175)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_83),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_14),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_86),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_87),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_88),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_89),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_90),
.Y(n_201)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_92),
.Y(n_206)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_93),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_21),
.B(n_15),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_59),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_109),
.Y(n_145)
);

CKINVDCx9p33_ASAP7_75t_R g96 ( 
.A(n_55),
.Y(n_96)
);

INVx13_ASAP7_75t_L g220 ( 
.A(n_96),
.Y(n_220)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_98),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_21),
.B(n_15),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_99),
.B(n_127),
.Y(n_195)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_100),
.Y(n_181)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_102),
.Y(n_215)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_103),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_104),
.Y(n_172)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_43),
.Y(n_105)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_105),
.Y(n_187)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_106),
.Y(n_223)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_22),
.Y(n_107)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_108),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_59),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_33),
.Y(n_111)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_28),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_112),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_34),
.Y(n_113)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_33),
.Y(n_114)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

INVx4_ASAP7_75t_SL g115 ( 
.A(n_34),
.Y(n_115)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_33),
.Y(n_116)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_116),
.Y(n_213)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_117),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_27),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_124),
.Y(n_161)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_36),
.Y(n_119)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_40),
.Y(n_120)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_123),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_27),
.B(n_53),
.Y(n_124)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_125),
.Y(n_189)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_40),
.Y(n_126)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_38),
.B(n_11),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_32),
.Y(n_128)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_128),
.Y(n_216)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_28),
.Y(n_129)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_129),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_30),
.Y(n_130)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_32),
.Y(n_131)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_51),
.Y(n_132)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_132),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_131),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_134),
.Y(n_291)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_136),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_112),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_137),
.B(n_139),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_114),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_88),
.A2(n_41),
.B1(n_29),
.B2(n_25),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_143),
.A2(n_166),
.B1(n_23),
.B2(n_31),
.Y(n_248)
);

NAND3xp33_ASAP7_75t_SL g147 ( 
.A(n_84),
.B(n_57),
.C(n_32),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_147),
.B(n_192),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_94),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_154),
.B(n_162),
.Y(n_239)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_158),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_79),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_90),
.A2(n_29),
.B1(n_41),
.B2(n_25),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_68),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_168),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_44),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_170),
.B(n_179),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_122),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_178),
.B(n_203),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_130),
.B(n_44),
.Y(n_179)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_76),
.Y(n_183)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_183),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_65),
.A2(n_58),
.B1(n_54),
.B2(n_37),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_188),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_125),
.B(n_86),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_115),
.A2(n_25),
.B1(n_41),
.B2(n_29),
.Y(n_197)
);

OA22x2_ASAP7_75t_L g280 ( 
.A1(n_197),
.A2(n_8),
.B1(n_9),
.B2(n_166),
.Y(n_280)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_130),
.B(n_38),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_202),
.B(n_209),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_83),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_116),
.Y(n_205)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_67),
.B(n_53),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_72),
.B(n_56),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_211),
.B(n_218),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_81),
.B(n_58),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_91),
.Y(n_219)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_107),
.Y(n_221)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_108),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_230),
.Y(n_249)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_74),
.Y(n_225)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_87),
.B(n_56),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_227),
.B(n_142),
.Y(n_314)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_92),
.Y(n_229)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_229),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_102),
.B(n_54),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_192),
.A2(n_23),
.B1(n_37),
.B2(n_31),
.Y(n_231)
);

A2O1A1Ixp33_ASAP7_75t_SL g365 ( 
.A1(n_231),
.A2(n_258),
.B(n_276),
.C(n_280),
.Y(n_365)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_133),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_233),
.Y(n_355)
);

BUFx12_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_234),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_168),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_236),
.B(n_238),
.Y(n_318)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_133),
.Y(n_237)
);

INVx5_ASAP7_75t_L g349 ( 
.A(n_237),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_145),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g240 ( 
.A(n_163),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_240),
.Y(n_319)
);

BUFx12f_ASAP7_75t_L g241 ( 
.A(n_163),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_241),
.Y(n_347)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_152),
.Y(n_247)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_247),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_248),
.A2(n_263),
.B1(n_272),
.B2(n_215),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_177),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_250),
.B(n_266),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_144),
.Y(n_252)
);

INVx8_ASAP7_75t_L g376 ( 
.A(n_252),
.Y(n_376)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_207),
.Y(n_254)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_254),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_214),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_255),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_161),
.B(n_30),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_256),
.B(n_259),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_182),
.A2(n_23),
.B1(n_106),
.B2(n_3),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_217),
.B(n_1),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_262),
.A2(n_136),
.B1(n_215),
.B2(n_206),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_159),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_167),
.B(n_11),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_264),
.B(n_270),
.Y(n_322)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_144),
.Y(n_265)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_265),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_220),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_140),
.Y(n_267)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_267),
.Y(n_321)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_160),
.Y(n_268)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_268),
.Y(n_372)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_151),
.Y(n_269)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_269),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_177),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_138),
.B(n_2),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_271),
.B(n_275),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_143),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_195),
.B(n_10),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_273),
.B(n_278),
.Y(n_333)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_181),
.Y(n_274)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_274),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_149),
.B(n_4),
.Y(n_275)
);

AO22x2_ASAP7_75t_L g276 ( 
.A1(n_190),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_187),
.Y(n_277)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_277),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_227),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_180),
.Y(n_279)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_279),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_182),
.A2(n_8),
.B1(n_9),
.B2(n_173),
.Y(n_281)
);

OA22x2_ASAP7_75t_L g342 ( 
.A1(n_281),
.A2(n_284),
.B1(n_165),
.B2(n_157),
.Y(n_342)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_176),
.Y(n_282)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_282),
.Y(n_343)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_200),
.Y(n_283)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_283),
.Y(n_377)
);

OA22x2_ASAP7_75t_L g284 ( 
.A1(n_197),
.A2(n_9),
.B1(n_155),
.B2(n_191),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_198),
.B(n_9),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_285),
.B(n_298),
.Y(n_366)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_153),
.Y(n_286)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_286),
.Y(n_348)
);

CKINVDCx12_ASAP7_75t_R g287 ( 
.A(n_220),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_287),
.B(n_290),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_193),
.Y(n_288)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_288),
.Y(n_357)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_212),
.Y(n_289)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_289),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_146),
.B(n_188),
.Y(n_290)
);

INVx8_ASAP7_75t_L g292 ( 
.A(n_189),
.Y(n_292)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_292),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_135),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_293),
.B(n_174),
.Y(n_364)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_204),
.Y(n_294)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_294),
.Y(n_361)
);

BUFx12f_ASAP7_75t_L g295 ( 
.A(n_223),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_305),
.Y(n_323)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_194),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_296),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_210),
.B(n_142),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_226),
.Y(n_299)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_299),
.Y(n_363)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_156),
.Y(n_300)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_300),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_180),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_301),
.B(n_307),
.Y(n_369)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_189),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_308),
.Y(n_324)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_194),
.Y(n_305)
);

INVx6_ASAP7_75t_L g307 ( 
.A(n_185),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_175),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_185),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_309),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_193),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_310),
.B(n_312),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_186),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_311),
.Y(n_350)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_186),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_156),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_306),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_315),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_214),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_262),
.A2(n_150),
.B1(n_171),
.B2(n_228),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_316),
.A2(n_328),
.B1(n_279),
.B2(n_311),
.Y(n_409)
);

AOI32xp33_ASAP7_75t_L g317 ( 
.A1(n_239),
.A2(n_172),
.A3(n_169),
.B1(n_147),
.B2(n_213),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_317),
.B(n_344),
.Y(n_379)
);

CKINVDCx14_ASAP7_75t_R g422 ( 
.A(n_320),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_249),
.B(n_222),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_325),
.B(n_371),
.Y(n_381)
);

AO22x2_ASAP7_75t_L g329 ( 
.A1(n_280),
.A2(n_284),
.B1(n_272),
.B2(n_257),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_329),
.B(n_337),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_196),
.C(n_208),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_330),
.B(n_303),
.C(n_242),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_257),
.A2(n_216),
.B(n_222),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_331),
.A2(n_352),
.B(n_258),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_251),
.B(n_164),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_334),
.B(n_364),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_148),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_335),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_SL g406 ( 
.A1(n_342),
.A2(n_351),
.B1(n_315),
.B2(n_241),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_297),
.B(n_194),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_260),
.A2(n_245),
.B1(n_280),
.B2(n_231),
.Y(n_351)
);

OAI21xp33_ASAP7_75t_L g352 ( 
.A1(n_253),
.A2(n_223),
.B(n_228),
.Y(n_352)
);

OA22x2_ASAP7_75t_L g360 ( 
.A1(n_284),
.A2(n_174),
.B1(n_213),
.B2(n_157),
.Y(n_360)
);

AO22x2_ASAP7_75t_L g427 ( 
.A1(n_360),
.A2(n_242),
.B1(n_234),
.B2(n_141),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_304),
.A2(n_165),
.B1(n_184),
.B2(n_201),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_368),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_255),
.A2(n_184),
.B1(n_201),
.B2(n_206),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_370),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_291),
.B(n_150),
.Y(n_371)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_324),
.Y(n_378)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_378),
.Y(n_439)
);

AND2x6_ASAP7_75t_L g380 ( 
.A(n_352),
.B(n_296),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_380),
.B(n_388),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_355),
.Y(n_382)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_382),
.Y(n_462)
);

OAI32xp33_ASAP7_75t_L g383 ( 
.A1(n_362),
.A2(n_276),
.A3(n_232),
.B1(n_235),
.B2(n_244),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_383),
.B(n_411),
.Y(n_454)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_321),
.Y(n_384)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_384),
.Y(n_440)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_348),
.Y(n_385)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_385),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_318),
.B(n_366),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_386),
.B(n_387),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_334),
.B(n_243),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_326),
.B(n_261),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_361),
.Y(n_389)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_389),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_355),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_390),
.Y(n_442)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_367),
.Y(n_391)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_391),
.Y(n_446)
);

INVx6_ASAP7_75t_L g392 ( 
.A(n_376),
.Y(n_392)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_392),
.Y(n_452)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_324),
.Y(n_394)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_394),
.Y(n_453)
);

AND2x6_ASAP7_75t_L g395 ( 
.A(n_325),
.B(n_276),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_395),
.B(n_397),
.Y(n_461)
);

INVx11_ASAP7_75t_L g396 ( 
.A(n_327),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g447 ( 
.A1(n_396),
.A2(n_407),
.B1(n_408),
.B2(n_412),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_330),
.B(n_288),
.Y(n_397)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_377),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_399),
.Y(n_437)
);

INVx6_ASAP7_75t_L g400 ( 
.A(n_376),
.Y(n_400)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_400),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_333),
.B(n_310),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_401),
.B(n_404),
.Y(n_464)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_358),
.Y(n_402)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_402),
.Y(n_467)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_324),
.Y(n_403)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_403),
.Y(n_469)
);

BUFx4f_ASAP7_75t_SL g404 ( 
.A(n_357),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_346),
.B(n_292),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_405),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_406),
.A2(n_413),
.B(n_410),
.Y(n_445)
);

INVx13_ASAP7_75t_L g407 ( 
.A(n_339),
.Y(n_407)
);

INVx13_ASAP7_75t_L g408 ( 
.A(n_339),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_409),
.A2(n_423),
.B1(n_424),
.B2(n_350),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_371),
.B(n_312),
.Y(n_411)
);

INVx8_ASAP7_75t_L g412 ( 
.A(n_345),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_329),
.B(n_265),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_414),
.B(n_416),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g416 ( 
.A(n_331),
.B(n_241),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_417),
.B(n_332),
.C(n_359),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_329),
.B(n_233),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_419),
.B(n_398),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_322),
.B(n_246),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_420),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_337),
.A2(n_171),
.B1(n_281),
.B2(n_307),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_421),
.A2(n_415),
.B1(n_393),
.B2(n_409),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_316),
.A2(n_301),
.B1(n_252),
.B2(n_309),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_363),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_365),
.A2(n_303),
.B(n_246),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_425),
.A2(n_365),
.B(n_342),
.Y(n_430)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_354),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_426),
.B(n_427),
.Y(n_434)
);

AND2x2_ASAP7_75t_SL g428 ( 
.A(n_381),
.B(n_335),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_428),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_429),
.A2(n_433),
.B1(n_436),
.B2(n_449),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_430),
.A2(n_347),
.B(n_319),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_413),
.A2(n_365),
.B(n_374),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_431),
.A2(n_445),
.B(n_448),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_393),
.A2(n_329),
.B1(n_365),
.B2(n_360),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_381),
.B(n_335),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_435),
.B(n_450),
.C(n_451),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_393),
.A2(n_414),
.B1(n_419),
.B2(n_421),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_425),
.A2(n_360),
.B1(n_342),
.B2(n_368),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_438),
.A2(n_430),
.B1(n_433),
.B2(n_431),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_444),
.A2(n_349),
.B1(n_372),
.B2(n_341),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_418),
.A2(n_332),
.B(n_320),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_422),
.A2(n_370),
.B1(n_360),
.B2(n_369),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_332),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_379),
.A2(n_342),
.B(n_338),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_457),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_415),
.A2(n_375),
.B1(n_349),
.B2(n_373),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_458),
.A2(n_396),
.B1(n_399),
.B2(n_373),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_398),
.B(n_411),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_460),
.B(n_372),
.C(n_354),
.Y(n_503)
);

NOR2x1_ASAP7_75t_L g488 ( 
.A(n_463),
.B(n_465),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_383),
.A2(n_323),
.B(n_319),
.Y(n_465)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_443),
.Y(n_470)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_470),
.Y(n_518)
);

AOI22x1_ASAP7_75t_SL g471 ( 
.A1(n_454),
.A2(n_380),
.B1(n_416),
.B2(n_395),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_471),
.A2(n_472),
.B1(n_479),
.B2(n_493),
.Y(n_541)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_462),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_474),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_432),
.B(n_426),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_475),
.B(n_478),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_466),
.B(n_378),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_476),
.B(n_480),
.Y(n_510)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_443),
.Y(n_477)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_477),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_432),
.B(n_353),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_436),
.A2(n_410),
.B1(n_423),
.B2(n_403),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_466),
.B(n_353),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_437),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_481),
.B(n_486),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_454),
.A2(n_394),
.B1(n_427),
.B2(n_412),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_482),
.A2(n_487),
.B1(n_497),
.B2(n_434),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_459),
.B(n_377),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_483),
.B(n_499),
.Y(n_513)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_440),
.Y(n_484)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_484),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_437),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_468),
.A2(n_427),
.B1(n_400),
.B2(n_392),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_439),
.B(n_404),
.Y(n_489)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_489),
.Y(n_528)
);

INVx13_ASAP7_75t_L g490 ( 
.A(n_447),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_490),
.Y(n_524)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_440),
.Y(n_491)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_491),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_439),
.B(n_404),
.Y(n_492)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_492),
.Y(n_540)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_441),
.Y(n_494)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_494),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_462),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_495),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_434),
.A2(n_427),
.B1(n_390),
.B2(n_382),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_453),
.B(n_375),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_498),
.B(n_507),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g499 ( 
.A(n_464),
.Y(n_499)
);

OAI21xp33_ASAP7_75t_L g500 ( 
.A1(n_448),
.A2(n_340),
.B(n_336),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_500),
.B(n_502),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_459),
.B(n_455),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_503),
.B(n_506),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_505),
.A2(n_445),
.B(n_465),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_451),
.B(n_343),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_460),
.B(n_347),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_508),
.B(n_450),
.C(n_463),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_476),
.B(n_461),
.Y(n_509)
);

CKINVDCx16_ASAP7_75t_R g551 ( 
.A(n_509),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_514),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_515),
.B(n_543),
.Y(n_562)
);

NOR2x1_ASAP7_75t_L g521 ( 
.A(n_488),
.B(n_435),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_521),
.B(n_539),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_481),
.B(n_469),
.Y(n_522)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_522),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_486),
.B(n_469),
.Y(n_523)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_523),
.Y(n_560)
);

XNOR2x1_ASAP7_75t_L g526 ( 
.A(n_508),
.B(n_468),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_SL g559 ( 
.A(n_526),
.B(n_531),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_473),
.B(n_446),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_529),
.B(n_532),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_504),
.A2(n_434),
.B1(n_438),
.B2(n_457),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_530),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_SL g531 ( 
.A(n_473),
.B(n_428),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_504),
.B(n_446),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_488),
.B(n_441),
.Y(n_534)
);

CKINVDCx16_ASAP7_75t_R g553 ( 
.A(n_534),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_536),
.A2(n_472),
.B1(n_497),
.B2(n_479),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_506),
.B(n_428),
.C(n_453),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_537),
.B(n_496),
.C(n_498),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_503),
.B(n_467),
.Y(n_538)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_538),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_470),
.B(n_467),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_501),
.B(n_429),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_501),
.B(n_434),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_544),
.B(n_523),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_477),
.B(n_456),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_545),
.B(n_452),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_489),
.B(n_456),
.Y(n_546)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_546),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_522),
.B(n_492),
.Y(n_547)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_547),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_549),
.A2(n_519),
.B1(n_524),
.B2(n_525),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_550),
.B(n_537),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_531),
.B(n_496),
.C(n_485),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_552),
.B(n_571),
.C(n_578),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_514),
.A2(n_505),
.B(n_482),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_561),
.Y(n_589)
);

MAJx2_ASAP7_75t_L g584 ( 
.A(n_563),
.B(n_565),
.C(n_573),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_510),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_564),
.B(n_568),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_SL g565 ( 
.A(n_515),
.B(n_471),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_536),
.A2(n_487),
.B1(n_494),
.B2(n_491),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_566),
.A2(n_569),
.B1(n_528),
.B2(n_544),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_518),
.Y(n_567)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_567),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_512),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_530),
.A2(n_484),
.B1(n_490),
.B2(n_452),
.Y(n_569)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_570),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_517),
.B(n_442),
.C(n_474),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_511),
.B(n_341),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_572),
.B(n_577),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_517),
.B(n_407),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_546),
.B(n_495),
.Y(n_574)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_574),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_512),
.B(n_495),
.Y(n_576)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_576),
.Y(n_605)
);

FAx1_ASAP7_75t_SL g577 ( 
.A(n_521),
.B(n_408),
.CI(n_240),
.CON(n_577),
.SN(n_577)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_526),
.B(n_356),
.C(n_240),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_528),
.B(n_237),
.Y(n_579)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_579),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_581),
.B(n_585),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_562),
.B(n_573),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_582),
.B(n_578),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_550),
.B(n_543),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g586 ( 
.A1(n_553),
.A2(n_527),
.B1(n_524),
.B2(n_540),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_586),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_551),
.B(n_513),
.Y(n_590)
);

CKINVDCx14_ASAP7_75t_R g610 ( 
.A(n_590),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_571),
.B(n_541),
.C(n_540),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_591),
.B(n_595),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_SL g614 ( 
.A1(n_593),
.A2(n_600),
.B1(n_561),
.B2(n_560),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_562),
.B(n_516),
.C(n_542),
.Y(n_595)
);

BUFx24_ASAP7_75t_SL g596 ( 
.A(n_557),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_SL g616 ( 
.A(n_596),
.B(n_601),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_552),
.B(n_519),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_599),
.B(n_569),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_558),
.B(n_542),
.Y(n_601)
);

XOR2x1_ASAP7_75t_SL g602 ( 
.A(n_577),
.B(n_520),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_SL g617 ( 
.A1(n_602),
.A2(n_555),
.B(n_575),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_549),
.A2(n_520),
.B1(n_525),
.B2(n_535),
.Y(n_603)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_603),
.Y(n_620)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_547),
.Y(n_604)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_604),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_608),
.B(n_613),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_SL g611 ( 
.A1(n_598),
.A2(n_556),
.B(n_548),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_611),
.B(n_625),
.Y(n_634)
);

XOR2xp5_ASAP7_75t_L g640 ( 
.A(n_612),
.B(n_584),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_595),
.B(n_565),
.C(n_563),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_614),
.Y(n_635)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_617),
.Y(n_628)
);

BUFx12_ASAP7_75t_L g618 ( 
.A(n_591),
.Y(n_618)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_618),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_587),
.B(n_574),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_619),
.B(n_621),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_594),
.B(n_576),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_588),
.B(n_567),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_622),
.B(n_624),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_580),
.A2(n_566),
.B1(n_554),
.B2(n_560),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_623),
.A2(n_626),
.B1(n_614),
.B2(n_607),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_605),
.B(n_554),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_599),
.B(n_579),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_589),
.A2(n_548),
.B(n_556),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_581),
.B(n_518),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_627),
.B(n_559),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_606),
.B(n_583),
.C(n_585),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_632),
.B(n_633),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_616),
.B(n_583),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_606),
.B(n_582),
.C(n_584),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_636),
.B(n_638),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_SL g637 ( 
.A1(n_609),
.A2(n_592),
.B1(n_597),
.B2(n_533),
.Y(n_637)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_637),
.Y(n_649)
);

CKINVDCx16_ASAP7_75t_R g638 ( 
.A(n_622),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_639),
.B(n_641),
.Y(n_659)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_640),
.B(n_613),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_609),
.B(n_600),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_610),
.B(n_535),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_642),
.B(n_643),
.Y(n_655)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_615),
.B(n_559),
.C(n_602),
.Y(n_643)
);

INVxp33_ASAP7_75t_L g661 ( 
.A(n_644),
.Y(n_661)
);

XOR2xp5_ASAP7_75t_L g646 ( 
.A(n_612),
.B(n_577),
.Y(n_646)
);

XNOR2xp5_ASAP7_75t_L g656 ( 
.A(n_646),
.B(n_617),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_SL g647 ( 
.A1(n_628),
.A2(n_620),
.B1(n_607),
.B2(n_621),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_SL g670 ( 
.A1(n_647),
.A2(n_644),
.B1(n_631),
.B2(n_533),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_SL g667 ( 
.A(n_648),
.B(n_652),
.Y(n_667)
);

XOR2xp5_ASAP7_75t_L g651 ( 
.A(n_630),
.B(n_611),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_651),
.Y(n_666)
);

BUFx24_ASAP7_75t_SL g652 ( 
.A(n_629),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_632),
.B(n_618),
.C(n_626),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_653),
.B(n_654),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_635),
.B(n_618),
.C(n_623),
.Y(n_654)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_656),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_SL g657 ( 
.A1(n_634),
.A2(n_624),
.B(n_619),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_657),
.B(n_660),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_645),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_650),
.B(n_653),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_662),
.B(n_665),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_659),
.B(n_635),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_658),
.B(n_631),
.Y(n_669)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_669),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g675 ( 
.A1(n_670),
.A2(n_651),
.B1(n_640),
.B2(n_636),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_661),
.A2(n_646),
.B(n_643),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_671),
.A2(n_656),
.B(n_661),
.Y(n_673)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_654),
.Y(n_672)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_672),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_673),
.A2(n_674),
.B(n_679),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_SL g674 ( 
.A1(n_668),
.A2(n_655),
.B(n_649),
.Y(n_674)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_675),
.Y(n_681)
);

XNOR2xp5_ASAP7_75t_L g677 ( 
.A(n_671),
.B(n_516),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_677),
.B(n_666),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_664),
.B(n_663),
.Y(n_679)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_680),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_682),
.Y(n_685)
);

AOI322xp5_ASAP7_75t_L g686 ( 
.A1(n_684),
.A2(n_679),
.A3(n_666),
.B1(n_676),
.B2(n_678),
.C1(n_667),
.C2(n_295),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_686),
.B(n_683),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_SL g688 ( 
.A1(n_687),
.A2(n_685),
.B(n_681),
.Y(n_688)
);

BUFx24_ASAP7_75t_SL g689 ( 
.A(n_688),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_689),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_690),
.A2(n_356),
.B(n_295),
.Y(n_691)
);


endmodule