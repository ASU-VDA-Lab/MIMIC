module fake_jpeg_11256_n_120 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_120);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_34),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_52),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_57),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_55),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_56),
.B(n_58),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_47),
.B1(n_38),
.B2(n_39),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_67),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_39),
.B1(n_40),
.B2(n_50),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_50),
.B1(n_46),
.B2(n_41),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_49),
.B1(n_48),
.B2(n_44),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_42),
.B1(n_46),
.B2(n_17),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_16),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_1),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_74),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_1),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_8),
.B(n_9),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_2),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_77),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_2),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_3),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_80),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_3),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_4),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_82),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_6),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_65),
.Y(n_84)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_69),
.B(n_59),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_88),
.B(n_91),
.Y(n_105)
);

OR2x2_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_72),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_70),
.B(n_7),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_25),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_102),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_36),
.C(n_14),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_106),
.C(n_108),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_10),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_103),
.B(n_107),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_35),
.C(n_18),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_15),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_19),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_96),
.B(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_100),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_114),
.C(n_111),
.Y(n_115)
);

OAI322xp33_ASAP7_75t_L g114 ( 
.A1(n_110),
.A2(n_106),
.A3(n_101),
.B1(n_87),
.B2(n_104),
.C1(n_96),
.C2(n_30),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_112),
.C(n_104),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_85),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_21),
.C(n_22),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_27),
.B(n_28),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_29),
.Y(n_120)
);


endmodule