module fake_jpeg_31805_n_115 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_115);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_115;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_5),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_5),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_7),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_21),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_7),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_37),
.B(n_49),
.Y(n_62)
);

XNOR2x1_ASAP7_75t_SL g38 ( 
.A(n_35),
.B(n_19),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_50),
.Y(n_65)
);

AO22x2_ASAP7_75t_L g41 ( 
.A1(n_27),
.A2(n_16),
.B1(n_25),
.B2(n_13),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_42),
.B1(n_44),
.B2(n_50),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_31),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_19),
.B(n_20),
.C(n_17),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_13),
.B(n_31),
.Y(n_57)
);

AO22x2_ASAP7_75t_L g50 ( 
.A1(n_28),
.A2(n_13),
.B1(n_12),
.B2(n_3),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_56),
.Y(n_75)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_41),
.B1(n_47),
.B2(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_50),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_20),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_10),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_8),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_31),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_65),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_0),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_69),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_0),
.Y(n_69)
);

AND2x6_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_57),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_74),
.B(n_69),
.C(n_56),
.Y(n_86)
);

AND2x6_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_38),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_64),
.B(n_68),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_81),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_87),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_90),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_80),
.A2(n_45),
.B1(n_39),
.B2(n_54),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_75),
.B1(n_71),
.B2(n_4),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_72),
.B(n_12),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_1),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_91),
.B(n_4),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_70),
.B1(n_72),
.B2(n_74),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_93),
.A2(n_86),
.B1(n_90),
.B2(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_91),
.C(n_89),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_101),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_92),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_102),
.B(n_103),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_88),
.C(n_84),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_96),
.B1(n_92),
.B2(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_8),
.Y(n_109)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

AO21x1_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_98),
.B(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_109),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_106),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_111),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_11),
.Y(n_115)
);


endmodule