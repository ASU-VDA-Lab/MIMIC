module fake_jpeg_25006_n_297 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_20),
.B(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_41),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_32),
.B1(n_25),
.B2(n_27),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_43),
.A2(n_29),
.B1(n_27),
.B2(n_34),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_55),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_47),
.B(n_16),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_20),
.B1(n_30),
.B2(n_16),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_21),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_29),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_56),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_27),
.B1(n_32),
.B2(n_25),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_29),
.B1(n_40),
.B2(n_36),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_55),
.B1(n_54),
.B2(n_52),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_71),
.B1(n_84),
.B2(n_86),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_65),
.A2(n_69),
.B1(n_22),
.B2(n_23),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_30),
.B1(n_21),
.B2(n_26),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_76),
.Y(n_95)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_24),
.Y(n_76)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_57),
.B1(n_19),
.B2(n_46),
.Y(n_102)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_37),
.B(n_26),
.C(n_42),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_61),
.B(n_46),
.C(n_51),
.Y(n_114)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_56),
.B1(n_58),
.B2(n_48),
.Y(n_84)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_88),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_68),
.B(n_28),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_90),
.B(n_92),
.Y(n_123)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_91),
.B(n_97),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_68),
.B(n_28),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_35),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_96),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_65),
.B(n_24),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_57),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_101),
.B(n_110),
.Y(n_140)
);

AO21x1_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_107),
.B(n_112),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_65),
.A2(n_78),
.B1(n_75),
.B2(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_39),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_79),
.Y(n_141)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_SL g112 ( 
.A(n_71),
.B(n_28),
.C(n_31),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_61),
.B(n_53),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_139),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_78),
.C(n_83),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_122),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_86),
.B1(n_84),
.B2(n_64),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_117),
.A2(n_118),
.B1(n_89),
.B2(n_108),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_64),
.B1(n_80),
.B2(n_67),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_0),
.B(n_1),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_120),
.A2(n_121),
.B(n_96),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_101),
.B(n_94),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_44),
.C(n_51),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_124),
.B(n_134),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_98),
.B(n_28),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_136),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_66),
.B1(n_67),
.B2(n_87),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_131),
.B1(n_137),
.B2(n_142),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_111),
.A2(n_66),
.B1(n_77),
.B2(n_79),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_SL g161 ( 
.A(n_130),
.B(n_103),
.C(n_108),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_19),
.B1(n_73),
.B2(n_31),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_141),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_53),
.C(n_44),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_100),
.A2(n_31),
.B1(n_33),
.B2(n_18),
.Y(n_137)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_31),
.B1(n_33),
.B2(n_18),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_102),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_143),
.A2(n_146),
.B(n_156),
.Y(n_191)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_145),
.Y(n_186)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_98),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_95),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_149),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_125),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_151),
.B(n_15),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_167),
.B1(n_172),
.B2(n_142),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_154),
.A2(n_160),
.B(n_161),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_129),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_155),
.B(n_157),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_121),
.A2(n_99),
.B(n_89),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_166),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_138),
.B(n_13),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_170),
.Y(n_190)
);

AOI32xp33_ASAP7_75t_L g160 ( 
.A1(n_128),
.A2(n_112),
.A3(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_113),
.B1(n_33),
.B2(n_18),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_113),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_134),
.A2(n_33),
.B1(n_18),
.B2(n_79),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_120),
.A2(n_77),
.B(n_1),
.Y(n_168)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_116),
.B(n_0),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_171),
.A2(n_138),
.B1(n_122),
.B2(n_119),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_132),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_169),
.A2(n_132),
.B1(n_130),
.B2(n_133),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_181),
.B1(n_198),
.B2(n_172),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_174),
.A2(n_193),
.B1(n_196),
.B2(n_144),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_176),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_123),
.C(n_125),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_123),
.C(n_131),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_180),
.Y(n_203)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_170),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_187),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_126),
.C(n_137),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_164),
.A2(n_133),
.B1(n_119),
.B2(n_2),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_133),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_182),
.A2(n_143),
.B(n_146),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_177),
.Y(n_200)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_188),
.B(n_151),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_145),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_152),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_195),
.A2(n_162),
.B1(n_163),
.B2(n_171),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_165),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_198)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_200),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_201),
.A2(n_211),
.B(n_213),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_173),
.A2(n_143),
.B1(n_153),
.B2(n_158),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_202),
.A2(n_184),
.B1(n_192),
.B2(n_183),
.Y(n_231)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_157),
.Y(n_206)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_197),
.B(n_159),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_207),
.B(n_221),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_208),
.A2(n_210),
.B1(n_181),
.B2(n_184),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_216),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_182),
.A2(n_156),
.B(n_154),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_220),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_174),
.A2(n_162),
.B1(n_168),
.B2(n_160),
.Y(n_215)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_150),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_217),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_195),
.A2(n_168),
.B1(n_161),
.B2(n_167),
.Y(n_218)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_146),
.Y(n_219)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_182),
.Y(n_220)
);

NAND3xp33_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_12),
.C(n_11),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_178),
.C(n_180),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_216),
.C(n_203),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_227),
.A2(n_201),
.B1(n_194),
.B2(n_213),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_192),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_236),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_231),
.A2(n_208),
.B1(n_183),
.B2(n_194),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_191),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_237),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_185),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_240),
.Y(n_254)
);

O2A1O1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_220),
.B(n_191),
.C(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_244),
.B(n_245),
.Y(n_265)
);

BUFx24_ASAP7_75t_SL g246 ( 
.A(n_235),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_246),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_199),
.Y(n_247)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_253),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_211),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_251),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_238),
.A2(n_202),
.B1(n_205),
.B2(n_204),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_212),
.C(n_187),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_228),
.C(n_226),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_R g257 ( 
.A1(n_243),
.A2(n_239),
.B(n_228),
.Y(n_257)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_262),
.C(n_248),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_226),
.B(n_231),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_229),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_236),
.C(n_232),
.Y(n_262)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_264),
.Y(n_269)
);

OAI21x1_ASAP7_75t_SL g266 ( 
.A1(n_258),
.A2(n_251),
.B(n_250),
.Y(n_266)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_266),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_268),
.C(n_274),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_262),
.C(n_261),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_254),
.A2(n_233),
.B1(n_241),
.B2(n_249),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_270),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_260),
.A2(n_227),
.B1(n_179),
.B2(n_249),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_273),
.Y(n_280)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_256),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_229),
.C(n_209),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_275),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_271),
.A2(n_265),
.B1(n_260),
.B2(n_263),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_279),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_274),
.A2(n_261),
.B(n_263),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_10),
.Y(n_288)
);

A2O1A1O1Ixp25_ASAP7_75t_L g279 ( 
.A1(n_269),
.A2(n_259),
.B(n_264),
.C(n_198),
.D(n_10),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_269),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_285),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_282),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_280),
.B(n_278),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_288),
.C(n_281),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_289),
.A2(n_290),
.B(n_12),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_12),
.C(n_5),
.Y(n_290)
);

OAI311xp33_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_291),
.A3(n_5),
.B1(n_7),
.C1(n_8),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_4),
.C(n_5),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_7),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_9),
.B(n_7),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_8),
.C(n_9),
.Y(n_297)
);


endmodule