module real_jpeg_24977_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_1),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_1),
.A2(n_58),
.B1(n_61),
.B2(n_66),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_1),
.A2(n_38),
.B1(n_40),
.B2(n_58),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_1),
.A2(n_26),
.B1(n_32),
.B2(n_58),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_2),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_2),
.A2(n_37),
.B1(n_61),
.B2(n_66),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_2),
.A2(n_26),
.B1(n_32),
.B2(n_37),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_6),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_6),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_6),
.A2(n_61),
.B1(n_66),
.B2(n_72),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_6),
.A2(n_38),
.B1(n_40),
.B2(n_72),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_6),
.A2(n_26),
.B1(n_32),
.B2(n_72),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_7),
.A2(n_56),
.B1(n_131),
.B2(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_7),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_7),
.A2(n_61),
.B1(n_66),
.B2(n_145),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_7),
.A2(n_38),
.B1(n_40),
.B2(n_145),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_7),
.A2(n_26),
.B1(n_32),
.B2(n_145),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_8),
.A2(n_38),
.B1(n_40),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_8),
.A2(n_26),
.B1(n_32),
.B2(n_47),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_8),
.A2(n_47),
.B1(n_61),
.B2(n_66),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_11),
.B(n_54),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_11),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_11),
.B(n_60),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_11),
.B(n_38),
.C(n_81),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_11),
.A2(n_61),
.B1(n_66),
.B2(n_198),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_11),
.B(n_122),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_11),
.A2(n_38),
.B1(n_40),
.B2(n_198),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_11),
.B(n_26),
.C(n_43),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_11),
.A2(n_25),
.B(n_259),
.Y(n_284)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_13),
.A2(n_56),
.B1(n_71),
.B2(n_107),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_13),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_13),
.A2(n_61),
.B1(n_66),
.B2(n_107),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_13),
.A2(n_38),
.B1(n_40),
.B2(n_107),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_13),
.A2(n_26),
.B1(n_32),
.B2(n_107),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_14),
.A2(n_61),
.B1(n_66),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_14),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_14),
.A2(n_38),
.B1(n_40),
.B2(n_85),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_14),
.A2(n_56),
.B1(n_85),
.B2(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_14),
.A2(n_26),
.B1(n_32),
.B2(n_85),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_15),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_15),
.A2(n_33),
.B1(n_38),
.B2(n_40),
.Y(n_90)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_16),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_16),
.A2(n_167),
.B1(n_271),
.B2(n_273),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_135),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_133),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_111),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_21),
.B(n_111),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_76),
.C(n_92),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_22),
.A2(n_76),
.B1(n_77),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_22),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_49),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_23),
.A2(n_24),
.B(n_51),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_24),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_24),
.A2(n_34),
.B1(n_35),
.B2(n_50),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B(n_31),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_25),
.A2(n_28),
.B1(n_31),
.B2(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_25),
.A2(n_28),
.B1(n_97),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_25),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_25),
.A2(n_169),
.B1(n_171),
.B2(n_207),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_25),
.B(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_25),
.A2(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_26),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_45)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_27),
.Y(n_227)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_30),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_30),
.B(n_198),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_32),
.B(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_41),
.B1(n_46),
.B2(n_48),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_36),
.A2(n_41),
.B1(n_48),
.B2(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_38),
.A2(n_40),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_38),
.B(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_41),
.A2(n_48),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_41),
.B(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_41),
.A2(n_48),
.B1(n_231),
.B2(n_233),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.Y(n_41)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_45),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_45),
.A2(n_88),
.B1(n_101),
.B2(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_45),
.A2(n_155),
.B(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_45),
.A2(n_194),
.B(n_232),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_45),
.B(n_198),
.Y(n_278)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_48),
.B(n_195),
.Y(n_247)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_59),
.B(n_67),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_53),
.A2(n_59),
.B1(n_108),
.B2(n_130),
.Y(n_129)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_64),
.B1(n_65),
.B2(n_71),
.Y(n_75)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_59),
.B(n_69),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_59),
.A2(n_67),
.B(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_60),
.A2(n_74),
.B1(n_106),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_60)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_66),
.B1(n_81),
.B2(n_82),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g175 ( 
.A(n_61),
.B(n_65),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_61),
.B(n_222),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI32xp33_ASAP7_75t_L g173 ( 
.A1(n_64),
.A2(n_66),
.A3(n_71),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_74),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g197 ( 
.A1(n_73),
.A2(n_198),
.B(n_199),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_74),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_74),
.A2(n_110),
.B(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_87),
.B(n_91),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_87),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_86),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_103),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_79),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_79),
.A2(n_162),
.B(n_164),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g235 ( 
.A1(n_79),
.A2(n_164),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_80),
.A2(n_103),
.B(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_80),
.A2(n_148),
.B(n_203),
.Y(n_202)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_86),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_88),
.A2(n_246),
.B(n_247),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_88),
.A2(n_247),
.B(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_90),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_92),
.A2(n_93),
.B1(n_310),
.B2(n_312),
.Y(n_309)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_102),
.C(n_104),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_94),
.A2(n_95),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_96),
.A2(n_98),
.B1(n_99),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_96),
.Y(n_157)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_102),
.B(n_104),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B(n_109),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_129),
.B2(n_132),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_125),
.B1(n_126),
.B2(n_128),
.Y(n_118)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_121),
.A2(n_122),
.B1(n_163),
.B2(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_122),
.B(n_149),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_129),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_308),
.B(n_314),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_183),
.B(n_307),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_176),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_138),
.B(n_176),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_156),
.C(n_158),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_139),
.A2(n_140),
.B1(n_156),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_150),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_147),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_146),
.C(n_150),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_151),
.B(n_154),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_167),
.B1(n_168),
.B2(n_170),
.Y(n_166)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_156),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_158),
.B(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.C(n_165),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_159),
.B(n_161),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_165),
.B(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_173),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_173),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_171),
.A2(n_272),
.B(n_280),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_174),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_182),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_178),
.B(n_179),
.C(n_182),
.Y(n_313)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_214),
.B(n_301),
.C(n_306),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_208),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_208),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_200),
.C(n_201),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_186),
.A2(n_187),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_196),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_192),
.C(n_196),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_191),
.Y(n_203)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_200),
.B(n_201),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.C(n_206),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_241),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_206),
.Y(n_241)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_209),
.B(n_212),
.C(n_213),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_295),
.B(n_300),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_248),
.B(n_294),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_237),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_219),
.B(n_237),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_230),
.C(n_234),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_220),
.B(n_290),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_223),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B(n_228),
.Y(n_223)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_228),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_229),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_230),
.A2(n_234),
.B1(n_235),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_230),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_233),
.Y(n_246)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_242),
.B2(n_243),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_238),
.B(n_244),
.C(n_245),
.Y(n_299)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_288),
.B(n_293),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_268),
.B(n_287),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_262),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_262),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_257),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_253),
.B(n_256),
.C(n_257),
.Y(n_292)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_258),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_266),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_266),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_276),
.B(n_286),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_274),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_274),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_281),
.B(n_285),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_279),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_292),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_292),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_299),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_299),
.Y(n_300)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_303),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_313),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_313),
.Y(n_314)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_310),
.Y(n_312)
);


endmodule