module fake_jpeg_17760_n_49 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_2),
.B(n_4),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_6),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_7),
.B(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_17),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_9),
.A2(n_11),
.B1(n_13),
.B2(n_7),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_16),
.B(n_18),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_0),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_13),
.B1(n_8),
.B2(n_14),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_0),
.Y(n_19)
);

AND2x2_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_20),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_1),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_8),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_22),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_12),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_15),
.B(n_3),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_12),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_21),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_17),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_27),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_22),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_16),
.B1(n_18),
.B2(n_6),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_26),
.B(n_6),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_37),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_31),
.C(n_10),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_42),
.B(n_35),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_37),
.B1(n_43),
.B2(n_42),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_40),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_46),
.B(n_44),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_48),
.Y(n_49)
);


endmodule