module fake_jpeg_6292_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_14),
.B(n_5),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_42),
.Y(n_47)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_38),
.A2(n_40),
.B1(n_20),
.B2(n_21),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_39),
.Y(n_56)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_43),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_0),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_19),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_22),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_54),
.Y(n_99)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_22),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_58),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_21),
.B1(n_33),
.B2(n_20),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_67),
.B1(n_72),
.B2(n_28),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_20),
.B1(n_33),
.B2(n_21),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_62),
.A2(n_24),
.B(n_26),
.C(n_29),
.Y(n_97)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_66),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_37),
.A2(n_20),
.B1(n_33),
.B2(n_22),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_45),
.B1(n_28),
.B2(n_25),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_28),
.B1(n_25),
.B2(n_27),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_40),
.B1(n_45),
.B2(n_23),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_86),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_78),
.B(n_29),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_41),
.C(n_44),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_41),
.C(n_23),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_32),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_32),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_24),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_29),
.B(n_24),
.Y(n_128)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_88),
.Y(n_104)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_90),
.A2(n_57),
.B1(n_19),
.B2(n_27),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_55),
.A2(n_25),
.B1(n_23),
.B2(n_27),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_96),
.Y(n_112)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_19),
.B(n_51),
.C(n_62),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_108),
.B(n_128),
.Y(n_134)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_101),
.B(n_103),
.Y(n_145)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_52),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_107),
.Y(n_129)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_106),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_49),
.Y(n_107)
);

AO22x1_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_51),
.B1(n_36),
.B2(n_34),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_82),
.C(n_99),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_111),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_69),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_83),
.Y(n_113)
);

INVx3_ASAP7_75t_SL g143 ( 
.A(n_113),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_92),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_114),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_70),
.Y(n_115)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_46),
.Y(n_116)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_69),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_125),
.Y(n_136)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_118),
.A2(n_120),
.B1(n_122),
.B2(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_26),
.Y(n_140)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_124),
.B1(n_82),
.B2(n_84),
.Y(n_137)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_86),
.A2(n_36),
.B(n_57),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_39),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_92),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_113),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_122),
.B1(n_103),
.B2(n_104),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_133),
.A2(n_100),
.B1(n_123),
.B2(n_120),
.Y(n_157)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_135),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_114),
.B1(n_83),
.B2(n_98),
.Y(n_170)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_139),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_127),
.Y(n_167)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_144),
.B(n_146),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_102),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_147),
.B(n_106),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_84),
.C(n_91),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_153),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_119),
.A2(n_64),
.B1(n_63),
.B2(n_46),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_91),
.C(n_93),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_154),
.A2(n_124),
.B(n_101),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_164),
.Y(n_206)
);

AO22x1_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_124),
.B1(n_128),
.B2(n_121),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_159),
.A2(n_183),
.B(n_140),
.Y(n_199)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_160),
.B(n_161),
.Y(n_209)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_137),
.A2(n_124),
.B1(n_117),
.B2(n_125),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_163),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_165),
.B(n_169),
.Y(n_197)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_166),
.B(n_167),
.CI(n_178),
.CON(n_211),
.SN(n_211)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_176),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_98),
.B1(n_93),
.B2(n_89),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_150),
.A2(n_118),
.B1(n_36),
.B2(n_65),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_144),
.A2(n_73),
.B1(n_65),
.B2(n_26),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_180),
.A2(n_142),
.B1(n_153),
.B2(n_149),
.Y(n_187)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_39),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_187),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_157),
.A2(n_156),
.B1(n_134),
.B2(n_145),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_188),
.A2(n_198),
.B1(n_210),
.B2(n_168),
.Y(n_223)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_189),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_136),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_191),
.C(n_196),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_136),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_162),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_192),
.B(n_200),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_131),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_159),
.A2(n_134),
.B1(n_142),
.B2(n_146),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_204),
.B(n_206),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_182),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_203),
.Y(n_212)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_159),
.A2(n_140),
.B(n_152),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_39),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_179),
.A2(n_138),
.B1(n_141),
.B2(n_135),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_228),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_202),
.A2(n_179),
.B1(n_169),
.B2(n_165),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_214),
.A2(n_221),
.B1(n_225),
.B2(n_237),
.Y(n_243)
);

BUFx12_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_216),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_193),
.B(n_161),
.Y(n_219)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_219),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_210),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_220),
.B(n_232),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_168),
.B1(n_184),
.B2(n_160),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_163),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_226),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_223),
.A2(n_231),
.B1(n_189),
.B2(n_56),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_205),
.B(n_178),
.Y(n_224)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_194),
.A2(n_176),
.B1(n_178),
.B2(n_81),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_39),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_229),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_81),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_199),
.A2(n_204),
.B(n_198),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_234),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_195),
.A2(n_56),
.B(n_39),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_0),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_188),
.A2(n_211),
.B(n_185),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_222),
.B(n_211),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_240),
.B(n_249),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_196),
.C(n_211),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_246),
.C(n_248),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_245),
.A2(n_215),
.B1(n_214),
.B2(n_233),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_56),
.C(n_16),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_227),
.B(n_10),
.Y(n_247)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_247),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_16),
.C(n_30),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_230),
.B(n_16),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_30),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_253),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_216),
.Y(n_252)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_30),
.Y(n_253)
);

NAND3xp33_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_16),
.C(n_18),
.Y(n_256)
);

AO21x1_ASAP7_75t_L g261 ( 
.A1(n_256),
.A2(n_258),
.B(n_259),
.Y(n_261)
);

XOR2x1_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_16),
.Y(n_258)
);

NAND3xp33_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_16),
.C(n_8),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_74),
.C(n_1),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_232),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_263),
.A2(n_274),
.B1(n_218),
.B2(n_249),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_275),
.C(n_250),
.Y(n_283)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_257),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_216),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_243),
.A2(n_215),
.B1(n_237),
.B2(n_212),
.Y(n_266)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_258),
.A2(n_212),
.B1(n_231),
.B2(n_219),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_267),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_228),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_273),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_239),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_276),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_225),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_254),
.A2(n_259),
.B1(n_218),
.B2(n_235),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_236),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_238),
.Y(n_276)
);

OAI21x1_ASAP7_75t_L g278 ( 
.A1(n_256),
.A2(n_229),
.B(n_216),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_278),
.A2(n_7),
.B(n_14),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_255),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_8),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_240),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_277),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_291),
.C(n_294),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_264),
.B(n_260),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_284),
.B(n_288),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_272),
.Y(n_285)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_286),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_263),
.A2(n_244),
.B1(n_74),
.B2(n_2),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_290),
.A2(n_295),
.B(n_261),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_273),
.C(n_269),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_7),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_292),
.B(n_2),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_261),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_0),
.C(n_1),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_270),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_296),
.A2(n_300),
.B(n_302),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_298),
.B(n_6),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_262),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_262),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_303),
.A2(n_309),
.B(n_4),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_307),
.C(n_308),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_3),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_282),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_277),
.C(n_4),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_294),
.B(n_3),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_290),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_312),
.Y(n_322)
);

AO21x1_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_283),
.B(n_301),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_314),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_287),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_297),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_15),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_4),
.C(n_5),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_12),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_319),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_307),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_6),
.Y(n_324)
);

NOR3xp33_ASAP7_75t_SL g321 ( 
.A(n_315),
.B(n_304),
.C(n_11),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_324),
.Y(n_333)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_326),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_316),
.B(n_12),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_328),
.C(n_310),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_330),
.C(n_332),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_311),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_13),
.Y(n_332)
);

AOI321xp33_ASAP7_75t_L g335 ( 
.A1(n_333),
.A2(n_13),
.A3(n_15),
.B1(n_325),
.B2(n_327),
.C(n_331),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_335),
.Y(n_336)
);

AO21x1_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_333),
.B(n_334),
.Y(n_337)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_337),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_13),
.Y(n_339)
);


endmodule