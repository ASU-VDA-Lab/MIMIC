module fake_jpeg_8278_n_227 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_44),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_20),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_25),
.B1(n_18),
.B2(n_34),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_62),
.B1(n_70),
.B2(n_19),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_32),
.B(n_18),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_33),
.B(n_28),
.C(n_27),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_50),
.B(n_63),
.Y(n_89)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_57),
.Y(n_71)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_58),
.B(n_59),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_60),
.B(n_0),
.Y(n_94)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

OR2x2_ASAP7_75t_SL g99 ( 
.A(n_61),
.B(n_67),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_25),
.B1(n_19),
.B2(n_34),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_30),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_31),
.C(n_20),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_26),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_35),
.A2(n_33),
.B1(n_28),
.B2(n_19),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_72),
.A2(n_51),
.B1(n_67),
.B2(n_65),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_27),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_74),
.B(n_77),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_38),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_93),
.Y(n_106)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_78),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_30),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_80),
.Y(n_116)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_81),
.A2(n_85),
.B1(n_87),
.B2(n_56),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_31),
.Y(n_82)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_51),
.Y(n_83)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_29),
.B1(n_17),
.B2(n_22),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_24),
.B(n_1),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_5),
.B(n_8),
.C(n_9),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_56),
.A2(n_29),
.B1(n_24),
.B2(n_2),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_24),
.B1(n_1),
.B2(n_3),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_3),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_96),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_4),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_48),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_101),
.B1(n_10),
.B2(n_15),
.Y(n_121)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_55),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_53),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_102),
.B(n_121),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_104),
.A2(n_71),
.B(n_92),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_81),
.A2(n_75),
.B1(n_86),
.B2(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_8),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_115),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_8),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_9),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_125),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_72),
.A2(n_54),
.B1(n_12),
.B2(n_14),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_87),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_10),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_120),
.A2(n_92),
.B(n_96),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_85),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_99),
.Y(n_126)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_137),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_130),
.B(n_136),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_148),
.B1(n_105),
.B2(n_91),
.Y(n_155)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_99),
.Y(n_132)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_132),
.A2(n_120),
.B(n_117),
.C(n_105),
.D(n_76),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_77),
.Y(n_134)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_145),
.B(n_117),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_93),
.Y(n_139)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_109),
.A2(n_106),
.B(n_110),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_140),
.A2(n_120),
.B(n_104),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_116),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_142),
.B(n_144),
.Y(n_165)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_92),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_147),
.Y(n_168)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_124),
.C(n_118),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_154),
.C(n_157),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_164),
.B(n_145),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_153),
.B(n_159),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_123),
.C(n_121),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_155),
.A2(n_135),
.B1(n_143),
.B2(n_142),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_123),
.C(n_103),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_137),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_147),
.C(n_133),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_136),
.C(n_133),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_141),
.B(n_113),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_141),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_152),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_138),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_165),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_181),
.Y(n_190)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_171),
.A2(n_183),
.B1(n_184),
.B2(n_153),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_154),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_180),
.C(n_182),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_163),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_160),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_177),
.B(n_178),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_149),
.B(n_130),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_132),
.C(n_143),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_157),
.C(n_164),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_167),
.A2(n_135),
.B1(n_148),
.B2(n_126),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_175),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_185),
.B(n_189),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_191),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_184),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_150),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_166),
.C(n_168),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_194),
.C(n_173),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_114),
.B1(n_80),
.B2(n_128),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_179),
.A2(n_151),
.B1(n_156),
.B2(n_137),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_195),
.A2(n_170),
.B(n_171),
.Y(n_198)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_198),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_190),
.A2(n_180),
.B(n_176),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_202),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_187),
.B(n_174),
.Y(n_202)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_172),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_198),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_114),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_192),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_196),
.A2(n_128),
.B(n_96),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_199),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_191),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_206),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

AOI31xp67_ASAP7_75t_SL g213 ( 
.A1(n_201),
.A2(n_194),
.A3(n_186),
.B(n_197),
.Y(n_213)
);

AO21x1_ASAP7_75t_L g217 ( 
.A1(n_213),
.A2(n_203),
.B(n_78),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_186),
.C(n_199),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_214),
.B(n_216),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_215),
.Y(n_219)
);

NOR2x1_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_207),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_207),
.C(n_210),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_220),
.A2(n_218),
.B(n_84),
.Y(n_223)
);

OAI21x1_ASAP7_75t_L g224 ( 
.A1(n_221),
.A2(n_100),
.B(n_220),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_224),
.Y(n_225)
);

NOR3xp33_ASAP7_75t_SL g226 ( 
.A(n_225),
.B(n_222),
.C(n_221),
.Y(n_226)
);

FAx1_ASAP7_75t_SL g227 ( 
.A(n_226),
.B(n_219),
.CI(n_221),
.CON(n_227),
.SN(n_227)
);


endmodule