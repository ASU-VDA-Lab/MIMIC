module fake_jpeg_9649_n_297 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_40),
.B(n_35),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_44),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_19),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_51),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_38),
.B1(n_18),
.B2(n_40),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_70),
.B1(n_30),
.B2(n_22),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_19),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_35),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_52),
.B(n_61),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_18),
.B1(n_29),
.B2(n_23),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_53),
.A2(n_69),
.B1(n_34),
.B2(n_25),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_26),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_59),
.B(n_67),
.Y(n_97)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_30),
.Y(n_78)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_SL g66 ( 
.A1(n_36),
.A2(n_26),
.B(n_23),
.Y(n_66)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_68),
.B(n_34),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_36),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_39),
.A2(n_18),
.B1(n_29),
.B2(n_32),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_37),
.A2(n_29),
.B1(n_21),
.B2(n_32),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_27),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_47),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_72),
.A2(n_99),
.B1(n_65),
.B2(n_61),
.Y(n_109)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_74),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_77),
.Y(n_124)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_107),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_31),
.B(n_25),
.C(n_27),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_SL g119 ( 
.A(n_79),
.B(n_87),
.C(n_1),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_80),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_95),
.B1(n_98),
.B2(n_28),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_31),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_84),
.B(n_90),
.Y(n_121)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_86),
.Y(n_132)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_0),
.B(n_1),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_19),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_91),
.B(n_96),
.Y(n_134)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_50),
.A2(n_33),
.B1(n_20),
.B2(n_19),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_64),
.A2(n_33),
.B1(n_19),
.B2(n_17),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_58),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_64),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_17),
.Y(n_104)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_33),
.C(n_28),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_109),
.A2(n_114),
.B1(n_116),
.B2(n_130),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_111),
.B(n_94),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_72),
.A2(n_65),
.B1(n_28),
.B2(n_3),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_1),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_131),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_71),
.A2(n_99),
.B1(n_95),
.B2(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_117),
.B(n_82),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_119),
.A2(n_6),
.B(n_7),
.Y(n_162)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_129),
.B(n_89),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_106),
.A2(n_28),
.B1(n_3),
.B2(n_5),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_2),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_87),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_135),
.A2(n_96),
.B(n_105),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_119),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_152),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_107),
.C(n_103),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_147),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_139),
.A2(n_158),
.B(n_118),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_131),
.B(n_79),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_140),
.B(n_141),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_112),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_124),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_146),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_115),
.B(n_116),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_143),
.B(n_144),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_78),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_85),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_101),
.C(n_102),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_83),
.C(n_100),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_148),
.B(n_11),
.Y(n_196)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_150),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_109),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_121),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_8),
.Y(n_182)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_157),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_154),
.A2(n_162),
.B(n_123),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_80),
.B(n_108),
.C(n_89),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_156),
.A2(n_113),
.B1(n_120),
.B2(n_10),
.Y(n_184)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_135),
.A2(n_93),
.B(n_108),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_77),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_159),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_160),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_161),
.B(n_118),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_125),
.B(n_7),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_164),
.Y(n_180)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_129),
.B(n_127),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_165),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_126),
.B(n_7),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_8),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_150),
.A2(n_130),
.B1(n_136),
.B2(n_127),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_168),
.A2(n_185),
.B1(n_155),
.B2(n_144),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_173),
.B(n_145),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_139),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_178),
.B(n_186),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_113),
.B(n_123),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_181),
.A2(n_192),
.B(n_162),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_187),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_191),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_152),
.A2(n_120),
.B1(n_9),
.B2(n_10),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_189),
.Y(n_204)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_143),
.A2(n_14),
.B(n_11),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_8),
.Y(n_193)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_183),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_145),
.C(n_138),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_198),
.A2(n_177),
.B(n_169),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_199),
.B(n_211),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_207),
.Y(n_226)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_202),
.B(n_206),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_172),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_170),
.B(n_148),
.C(n_167),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_218),
.C(n_193),
.Y(n_229)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_175),
.B(n_174),
.Y(n_236)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_141),
.Y(n_213)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_214),
.A2(n_216),
.B1(n_219),
.B2(n_220),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_142),
.Y(n_215)
);

INVxp33_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_217),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_173),
.B(n_155),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_191),
.A2(n_154),
.B1(n_140),
.B2(n_149),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_170),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_229),
.C(n_238),
.Y(n_245)
);

AO21x1_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_232),
.B(n_192),
.Y(n_248)
);

AO21x1_ASAP7_75t_L g232 ( 
.A1(n_197),
.A2(n_169),
.B(n_178),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_196),
.C(n_187),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_233),
.B(n_182),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_217),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_188),
.Y(n_254)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_168),
.B1(n_186),
.B2(n_195),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_219),
.B1(n_204),
.B2(n_198),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_195),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_211),
.B(n_181),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_205),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_222),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_241),
.B(n_242),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_223),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_243),
.A2(n_255),
.B(n_189),
.Y(n_265)
);

INVxp33_ASAP7_75t_SL g244 ( 
.A(n_235),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_249),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_230),
.B(n_207),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_246),
.B(n_251),
.Y(n_262)
);

NAND4xp25_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_184),
.C(n_175),
.D(n_185),
.Y(n_247)
);

O2A1O1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_247),
.A2(n_248),
.B(n_253),
.C(n_200),
.Y(n_261)
);

INVxp33_ASAP7_75t_SL g249 ( 
.A(n_235),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_225),
.B(n_151),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_254),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_204),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_227),
.C(n_226),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_259),
.C(n_222),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_221),
.B1(n_179),
.B2(n_200),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_258),
.A2(n_267),
.B(n_247),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_229),
.C(n_201),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_261),
.A2(n_203),
.B1(n_163),
.B2(n_208),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_253),
.B(n_182),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_203),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_265),
.A2(n_268),
.B(n_166),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_257),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_240),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_243),
.A2(n_194),
.B(n_239),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_269),
.B(n_271),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_264),
.A2(n_248),
.B1(n_137),
.B2(n_166),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_270),
.A2(n_272),
.B(n_276),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_R g272 ( 
.A(n_261),
.B(n_137),
.C(n_238),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_274),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_275),
.B(n_277),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_11),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_267),
.B1(n_262),
.B2(n_256),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_278),
.B(n_12),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_266),
.Y(n_279)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_279),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_272),
.Y(n_281)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_12),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_283),
.A2(n_282),
.B(n_280),
.Y(n_286)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_286),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_289),
.B(n_290),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_271),
.B(n_275),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_13),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_13),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_295),
.C(n_293),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_291),
.A2(n_288),
.B(n_14),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_292),
.Y(n_297)
);


endmodule