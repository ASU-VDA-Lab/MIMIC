module fake_jpeg_30791_n_243 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_243);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_243;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_8),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_25),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_23),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_26),
.B(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_2),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_16),
.B1(n_18),
.B2(n_21),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_54),
.B1(n_60),
.B2(n_62),
.Y(n_71)
);

AO22x1_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_31),
.B1(n_26),
.B2(n_28),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_47),
.A2(n_40),
.B1(n_44),
.B2(n_42),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_16),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_57),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_30),
.B1(n_32),
.B2(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_55),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_59),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_16),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_37),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_30),
.B1(n_32),
.B2(n_22),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_24),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_63),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_35),
.A2(n_21),
.B1(n_25),
.B2(n_22),
.Y(n_62)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_19),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_66),
.B(n_85),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_75),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_63),
.A2(n_35),
.B1(n_34),
.B2(n_43),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_70),
.A2(n_76),
.B1(n_83),
.B2(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_19),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_36),
.B1(n_34),
.B2(n_43),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVxp67_ASAP7_75t_SL g79 ( 
.A(n_51),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_91),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_34),
.B1(n_43),
.B2(n_44),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_50),
.A2(n_36),
.B(n_24),
.C(n_17),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_56),
.B(n_17),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_86),
.B(n_87),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_55),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_89),
.A2(n_60),
.B1(n_42),
.B2(n_53),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_50),
.A2(n_32),
.B1(n_29),
.B2(n_15),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_28),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_93),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_L g93 ( 
.A(n_47),
.B(n_2),
.C(n_3),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_47),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_40),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_96),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_45),
.B(n_39),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_52),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_54),
.A2(n_31),
.B(n_4),
.C(n_5),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_98),
.B(n_4),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_58),
.B(n_3),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_5),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_101),
.A2(n_112),
.B1(n_70),
.B2(n_83),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_42),
.B(n_29),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_121),
.B(n_69),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_84),
.B1(n_73),
.B2(n_72),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_71),
.A2(n_52),
.B1(n_33),
.B2(n_15),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_84),
.B(n_5),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_124),
.B(n_6),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_51),
.B1(n_39),
.B2(n_52),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_65),
.B1(n_67),
.B2(n_88),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_72),
.Y(n_131)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_143),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_106),
.A2(n_73),
.B1(n_99),
.B2(n_82),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_147),
.B1(n_149),
.B2(n_115),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_85),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_119),
.Y(n_172)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_121),
.B(n_153),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_80),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_137),
.B(n_138),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_116),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_124),
.B(n_78),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_142),
.B(n_132),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_77),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_97),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_108),
.C(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_101),
.A2(n_89),
.B1(n_98),
.B2(n_53),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_106),
.A2(n_89),
.B1(n_64),
.B2(n_33),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_152),
.Y(n_159)
);

A2O1A1O1Ixp25_ASAP7_75t_L g151 ( 
.A1(n_117),
.A2(n_89),
.B(n_81),
.C(n_8),
.D(n_9),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_110),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_111),
.Y(n_152)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_148),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_172),
.C(n_141),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_156),
.B(n_162),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_158),
.A2(n_167),
.B(n_166),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_118),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_SL g183 ( 
.A1(n_164),
.A2(n_154),
.B(n_113),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_166),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_129),
.B1(n_109),
.B2(n_128),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_136),
.A2(n_114),
.B(n_110),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_127),
.Y(n_168)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_168),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_186),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_164),
.A2(n_151),
.B(n_147),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_183),
.B(n_160),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_174),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_180),
.A2(n_192),
.B(n_170),
.Y(n_201)
);

INVxp67_ASAP7_75t_SL g181 ( 
.A(n_159),
.Y(n_181)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_144),
.C(n_134),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_162),
.C(n_175),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_140),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_185),
.B(n_157),
.Y(n_199)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_193),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_135),
.B1(n_130),
.B2(n_102),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_189),
.A2(n_192),
.B1(n_169),
.B2(n_173),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_114),
.B(n_119),
.Y(n_192)
);

OAI321xp33_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_127),
.A3(n_113),
.B1(n_120),
.B2(n_10),
.C(n_11),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_191),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_197),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_201),
.B(n_180),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_191),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_156),
.B1(n_171),
.B2(n_172),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_198),
.A2(n_200),
.B1(n_184),
.B2(n_176),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_188),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_190),
.A2(n_170),
.B1(n_169),
.B2(n_173),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_202),
.A2(n_188),
.B1(n_189),
.B2(n_178),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_206),
.C(n_207),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_120),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_185),
.Y(n_208)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_210),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_206),
.B(n_182),
.Y(n_210)
);

BUFx24_ASAP7_75t_SL g225 ( 
.A(n_212),
.Y(n_225)
);

XNOR2x1_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_201),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_217),
.B1(n_202),
.B2(n_198),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_177),
.B(n_7),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_216),
.C(n_205),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_6),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_221),
.B(n_224),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_203),
.C(n_207),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_223),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_214),
.C(n_213),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_209),
.Y(n_228)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_228),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_225),
.A2(n_215),
.B1(n_211),
.B2(n_9),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_230),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_226),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_232),
.B(n_234),
.Y(n_237)
);

OAI221xp5_ASAP7_75t_L g235 ( 
.A1(n_229),
.A2(n_221),
.B1(n_12),
.B2(n_13),
.C(n_7),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_235),
.A2(n_229),
.B(n_12),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_231),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_236),
.B(n_238),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_240),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_239),
.Y(n_242)
);

BUFx24_ASAP7_75t_SL g243 ( 
.A(n_242),
.Y(n_243)
);


endmodule