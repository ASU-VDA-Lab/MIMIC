module fake_netlist_6_2517_n_1663 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1663);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1663;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_SL g159 ( 
.A(n_58),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_54),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_112),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_22),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_37),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_36),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_52),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_105),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_53),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_96),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_62),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_142),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_154),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_88),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_33),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_33),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_9),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_80),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_48),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_150),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_147),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_104),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_83),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_22),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_5),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_50),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_40),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_143),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_106),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_1),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_85),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_129),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_55),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_75),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_9),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_76),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_65),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_19),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_100),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_111),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_93),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_74),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_4),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_0),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_130),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_25),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_86),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_73),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_6),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_71),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_28),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_2),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_133),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_25),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_49),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_107),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_19),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_11),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_137),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_42),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_135),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_101),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_120),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_21),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_113),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_156),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_11),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_20),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_81),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_125),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_60),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_136),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_8),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g238 ( 
.A(n_47),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_144),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_128),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_127),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_10),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_99),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_21),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_110),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_2),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_92),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_5),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_72),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_56),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_8),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_59),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_90),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_0),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_42),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_66),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_139),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_29),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_63),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_95),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_35),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_103),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_138),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_15),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_1),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_36),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_20),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_41),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_7),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_122),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_27),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_117),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_116),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_43),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_141),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_27),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_4),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_28),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_98),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_114),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_37),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_109),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_23),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_67),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_38),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_108),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_40),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_121),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_14),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_78),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_41),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_82),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_13),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_68),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_35),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_131),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_6),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_3),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_61),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_32),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_45),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_39),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_152),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_97),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_44),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_149),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_51),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_87),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_13),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_140),
.Y(n_310)
);

BUFx10_ASAP7_75t_L g311 ( 
.A(n_7),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_31),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_39),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_158),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_12),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_266),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_170),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_266),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_276),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_184),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_281),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_276),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_190),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_283),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_193),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_283),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_246),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_254),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_254),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_315),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_165),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_174),
.Y(n_332)
);

INVxp33_ASAP7_75t_SL g333 ( 
.A(n_162),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_185),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_195),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_197),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_215),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_218),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_232),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_198),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_237),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_255),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_264),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_203),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_269),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_278),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_281),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_289),
.Y(n_348)
);

INVxp33_ASAP7_75t_SL g349 ( 
.A(n_162),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_187),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_295),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_302),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_193),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_194),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_271),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_204),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_271),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_211),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_226),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_226),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_262),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_262),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_163),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_212),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_168),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_173),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_305),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_214),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_178),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_217),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_220),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_166),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_281),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_179),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_180),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_225),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_229),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_219),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_191),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_233),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_196),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_235),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_305),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_312),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_247),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_249),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_200),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_201),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_205),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_209),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_227),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_318),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_318),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_324),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_377),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_367),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_324),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_367),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_383),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_365),
.Y(n_400)
);

OAI21x1_ASAP7_75t_L g401 ( 
.A1(n_383),
.A2(n_240),
.B(n_236),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_323),
.B(n_238),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_335),
.B(n_223),
.Y(n_403)
);

AND2x6_ASAP7_75t_L g404 ( 
.A(n_325),
.B(n_305),
.Y(n_404)
);

INVx6_ASAP7_75t_L g405 ( 
.A(n_354),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_382),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_386),
.Y(n_407)
);

AND2x2_ASAP7_75t_SL g408 ( 
.A(n_366),
.B(n_305),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_336),
.B(n_340),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_359),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_339),
.Y(n_411)
);

INVx6_ASAP7_75t_L g412 ( 
.A(n_354),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_344),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_356),
.B(n_223),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_353),
.B(n_194),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_325),
.B(n_234),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_358),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_364),
.B(n_234),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_359),
.Y(n_419)
);

XNOR2x2_ASAP7_75t_R g420 ( 
.A(n_317),
.B(n_3),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_369),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_339),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_360),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_328),
.B(n_230),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_368),
.B(n_304),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_369),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_360),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_325),
.B(n_304),
.Y(n_428)
);

OAI21x1_ASAP7_75t_L g429 ( 
.A1(n_361),
.A2(n_314),
.B(n_243),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_374),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_341),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_328),
.B(n_329),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_320),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_333),
.A2(n_313),
.B1(n_309),
.B2(n_300),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_370),
.B(n_159),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_371),
.B(n_241),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_376),
.Y(n_437)
);

INVx6_ASAP7_75t_L g438 ( 
.A(n_321),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_374),
.B(n_245),
.Y(n_439)
);

CKINVDCx11_ASAP7_75t_R g440 ( 
.A(n_347),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_341),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_361),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_375),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_362),
.Y(n_444)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_380),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_362),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_385),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_346),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_363),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_363),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_346),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_330),
.Y(n_452)
);

AND2x6_ASAP7_75t_L g453 ( 
.A(n_375),
.B(n_305),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_316),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_327),
.Y(n_455)
);

AND2x6_ASAP7_75t_L g456 ( 
.A(n_379),
.B(n_256),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_350),
.B(n_257),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_349),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_331),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_396),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_396),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_398),
.Y(n_462)
);

INVxp33_ASAP7_75t_L g463 ( 
.A(n_455),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_405),
.Y(n_464)
);

NAND3xp33_ASAP7_75t_L g465 ( 
.A(n_402),
.B(n_378),
.C(n_372),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_432),
.Y(n_466)
);

BUFx4f_ASAP7_75t_L g467 ( 
.A(n_456),
.Y(n_467)
);

INVxp33_ASAP7_75t_L g468 ( 
.A(n_424),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_428),
.B(n_260),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_432),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_398),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_400),
.Y(n_473)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_404),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_403),
.B(n_379),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_399),
.Y(n_476)
);

NOR2x1p5_ASAP7_75t_L g477 ( 
.A(n_445),
.B(n_163),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_398),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_433),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_408),
.B(n_263),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_414),
.B(n_381),
.Y(n_481)
);

AND3x2_ASAP7_75t_L g482 ( 
.A(n_449),
.B(n_293),
.C(n_261),
.Y(n_482)
);

OR2x6_ASAP7_75t_L g483 ( 
.A(n_445),
.B(n_329),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_427),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_427),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_427),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_427),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_433),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_427),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_R g490 ( 
.A(n_395),
.B(n_406),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_404),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_401),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_405),
.Y(n_493)
);

INVxp33_ASAP7_75t_L g494 ( 
.A(n_424),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_435),
.B(n_381),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_405),
.Y(n_496)
);

NOR2x1p5_ASAP7_75t_L g497 ( 
.A(n_445),
.B(n_175),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_421),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_408),
.B(n_387),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_425),
.B(n_373),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_426),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_444),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_408),
.B(n_387),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_405),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_444),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_418),
.B(n_384),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_416),
.B(n_351),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_444),
.Y(n_508)
);

AND2x6_ASAP7_75t_L g509 ( 
.A(n_428),
.B(n_416),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_430),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_443),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_395),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_452),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_415),
.B(n_388),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_444),
.Y(n_515)
);

OAI21xp33_ASAP7_75t_SL g516 ( 
.A1(n_457),
.A2(n_389),
.B(n_388),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_401),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_416),
.B(n_352),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_452),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_444),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g521 ( 
.A1(n_439),
.A2(n_391),
.B1(n_390),
.B2(n_389),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_442),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_412),
.Y(n_523)
);

BUFx6f_ASAP7_75t_SL g524 ( 
.A(n_428),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_436),
.B(n_390),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_416),
.B(n_391),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_409),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_442),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_442),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_410),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_459),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_410),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_419),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_428),
.B(n_456),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_456),
.B(n_189),
.Y(n_535)
);

OAI21xp33_ASAP7_75t_SL g536 ( 
.A1(n_429),
.A2(n_322),
.B(n_316),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_412),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_456),
.B(n_206),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_429),
.Y(n_539)
);

OR2x6_ASAP7_75t_L g540 ( 
.A(n_438),
.B(n_355),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_439),
.B(n_331),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_406),
.Y(n_542)
);

BUFx8_ASAP7_75t_SL g543 ( 
.A(n_407),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_419),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_439),
.B(n_275),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_454),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_412),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_423),
.Y(n_548)
);

NAND3xp33_ASAP7_75t_L g549 ( 
.A(n_415),
.B(n_222),
.C(n_192),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_454),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_407),
.Y(n_551)
);

AND2x2_ASAP7_75t_SL g552 ( 
.A(n_439),
.B(n_279),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_412),
.B(n_355),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_448),
.Y(n_554)
);

AND3x2_ASAP7_75t_L g555 ( 
.A(n_450),
.B(n_303),
.C(n_282),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_423),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_446),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_456),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_446),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_454),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_448),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_413),
.B(n_284),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_450),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_451),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_451),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_392),
.Y(n_566)
);

OR2x6_ASAP7_75t_L g567 ( 
.A(n_438),
.B(n_357),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_456),
.B(n_252),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_413),
.B(n_357),
.Y(n_569)
);

BUFx6f_ASAP7_75t_SL g570 ( 
.A(n_420),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_392),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_417),
.B(n_160),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_393),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_393),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_417),
.B(n_348),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_394),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_438),
.Y(n_577)
);

OAI21xp33_ASAP7_75t_SL g578 ( 
.A1(n_394),
.A2(n_319),
.B(n_322),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_397),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_456),
.B(n_250),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_397),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_411),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_411),
.Y(n_583)
);

OR2x6_ASAP7_75t_L g584 ( 
.A(n_438),
.B(n_332),
.Y(n_584)
);

AND3x2_ASAP7_75t_L g585 ( 
.A(n_420),
.B(n_292),
.C(n_345),
.Y(n_585)
);

AND3x2_ASAP7_75t_L g586 ( 
.A(n_422),
.B(n_348),
.C(n_345),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_422),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_431),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_437),
.B(n_253),
.Y(n_589)
);

INVx8_ASAP7_75t_L g590 ( 
.A(n_404),
.Y(n_590)
);

NOR3xp33_ASAP7_75t_L g591 ( 
.A(n_458),
.B(n_210),
.C(n_228),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_431),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_441),
.Y(n_593)
);

INVx5_ASAP7_75t_L g594 ( 
.A(n_404),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_441),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_404),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_404),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_458),
.Y(n_598)
);

NAND2xp33_ASAP7_75t_L g599 ( 
.A(n_404),
.B(n_160),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_453),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_453),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_453),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_437),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_453),
.B(n_270),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_575),
.B(n_447),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_534),
.A2(n_272),
.B(n_273),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_SL g607 ( 
.A1(n_506),
.A2(n_434),
.B1(n_447),
.B2(n_230),
.Y(n_607)
);

OAI22xp33_ASAP7_75t_L g608 ( 
.A1(n_468),
.A2(n_244),
.B1(n_298),
.B2(n_186),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_L g609 ( 
.A(n_509),
.B(n_274),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_525),
.B(n_453),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_495),
.B(n_453),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_552),
.B(n_280),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_478),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_468),
.B(n_161),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_494),
.B(n_440),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_552),
.B(n_286),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_513),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_467),
.B(n_499),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_563),
.B(n_332),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_478),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_494),
.B(n_475),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_503),
.B(n_453),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_480),
.A2(n_175),
.B1(n_176),
.B2(n_186),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_467),
.B(n_161),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_481),
.B(n_164),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_462),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_507),
.B(n_334),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_467),
.B(n_164),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_509),
.Y(n_629)
);

INVxp33_ASAP7_75t_L g630 ( 
.A(n_463),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_539),
.B(n_167),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_529),
.B(n_167),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_539),
.B(n_169),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_519),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_465),
.B(n_169),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_529),
.B(n_171),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_463),
.B(n_311),
.Y(n_637)
);

NAND3xp33_ASAP7_75t_L g638 ( 
.A(n_569),
.B(n_258),
.C(n_199),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_529),
.B(n_171),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_472),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_563),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_546),
.B(n_172),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_539),
.B(n_172),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_546),
.B(n_177),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_531),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_500),
.B(n_177),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_546),
.B(n_181),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_550),
.B(n_181),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_460),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_550),
.B(n_182),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_473),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_L g652 ( 
.A(n_509),
.B(n_182),
.Y(n_652)
);

AND2x6_ASAP7_75t_L g653 ( 
.A(n_492),
.B(n_337),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_539),
.B(n_183),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_509),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_550),
.B(n_183),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_514),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_572),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_526),
.B(n_239),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_558),
.B(n_239),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_488),
.B(n_337),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_558),
.B(n_290),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_558),
.B(n_290),
.Y(n_663)
);

NOR2x1p5_ASAP7_75t_L g664 ( 
.A(n_512),
.B(n_176),
.Y(n_664)
);

INVxp33_ASAP7_75t_L g665 ( 
.A(n_490),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_558),
.B(n_294),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_509),
.Y(n_667)
);

NAND3xp33_ASAP7_75t_L g668 ( 
.A(n_549),
.B(n_202),
.C(n_207),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_480),
.A2(n_294),
.B1(n_310),
.B2(n_296),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_562),
.B(n_296),
.Y(n_670)
);

AND2x6_ASAP7_75t_SL g671 ( 
.A(n_570),
.B(n_338),
.Y(n_671)
);

NAND2xp33_ASAP7_75t_SL g672 ( 
.A(n_477),
.B(n_188),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_474),
.B(n_299),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_562),
.B(n_299),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_493),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_541),
.B(n_507),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_514),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_541),
.B(n_301),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_540),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_540),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_498),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_SL g682 ( 
.A1(n_479),
.A2(n_188),
.B1(n_291),
.B2(n_297),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_541),
.B(n_301),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_507),
.B(n_306),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_474),
.B(n_597),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_461),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_598),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_561),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_518),
.B(n_306),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_501),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_510),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_518),
.B(n_307),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_589),
.B(n_511),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_466),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_603),
.B(n_311),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_540),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_474),
.B(n_308),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_597),
.B(n_308),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_509),
.B(n_310),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_524),
.A2(n_230),
.B1(n_259),
.B2(n_288),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_603),
.B(n_311),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_493),
.Y(n_702)
);

AOI22x1_ASAP7_75t_L g703 ( 
.A1(n_596),
.A2(n_343),
.B1(n_342),
.B2(n_338),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_584),
.B(n_343),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_470),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_540),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_582),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_537),
.B(n_342),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_597),
.B(n_259),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_589),
.B(n_208),
.Y(n_710)
);

AOI221xp5_ASAP7_75t_L g711 ( 
.A1(n_591),
.A2(n_291),
.B1(n_297),
.B2(n_309),
.C(n_300),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_547),
.B(n_213),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_464),
.B(n_265),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_464),
.B(n_216),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_598),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_496),
.B(n_267),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_588),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_479),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_565),
.Y(n_719)
);

O2A1O1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_516),
.A2(n_326),
.B(n_319),
.C(n_288),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_588),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_565),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_543),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_496),
.B(n_221),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_504),
.B(n_224),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_530),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_504),
.B(n_523),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_530),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_469),
.A2(n_268),
.B1(n_242),
.B2(n_287),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_532),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_532),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_483),
.B(n_231),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_523),
.A2(n_326),
.B(n_285),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_483),
.B(n_277),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_483),
.B(n_251),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_583),
.B(n_248),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_492),
.B(n_259),
.Y(n_737)
);

OR2x6_ASAP7_75t_L g738 ( 
.A(n_577),
.B(n_288),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_533),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_567),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_533),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_587),
.B(n_64),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_544),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_469),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_483),
.B(n_15),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_524),
.A2(n_77),
.B1(n_153),
.B2(n_151),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_567),
.B(n_16),
.Y(n_747)
);

INVx4_ASAP7_75t_L g748 ( 
.A(n_590),
.Y(n_748)
);

AND2x6_ASAP7_75t_L g749 ( 
.A(n_492),
.B(n_69),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_R g750 ( 
.A(n_512),
.B(n_70),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_492),
.B(n_57),
.Y(n_751)
);

NOR2xp67_ASAP7_75t_L g752 ( 
.A(n_577),
.B(n_535),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_544),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_517),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_584),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_517),
.B(n_79),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_593),
.Y(n_757)
);

INVx8_ASAP7_75t_L g758 ( 
.A(n_584),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_517),
.B(n_46),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_517),
.B(n_84),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_707),
.Y(n_761)
);

BUFx2_ASAP7_75t_L g762 ( 
.A(n_641),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_621),
.B(n_592),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_717),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_621),
.B(n_576),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_658),
.B(n_522),
.Y(n_766)
);

AND2x6_ASAP7_75t_L g767 ( 
.A(n_629),
.B(n_602),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_649),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_646),
.B(n_522),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_721),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_723),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_702),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_641),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_657),
.B(n_584),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_646),
.B(n_528),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_754),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_693),
.B(n_528),
.Y(n_777)
);

INVx1_ASAP7_75t_SL g778 ( 
.A(n_630),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_619),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_757),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_687),
.B(n_527),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_693),
.B(n_560),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_702),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_718),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_677),
.B(n_567),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_625),
.B(n_560),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_710),
.A2(n_524),
.B1(n_568),
.B2(n_538),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_605),
.B(n_527),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_627),
.B(n_497),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_686),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_702),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_688),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_754),
.B(n_491),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_754),
.B(n_491),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_702),
.Y(n_795)
);

INVxp33_ASAP7_75t_L g796 ( 
.A(n_637),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_715),
.B(n_527),
.Y(n_797)
);

OAI22xp33_ASAP7_75t_L g798 ( 
.A1(n_694),
.A2(n_542),
.B1(n_551),
.B2(n_595),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_710),
.B(n_521),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_754),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_627),
.B(n_542),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_704),
.B(n_551),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_695),
.B(n_553),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_617),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_634),
.B(n_545),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_670),
.B(n_482),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_701),
.B(n_585),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_675),
.B(n_586),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_661),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_614),
.B(n_555),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_712),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_713),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_629),
.B(n_491),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_676),
.A2(n_469),
.B1(n_545),
.B2(n_580),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_618),
.A2(n_622),
.B(n_685),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_614),
.B(n_670),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_719),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_722),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_645),
.B(n_595),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_705),
.B(n_564),
.Y(n_820)
);

HB1xp67_ASAP7_75t_L g821 ( 
.A(n_755),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_SL g822 ( 
.A1(n_607),
.A2(n_570),
.B1(n_543),
.B2(n_601),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_655),
.B(n_491),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_750),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_674),
.B(n_554),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_750),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_674),
.B(n_469),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_679),
.B(n_680),
.Y(n_828)
);

NOR3xp33_ASAP7_75t_SL g829 ( 
.A(n_682),
.B(n_608),
.C(n_711),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_671),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_696),
.B(n_706),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_SL g832 ( 
.A1(n_745),
.A2(n_570),
.B1(n_469),
.B2(n_599),
.Y(n_832)
);

NAND2x1p5_ASAP7_75t_L g833 ( 
.A(n_655),
.B(n_491),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_618),
.A2(n_536),
.B(n_590),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_665),
.B(n_566),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_651),
.B(n_469),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_631),
.A2(n_599),
.B1(n_604),
.B2(n_485),
.Y(n_837)
);

AO22x1_ASAP7_75t_L g838 ( 
.A1(n_745),
.A2(n_602),
.B1(n_600),
.B2(n_581),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_681),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_690),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_635),
.B(n_566),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_691),
.B(n_548),
.Y(n_842)
);

AND2x6_ASAP7_75t_SL g843 ( 
.A(n_615),
.B(n_16),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_631),
.A2(n_520),
.B1(n_485),
.B2(n_486),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_664),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_726),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_728),
.Y(n_847)
);

OR2x6_ASAP7_75t_L g848 ( 
.A(n_758),
.B(n_590),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_659),
.B(n_556),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_653),
.B(n_556),
.Y(n_850)
);

NOR2x2_ASAP7_75t_L g851 ( 
.A(n_738),
.B(n_623),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_755),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_730),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_653),
.B(n_557),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_667),
.B(n_594),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_653),
.B(n_557),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_749),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_731),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_667),
.B(n_594),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_653),
.B(n_559),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_739),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_741),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_653),
.B(n_559),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_635),
.B(n_573),
.Y(n_864)
);

NAND3xp33_ASAP7_75t_SL g865 ( 
.A(n_623),
.B(n_729),
.C(n_744),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_751),
.A2(n_571),
.B1(n_581),
.B2(n_579),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_611),
.A2(n_600),
.B(n_515),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_743),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_747),
.Y(n_869)
);

AND2x6_ASAP7_75t_L g870 ( 
.A(n_747),
.B(n_600),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_608),
.B(n_574),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_714),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_678),
.B(n_574),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_632),
.B(n_571),
.Y(n_874)
);

BUFx12f_ASAP7_75t_L g875 ( 
.A(n_738),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_753),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_610),
.B(n_594),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_636),
.B(n_579),
.Y(n_878)
);

NAND3xp33_ASAP7_75t_SL g879 ( 
.A(n_729),
.B(n_471),
.C(n_476),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_708),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_751),
.A2(n_471),
.B1(n_476),
.B2(n_578),
.Y(n_881)
);

CKINVDCx20_ASAP7_75t_R g882 ( 
.A(n_672),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_683),
.B(n_638),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_639),
.B(n_505),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_613),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_740),
.B(n_594),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_736),
.B(n_612),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_732),
.B(n_594),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_642),
.B(n_502),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_620),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_626),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_633),
.A2(n_502),
.B1(n_520),
.B2(n_515),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_675),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_758),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_633),
.A2(n_508),
.B1(n_505),
.B2(n_489),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_644),
.B(n_489),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_R g897 ( 
.A(n_758),
.B(n_590),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_643),
.A2(n_487),
.B(n_486),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_647),
.B(n_487),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_716),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_640),
.Y(n_901)
);

O2A1O1Ixp5_ASAP7_75t_L g902 ( 
.A1(n_643),
.A2(n_484),
.B(n_18),
.C(n_23),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_648),
.B(n_650),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_654),
.A2(n_484),
.B(n_18),
.C(n_24),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_612),
.B(n_17),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_756),
.B(n_91),
.Y(n_906)
);

OR2x2_ASAP7_75t_SL g907 ( 
.A(n_668),
.B(n_17),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_703),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_724),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_727),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_732),
.B(n_24),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_654),
.A2(n_94),
.B1(n_146),
.B2(n_124),
.Y(n_912)
);

OR2x6_ASAP7_75t_SL g913 ( 
.A(n_669),
.B(n_26),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_684),
.B(n_89),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_656),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_689),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_725),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_752),
.B(n_26),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_737),
.B(n_29),
.Y(n_919)
);

INVxp67_ASAP7_75t_SL g920 ( 
.A(n_685),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_734),
.B(n_30),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_737),
.B(n_30),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_738),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_749),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_756),
.B(n_115),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_692),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_749),
.Y(n_927)
);

INVx5_ASAP7_75t_L g928 ( 
.A(n_749),
.Y(n_928)
);

INVx5_ASAP7_75t_L g929 ( 
.A(n_749),
.Y(n_929)
);

AO22x1_ASAP7_75t_L g930 ( 
.A1(n_734),
.A2(n_735),
.B1(n_699),
.B2(n_742),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_759),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_759),
.Y(n_932)
);

OR2x6_ASAP7_75t_L g933 ( 
.A(n_720),
.B(n_31),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_748),
.B(n_118),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_760),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_804),
.Y(n_936)
);

INVx4_ASAP7_75t_L g937 ( 
.A(n_776),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_920),
.A2(n_748),
.B(n_609),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_R g939 ( 
.A(n_824),
.B(n_735),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_816),
.B(n_616),
.Y(n_940)
);

AO22x1_ASAP7_75t_L g941 ( 
.A1(n_905),
.A2(n_700),
.B1(n_760),
.B2(n_746),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_763),
.B(n_616),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_774),
.B(n_709),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_865),
.A2(n_666),
.B1(n_662),
.B2(n_663),
.Y(n_944)
);

OAI21xp33_ASAP7_75t_L g945 ( 
.A1(n_829),
.A2(n_666),
.B(n_662),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_765),
.B(n_660),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_887),
.A2(n_709),
.B(n_660),
.C(n_663),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_778),
.B(n_624),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_776),
.Y(n_949)
);

O2A1O1Ixp5_ASAP7_75t_L g950 ( 
.A1(n_930),
.A2(n_624),
.B(n_628),
.C(n_697),
.Y(n_950)
);

NOR2xp67_ASAP7_75t_L g951 ( 
.A(n_928),
.B(n_698),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_796),
.B(n_697),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_781),
.B(n_673),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_920),
.A2(n_652),
.B(n_628),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_827),
.A2(n_673),
.B(n_606),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_926),
.B(n_733),
.Y(n_956)
);

AND2x2_ASAP7_75t_SL g957 ( 
.A(n_911),
.B(n_34),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_834),
.A2(n_102),
.B(n_119),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_834),
.A2(n_123),
.B(n_157),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_839),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_762),
.Y(n_961)
);

O2A1O1Ixp5_ASAP7_75t_L g962 ( 
.A1(n_799),
.A2(n_887),
.B(n_883),
.C(n_925),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_931),
.A2(n_935),
.B1(n_932),
.B2(n_841),
.Y(n_963)
);

BUFx8_ASAP7_75t_L g964 ( 
.A(n_784),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_SL g965 ( 
.A1(n_882),
.A2(n_822),
.B1(n_900),
.B2(n_806),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_774),
.B(n_785),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_776),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_894),
.B(n_893),
.Y(n_968)
);

OAI21xp33_ASAP7_75t_L g969 ( 
.A1(n_829),
.A2(n_809),
.B(n_779),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_894),
.B(n_789),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_773),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_781),
.B(n_797),
.Y(n_972)
);

INVxp67_ASAP7_75t_L g973 ( 
.A(n_821),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_840),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_865),
.A2(n_922),
.B(n_919),
.C(n_916),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_915),
.B(n_916),
.Y(n_976)
);

NAND2x1p5_ASAP7_75t_L g977 ( 
.A(n_928),
.B(n_929),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_768),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_883),
.A2(n_921),
.B(n_873),
.C(n_871),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_776),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_798),
.B(n_797),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_880),
.B(n_917),
.Y(n_982)
);

BUFx8_ASAP7_75t_SL g983 ( 
.A(n_771),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_910),
.B(n_766),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_871),
.B(n_811),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_815),
.A2(n_903),
.B(n_782),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_869),
.A2(n_798),
.B(n_904),
.C(n_803),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_812),
.B(n_872),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_873),
.B(n_835),
.Y(n_989)
);

AOI22x1_ASAP7_75t_SL g990 ( 
.A1(n_830),
.A2(n_845),
.B1(n_826),
.B2(n_913),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_800),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_772),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_914),
.A2(n_806),
.B(n_805),
.C(n_815),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_800),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_864),
.B(n_825),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_914),
.A2(n_906),
.B(n_925),
.C(n_904),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_807),
.B(n_810),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_906),
.A2(n_787),
.B(n_775),
.C(n_769),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_777),
.A2(n_896),
.B(n_884),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_802),
.B(n_852),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_929),
.A2(n_924),
.B1(n_927),
.B2(n_814),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_761),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_909),
.A2(n_786),
.B(n_878),
.C(n_874),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_820),
.B(n_849),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_832),
.A2(n_912),
.B1(n_764),
.B2(n_770),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_SL g1006 ( 
.A1(n_907),
.A2(n_832),
.B1(n_875),
.B2(n_923),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_772),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_924),
.A2(n_857),
.B1(n_837),
.B2(n_881),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_902),
.A2(n_819),
.B(n_836),
.C(n_780),
.Y(n_1009)
);

BUFx12f_ASAP7_75t_L g1010 ( 
.A(n_843),
.Y(n_1010)
);

OR2x6_ASAP7_75t_L g1011 ( 
.A(n_848),
.B(n_857),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_790),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_792),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_852),
.B(n_801),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_828),
.B(n_831),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_789),
.B(n_808),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_808),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_842),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_889),
.A2(n_899),
.B(n_888),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_870),
.B(n_861),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_897),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_857),
.B(n_800),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_870),
.B(n_862),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_783),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_870),
.B(n_853),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_870),
.B(n_847),
.Y(n_1026)
);

AO22x1_ASAP7_75t_L g1027 ( 
.A1(n_870),
.A2(n_857),
.B1(n_851),
.B2(n_918),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_858),
.B(n_817),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_SL g1029 ( 
.A(n_848),
.B(n_934),
.Y(n_1029)
);

NOR2x1_ASAP7_75t_L g1030 ( 
.A(n_791),
.B(n_795),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_818),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_800),
.B(n_897),
.Y(n_1032)
);

BUFx12f_ASAP7_75t_L g1033 ( 
.A(n_933),
.Y(n_1033)
);

INVx5_ASAP7_75t_L g1034 ( 
.A(n_848),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_846),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_791),
.B(n_795),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_868),
.Y(n_1037)
);

O2A1O1Ixp5_ASAP7_75t_L g1038 ( 
.A1(n_838),
.A2(n_877),
.B(n_908),
.C(n_902),
.Y(n_1038)
);

INVxp67_ASAP7_75t_L g1039 ( 
.A(n_933),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_879),
.A2(n_876),
.B1(n_885),
.B2(n_890),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_891),
.B(n_901),
.Y(n_1041)
);

O2A1O1Ixp5_ASAP7_75t_L g1042 ( 
.A1(n_877),
.A2(n_898),
.B(n_867),
.C(n_856),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_813),
.A2(n_855),
.B(n_823),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_850),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_854),
.B(n_860),
.Y(n_1045)
);

BUFx4f_ASAP7_75t_L g1046 ( 
.A(n_933),
.Y(n_1046)
);

AOI221xp5_ASAP7_75t_L g1047 ( 
.A1(n_879),
.A2(n_881),
.B1(n_866),
.B2(n_886),
.C(n_863),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_813),
.A2(n_823),
.B(n_859),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_767),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_855),
.A2(n_859),
.B(n_793),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_844),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_892),
.A2(n_895),
.B(n_794),
.C(n_767),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_767),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_767),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_934),
.B(n_833),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_833),
.B(n_816),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_894),
.B(n_893),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_905),
.A2(n_816),
.B(n_799),
.C(n_865),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_920),
.A2(n_754),
.B(n_685),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_865),
.A2(n_816),
.B1(n_905),
.B2(n_799),
.Y(n_1060)
);

NAND3xp33_ASAP7_75t_L g1061 ( 
.A(n_829),
.B(n_646),
.C(n_670),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_778),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_816),
.A2(n_887),
.B1(n_865),
.B2(n_710),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_905),
.A2(n_816),
.B(n_799),
.C(n_865),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_804),
.Y(n_1065)
);

CKINVDCx16_ASAP7_75t_R g1066 ( 
.A(n_875),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_920),
.A2(n_816),
.B1(n_932),
.B2(n_931),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_816),
.B(n_621),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1028),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1068),
.B(n_989),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_997),
.B(n_957),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_972),
.B(n_985),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_1059),
.A2(n_938),
.B(n_1043),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_SL g1074 ( 
.A1(n_975),
.A2(n_987),
.B(n_1048),
.Y(n_1074)
);

NOR2xp67_ASAP7_75t_L g1075 ( 
.A(n_1062),
.B(n_971),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_983),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_964),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_1061),
.A2(n_1064),
.B(n_1058),
.C(n_1063),
.Y(n_1078)
);

INVx5_ASAP7_75t_L g1079 ( 
.A(n_949),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_1050),
.A2(n_986),
.B(n_955),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_979),
.A2(n_962),
.B(n_1060),
.C(n_953),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_995),
.B(n_984),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_1042),
.A2(n_954),
.B(n_1019),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_999),
.A2(n_1008),
.B(n_998),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1004),
.A2(n_947),
.B(n_1003),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_1038),
.A2(n_959),
.B(n_958),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_982),
.B(n_976),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_996),
.A2(n_993),
.B(n_1047),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_961),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1018),
.B(n_942),
.Y(n_1090)
);

INVxp67_ASAP7_75t_L g1091 ( 
.A(n_1014),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_956),
.A2(n_963),
.B(n_1009),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_940),
.B(n_946),
.Y(n_1093)
);

AOI221xp5_ASAP7_75t_SL g1094 ( 
.A1(n_981),
.A2(n_969),
.B1(n_945),
.B2(n_1006),
.C(n_1039),
.Y(n_1094)
);

O2A1O1Ixp5_ASAP7_75t_L g1095 ( 
.A1(n_941),
.A2(n_950),
.B(n_1027),
.C(n_1046),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1001),
.A2(n_1067),
.B(n_1045),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_1011),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1052),
.A2(n_943),
.B(n_951),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_1020),
.A2(n_1026),
.B(n_1025),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1060),
.B(n_952),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_948),
.B(n_988),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_1023),
.A2(n_1040),
.B(n_1056),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_939),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1040),
.A2(n_1044),
.B(n_1051),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_1030),
.A2(n_1036),
.B(n_1054),
.Y(n_1105)
);

NAND3x1_ASAP7_75t_L g1106 ( 
.A(n_1016),
.B(n_1015),
.C(n_1065),
.Y(n_1106)
);

OR2x2_ASAP7_75t_L g1107 ( 
.A(n_1000),
.B(n_973),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_944),
.A2(n_1005),
.B(n_1046),
.C(n_951),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1017),
.B(n_970),
.Y(n_1109)
);

AND2x6_ASAP7_75t_L g1110 ( 
.A(n_1049),
.B(n_1053),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_960),
.B(n_974),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1029),
.A2(n_1032),
.B(n_977),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_965),
.A2(n_966),
.B1(n_1033),
.B2(n_1021),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_944),
.A2(n_1005),
.B(n_1002),
.C(n_1035),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_968),
.B(n_1057),
.Y(n_1115)
);

NOR2x1_ASAP7_75t_L g1116 ( 
.A(n_1011),
.B(n_937),
.Y(n_1116)
);

AO31x2_ASAP7_75t_L g1117 ( 
.A1(n_978),
.A2(n_1012),
.A3(n_1013),
.B(n_1037),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1031),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1022),
.A2(n_1055),
.B(n_1011),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_968),
.B(n_1041),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_992),
.B(n_1024),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1066),
.A2(n_990),
.B1(n_1007),
.B2(n_1010),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1034),
.A2(n_991),
.B(n_967),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1034),
.A2(n_949),
.B(n_967),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_SL g1125 ( 
.A1(n_967),
.A2(n_980),
.B(n_994),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_1034),
.Y(n_1126)
);

AO21x1_ASAP7_75t_L g1127 ( 
.A1(n_980),
.A2(n_1064),
.B(n_1058),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_980),
.B(n_994),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_994),
.B(n_1068),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1028),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1068),
.B(n_816),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_986),
.A2(n_754),
.B(n_920),
.Y(n_1132)
);

AO21x2_ASAP7_75t_L g1133 ( 
.A1(n_954),
.A2(n_986),
.B(n_1063),
.Y(n_1133)
);

NAND3x1_ASAP7_75t_L g1134 ( 
.A(n_997),
.B(n_420),
.C(n_788),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_986),
.A2(n_754),
.B(n_920),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_972),
.B(n_658),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1061),
.A2(n_1064),
.B(n_1058),
.C(n_1063),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_972),
.B(n_605),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_986),
.A2(n_754),
.B(n_920),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1068),
.B(n_816),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1068),
.B(n_816),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1061),
.A2(n_605),
.B1(n_317),
.B2(n_788),
.Y(n_1142)
);

CKINVDCx20_ASAP7_75t_R g1143 ( 
.A(n_983),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1040),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1068),
.B(n_816),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1059),
.A2(n_938),
.B(n_815),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_1011),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_949),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1040),
.Y(n_1149)
);

AOI21x1_ASAP7_75t_SL g1150 ( 
.A1(n_942),
.A2(n_816),
.B(n_911),
.Y(n_1150)
);

O2A1O1Ixp5_ASAP7_75t_SL g1151 ( 
.A1(n_981),
.A2(n_737),
.B(n_633),
.C(n_643),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1068),
.B(n_816),
.Y(n_1152)
);

BUFx10_ASAP7_75t_L g1153 ( 
.A(n_1016),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1059),
.A2(n_938),
.B(n_815),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_1011),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_972),
.B(n_658),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_1011),
.Y(n_1157)
);

INVxp67_ASAP7_75t_SL g1158 ( 
.A(n_961),
.Y(n_1158)
);

BUFx2_ASAP7_75t_R g1159 ( 
.A(n_983),
.Y(n_1159)
);

CKINVDCx8_ASAP7_75t_R g1160 ( 
.A(n_1066),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1061),
.A2(n_962),
.B(n_979),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_997),
.B(n_788),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_936),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_947),
.A2(n_998),
.A3(n_1008),
.B(n_996),
.Y(n_1164)
);

NOR4xp25_ASAP7_75t_L g1165 ( 
.A(n_1061),
.B(n_865),
.C(n_1064),
.D(n_1058),
.Y(n_1165)
);

AO31x2_ASAP7_75t_L g1166 ( 
.A1(n_947),
.A2(n_998),
.A3(n_1008),
.B(n_996),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_964),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_972),
.B(n_658),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1068),
.B(n_816),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_947),
.A2(n_998),
.A3(n_1008),
.B(n_996),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_986),
.A2(n_754),
.B(n_920),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1068),
.B(n_816),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_986),
.A2(n_754),
.B(n_920),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_986),
.A2(n_754),
.B(n_920),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_997),
.B(n_788),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1059),
.A2(n_938),
.B(n_815),
.Y(n_1176)
);

CKINVDCx11_ASAP7_75t_R g1177 ( 
.A(n_1010),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_936),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1068),
.B(n_816),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_947),
.A2(n_998),
.A3(n_1008),
.B(n_996),
.Y(n_1180)
);

NAND3xp33_ASAP7_75t_SL g1181 ( 
.A(n_1061),
.B(n_542),
.C(n_512),
.Y(n_1181)
);

OR2x2_ASAP7_75t_L g1182 ( 
.A(n_1068),
.B(n_778),
.Y(n_1182)
);

OAI21xp33_ASAP7_75t_L g1183 ( 
.A1(n_1061),
.A2(n_463),
.B(n_670),
.Y(n_1183)
);

CKINVDCx14_ASAP7_75t_R g1184 ( 
.A(n_939),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_986),
.A2(n_754),
.B(n_920),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_972),
.B(n_658),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1059),
.A2(n_938),
.B(n_815),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_986),
.A2(n_754),
.B(n_920),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1061),
.A2(n_605),
.B1(n_317),
.B2(n_788),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1028),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1061),
.A2(n_962),
.B(n_979),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_972),
.B(n_658),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1040),
.Y(n_1193)
);

AO21x2_ASAP7_75t_L g1194 ( 
.A1(n_954),
.A2(n_986),
.B(n_1063),
.Y(n_1194)
);

INVx2_ASAP7_75t_SL g1195 ( 
.A(n_964),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_SL g1196 ( 
.A1(n_1108),
.A2(n_1081),
.B(n_1078),
.C(n_1137),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_1182),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1132),
.A2(n_1139),
.B(n_1135),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1136),
.A2(n_1186),
.B1(n_1168),
.B2(n_1156),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1097),
.Y(n_1200)
);

OA21x2_ASAP7_75t_L g1201 ( 
.A1(n_1088),
.A2(n_1084),
.B(n_1085),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1092),
.A2(n_1173),
.B(n_1171),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1071),
.B(n_1162),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1174),
.A2(n_1188),
.B(n_1185),
.Y(n_1204)
);

NAND2x1p5_ASAP7_75t_L g1205 ( 
.A(n_1097),
.B(n_1147),
.Y(n_1205)
);

AO21x2_ASAP7_75t_L g1206 ( 
.A1(n_1074),
.A2(n_1191),
.B(n_1161),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1111),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_SL g1208 ( 
.A1(n_1127),
.A2(n_1112),
.B(n_1119),
.Y(n_1208)
);

NAND2x1p5_ASAP7_75t_L g1209 ( 
.A(n_1147),
.B(n_1155),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1069),
.B(n_1130),
.Y(n_1210)
);

AO21x2_ASAP7_75t_L g1211 ( 
.A1(n_1083),
.A2(n_1073),
.B(n_1096),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1146),
.A2(n_1154),
.B(n_1176),
.Y(n_1212)
);

CKINVDCx6p67_ASAP7_75t_R g1213 ( 
.A(n_1143),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1133),
.A2(n_1194),
.B(n_1080),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1093),
.B(n_1072),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1115),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1070),
.B(n_1100),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1165),
.A2(n_1151),
.B(n_1114),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1098),
.A2(n_1095),
.B(n_1104),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1192),
.A2(n_1189),
.B1(n_1142),
.B2(n_1138),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1187),
.A2(n_1105),
.B(n_1086),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1099),
.A2(n_1150),
.B(n_1102),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1082),
.B(n_1090),
.Y(n_1223)
);

AOI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1181),
.A2(n_1175),
.B1(n_1183),
.B2(n_1106),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1190),
.B(n_1107),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1163),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1144),
.A2(n_1149),
.B(n_1193),
.Y(n_1227)
);

AO31x2_ASAP7_75t_L g1228 ( 
.A1(n_1193),
.A2(n_1180),
.A3(n_1164),
.B(n_1166),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1155),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1131),
.A2(n_1172),
.B1(n_1140),
.B2(n_1141),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1157),
.A2(n_1121),
.B(n_1124),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1115),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1123),
.A2(n_1116),
.B(n_1126),
.Y(n_1233)
);

OA21x2_ASAP7_75t_L g1234 ( 
.A1(n_1094),
.A2(n_1129),
.B(n_1178),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_1079),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1091),
.B(n_1101),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1117),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1117),
.Y(n_1238)
);

NOR2xp67_ASAP7_75t_L g1239 ( 
.A(n_1103),
.B(n_1089),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1117),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1118),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1087),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_1158),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1145),
.A2(n_1179),
.B1(n_1169),
.B2(n_1152),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1128),
.Y(n_1245)
);

OR2x6_ASAP7_75t_L g1246 ( 
.A(n_1126),
.B(n_1125),
.Y(n_1246)
);

NOR2xp67_ASAP7_75t_SL g1247 ( 
.A(n_1160),
.B(n_1076),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1166),
.A2(n_1180),
.B(n_1170),
.C(n_1113),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1109),
.B(n_1120),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1134),
.A2(n_1079),
.B1(n_1184),
.B2(n_1122),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1153),
.B(n_1075),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1110),
.A2(n_1079),
.B(n_1195),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1110),
.A2(n_1167),
.B(n_1077),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1110),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_1177),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1148),
.B(n_1159),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1088),
.A2(n_1061),
.B(n_1063),
.Y(n_1257)
);

AO31x2_ASAP7_75t_L g1258 ( 
.A1(n_1081),
.A2(n_1084),
.A3(n_1088),
.B(n_1127),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1088),
.A2(n_1084),
.B(n_1085),
.Y(n_1259)
);

AO31x2_ASAP7_75t_L g1260 ( 
.A1(n_1081),
.A2(n_1084),
.A3(n_1088),
.B(n_1127),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_R g1261 ( 
.A(n_1184),
.B(n_771),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1111),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1088),
.A2(n_865),
.B(n_1061),
.C(n_979),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1071),
.B(n_1162),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1111),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1132),
.A2(n_1139),
.B(n_1135),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1111),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_1143),
.Y(n_1268)
);

CKINVDCx11_ASAP7_75t_R g1269 ( 
.A(n_1160),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1088),
.A2(n_1084),
.B(n_1085),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1088),
.A2(n_1061),
.B(n_1063),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_SL g1272 ( 
.A1(n_1088),
.A2(n_957),
.B1(n_570),
.B2(n_1061),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1093),
.B(n_1072),
.Y(n_1273)
);

AO31x2_ASAP7_75t_L g1274 ( 
.A1(n_1081),
.A2(n_1084),
.A3(n_1088),
.B(n_1127),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1093),
.B(n_1072),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1132),
.A2(n_1139),
.B(n_1135),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1182),
.B(n_1069),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1132),
.A2(n_1139),
.B(n_1135),
.Y(n_1278)
);

CKINVDCx11_ASAP7_75t_R g1279 ( 
.A(n_1160),
.Y(n_1279)
);

INVx6_ASAP7_75t_L g1280 ( 
.A(n_1079),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1088),
.A2(n_1084),
.B(n_1085),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1088),
.A2(n_1061),
.B(n_1063),
.Y(n_1282)
);

AOI21xp33_ASAP7_75t_SL g1283 ( 
.A1(n_1136),
.A2(n_542),
.B(n_512),
.Y(n_1283)
);

BUFx10_ASAP7_75t_L g1284 ( 
.A(n_1076),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1132),
.A2(n_1139),
.B(n_1135),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1111),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1088),
.A2(n_1061),
.B(n_1063),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_1182),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1100),
.A2(n_865),
.B1(n_1061),
.B2(n_957),
.Y(n_1289)
);

INVx3_ASAP7_75t_SL g1290 ( 
.A(n_1103),
.Y(n_1290)
);

AOI21xp33_ASAP7_75t_L g1291 ( 
.A1(n_1100),
.A2(n_1064),
.B(n_1058),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1132),
.A2(n_1139),
.B(n_1135),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1132),
.A2(n_1139),
.B(n_1135),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1235),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1217),
.B(n_1215),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1199),
.A2(n_1272),
.B1(n_1289),
.B2(n_1220),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1197),
.B(n_1288),
.Y(n_1297)
);

O2A1O1Ixp5_ASAP7_75t_L g1298 ( 
.A1(n_1218),
.A2(n_1259),
.B(n_1271),
.C(n_1282),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1225),
.B(n_1277),
.Y(n_1299)
);

AOI211xp5_ASAP7_75t_L g1300 ( 
.A1(n_1196),
.A2(n_1287),
.B(n_1271),
.C(n_1282),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1203),
.B(n_1264),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1261),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1272),
.A2(n_1289),
.B1(n_1275),
.B2(n_1273),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1210),
.B(n_1243),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1230),
.A2(n_1244),
.B1(n_1223),
.B2(n_1242),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1256),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_1216),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_1226),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1248),
.B(n_1245),
.Y(n_1309)
);

OAI31xp33_ASAP7_75t_L g1310 ( 
.A1(n_1263),
.A2(n_1291),
.A3(n_1244),
.B(n_1230),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1248),
.B(n_1257),
.Y(n_1311)
);

CKINVDCx14_ASAP7_75t_R g1312 ( 
.A(n_1261),
.Y(n_1312)
);

AOI221xp5_ASAP7_75t_L g1313 ( 
.A1(n_1291),
.A2(n_1287),
.B1(n_1257),
.B2(n_1263),
.C(n_1218),
.Y(n_1313)
);

AOI211xp5_ASAP7_75t_L g1314 ( 
.A1(n_1283),
.A2(n_1250),
.B(n_1224),
.C(n_1219),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1250),
.A2(n_1208),
.B(n_1219),
.C(n_1265),
.Y(n_1315)
);

INVxp67_ASAP7_75t_L g1316 ( 
.A(n_1251),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_SL g1317 ( 
.A1(n_1235),
.A2(n_1270),
.B(n_1281),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1249),
.B(n_1232),
.Y(n_1318)
);

AND2x6_ASAP7_75t_L g1319 ( 
.A(n_1254),
.B(n_1235),
.Y(n_1319)
);

INVx3_ASAP7_75t_SL g1320 ( 
.A(n_1290),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_SL g1321 ( 
.A1(n_1255),
.A2(n_1251),
.B1(n_1290),
.B2(n_1268),
.Y(n_1321)
);

NAND3xp33_ASAP7_75t_L g1322 ( 
.A(n_1201),
.B(n_1281),
.C(n_1270),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1207),
.A2(n_1267),
.B1(n_1262),
.B2(n_1286),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1206),
.B(n_1258),
.Y(n_1324)
);

O2A1O1Ixp5_ASAP7_75t_L g1325 ( 
.A1(n_1253),
.A2(n_1202),
.B(n_1214),
.C(n_1252),
.Y(n_1325)
);

BUFx4f_ASAP7_75t_L g1326 ( 
.A(n_1213),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_SL g1327 ( 
.A1(n_1235),
.A2(n_1246),
.B(n_1252),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1241),
.B(n_1234),
.Y(n_1328)
);

OAI22x1_ASAP7_75t_L g1329 ( 
.A1(n_1234),
.A2(n_1209),
.B1(n_1205),
.B2(n_1229),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1228),
.B(n_1260),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1205),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_SL g1332 ( 
.A1(n_1246),
.A2(n_1239),
.B(n_1209),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1269),
.B(n_1279),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1233),
.B(n_1231),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1237),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_SL g1336 ( 
.A1(n_1280),
.A2(n_1240),
.B(n_1238),
.Y(n_1336)
);

INVx2_ASAP7_75t_SL g1337 ( 
.A(n_1284),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1269),
.B(n_1279),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1274),
.B(n_1280),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1274),
.B(n_1280),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_1284),
.Y(n_1341)
);

O2A1O1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1211),
.A2(n_1274),
.B(n_1247),
.C(n_1222),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1221),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1198),
.A2(n_1204),
.B1(n_1293),
.B2(n_1266),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1276),
.B(n_1292),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1278),
.B(n_1285),
.Y(n_1346)
);

O2A1O1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1212),
.A2(n_981),
.B(n_1061),
.C(n_979),
.Y(n_1347)
);

NAND2x1p5_ASAP7_75t_L g1348 ( 
.A(n_1227),
.B(n_1243),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1252),
.B(n_1200),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1199),
.A2(n_1272),
.B1(n_957),
.B2(n_1289),
.Y(n_1350)
);

OA21x2_ASAP7_75t_L g1351 ( 
.A1(n_1219),
.A2(n_1218),
.B(n_1214),
.Y(n_1351)
);

OA21x2_ASAP7_75t_L g1352 ( 
.A1(n_1219),
.A2(n_1218),
.B(n_1214),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1235),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1203),
.B(n_1264),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1197),
.B(n_1288),
.Y(n_1355)
);

INVx5_ASAP7_75t_L g1356 ( 
.A(n_1246),
.Y(n_1356)
);

INVxp67_ASAP7_75t_L g1357 ( 
.A(n_1236),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_SL g1358 ( 
.A1(n_1223),
.A2(n_865),
.B(n_979),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1243),
.Y(n_1359)
);

O2A1O1Ixp5_ASAP7_75t_L g1360 ( 
.A1(n_1218),
.A2(n_1088),
.B(n_941),
.C(n_1259),
.Y(n_1360)
);

AOI221x1_ASAP7_75t_SL g1361 ( 
.A1(n_1215),
.A2(n_608),
.B1(n_1061),
.B2(n_1156),
.C(n_1136),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_1235),
.Y(n_1362)
);

OA21x2_ASAP7_75t_L g1363 ( 
.A1(n_1219),
.A2(n_1218),
.B(n_1214),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1335),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1334),
.B(n_1345),
.Y(n_1365)
);

BUFx6f_ASAP7_75t_L g1366 ( 
.A(n_1345),
.Y(n_1366)
);

AOI21xp33_ASAP7_75t_L g1367 ( 
.A1(n_1296),
.A2(n_1310),
.B(n_1300),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1343),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1324),
.B(n_1330),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1322),
.A2(n_1298),
.B(n_1360),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1349),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1351),
.B(n_1352),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1328),
.Y(n_1373)
);

BUFx4f_ASAP7_75t_SL g1374 ( 
.A(n_1320),
.Y(n_1374)
);

BUFx2_ASAP7_75t_L g1375 ( 
.A(n_1348),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1305),
.B(n_1313),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1325),
.A2(n_1344),
.B(n_1346),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1329),
.Y(n_1378)
);

AO21x1_ASAP7_75t_SL g1379 ( 
.A1(n_1311),
.A2(n_1309),
.B(n_1295),
.Y(n_1379)
);

OR2x6_ASAP7_75t_L g1380 ( 
.A(n_1317),
.B(n_1336),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1363),
.B(n_1339),
.Y(n_1381)
);

BUFx12f_ASAP7_75t_L g1382 ( 
.A(n_1341),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1359),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1363),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1340),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1308),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1342),
.Y(n_1387)
);

INVx2_ASAP7_75t_SL g1388 ( 
.A(n_1356),
.Y(n_1388)
);

AO21x2_ASAP7_75t_L g1389 ( 
.A1(n_1296),
.A2(n_1358),
.B(n_1315),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1300),
.B(n_1310),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1301),
.B(n_1354),
.Y(n_1391)
);

BUFx4f_ASAP7_75t_SL g1392 ( 
.A(n_1306),
.Y(n_1392)
);

AO21x2_ASAP7_75t_L g1393 ( 
.A1(n_1347),
.A2(n_1350),
.B(n_1305),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1323),
.Y(n_1394)
);

AO21x2_ASAP7_75t_L g1395 ( 
.A1(n_1350),
.A2(n_1303),
.B(n_1323),
.Y(n_1395)
);

INVxp67_ASAP7_75t_L g1396 ( 
.A(n_1304),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1319),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1319),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1368),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1375),
.Y(n_1400)
);

AOI211xp5_ASAP7_75t_SL g1401 ( 
.A1(n_1367),
.A2(n_1314),
.B(n_1327),
.C(n_1332),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1369),
.B(n_1299),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1397),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1364),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1381),
.B(n_1357),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1386),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1381),
.B(n_1318),
.Y(n_1407)
);

OR2x2_ASAP7_75t_SL g1408 ( 
.A(n_1376),
.B(n_1331),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1365),
.B(n_1319),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1381),
.B(n_1314),
.Y(n_1410)
);

INVxp67_ASAP7_75t_L g1411 ( 
.A(n_1379),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1385),
.B(n_1316),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1386),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1385),
.B(n_1355),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1367),
.A2(n_1297),
.B1(n_1361),
.B2(n_1307),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1373),
.B(n_1361),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_1366),
.Y(n_1417)
);

NAND2x1_ASAP7_75t_L g1418 ( 
.A(n_1380),
.B(n_1353),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1404),
.Y(n_1419)
);

INVxp67_ASAP7_75t_SL g1420 ( 
.A(n_1406),
.Y(n_1420)
);

NAND2x1p5_ASAP7_75t_L g1421 ( 
.A(n_1418),
.B(n_1388),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1410),
.A2(n_1390),
.B1(n_1389),
.B2(n_1395),
.Y(n_1422)
);

AO21x2_ASAP7_75t_L g1423 ( 
.A1(n_1416),
.A2(n_1384),
.B(n_1372),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1410),
.A2(n_1390),
.B1(n_1389),
.B2(n_1395),
.Y(n_1424)
);

NAND4xp25_ASAP7_75t_L g1425 ( 
.A(n_1415),
.B(n_1390),
.C(n_1376),
.D(n_1338),
.Y(n_1425)
);

INVxp67_ASAP7_75t_L g1426 ( 
.A(n_1402),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1404),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1399),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1404),
.Y(n_1429)
);

AO21x2_ASAP7_75t_L g1430 ( 
.A1(n_1416),
.A2(n_1384),
.B(n_1372),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1410),
.B(n_1341),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1415),
.A2(n_1398),
.B1(n_1397),
.B2(n_1396),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1411),
.A2(n_1389),
.B1(n_1395),
.B2(n_1393),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1403),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1402),
.B(n_1337),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1411),
.A2(n_1389),
.B1(n_1395),
.B2(n_1393),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1417),
.Y(n_1437)
);

OAI221xp5_ASAP7_75t_L g1438 ( 
.A1(n_1401),
.A2(n_1396),
.B1(n_1378),
.B2(n_1387),
.C(n_1333),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1408),
.A2(n_1398),
.B1(n_1392),
.B2(n_1394),
.Y(n_1439)
);

INVxp67_ASAP7_75t_L g1440 ( 
.A(n_1402),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1405),
.B(n_1371),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1406),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1405),
.B(n_1371),
.Y(n_1443)
);

OAI21xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1401),
.A2(n_1312),
.B(n_1341),
.Y(n_1444)
);

NAND3xp33_ASAP7_75t_L g1445 ( 
.A(n_1413),
.B(n_1387),
.C(n_1370),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1403),
.Y(n_1446)
);

OA21x2_ASAP7_75t_L g1447 ( 
.A1(n_1399),
.A2(n_1377),
.B(n_1384),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1408),
.A2(n_1398),
.B1(n_1392),
.B2(n_1394),
.Y(n_1448)
);

BUFx3_ASAP7_75t_L g1449 ( 
.A(n_1403),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1413),
.B(n_1383),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1400),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1412),
.B(n_1414),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1405),
.B(n_1371),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_SL g1454 ( 
.A(n_1409),
.B(n_1374),
.Y(n_1454)
);

INVx4_ASAP7_75t_SL g1455 ( 
.A(n_1434),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1419),
.Y(n_1456)
);

INVx4_ASAP7_75t_SL g1457 ( 
.A(n_1434),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1450),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1426),
.B(n_1412),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1440),
.B(n_1412),
.Y(n_1460)
);

INVx5_ASAP7_75t_L g1461 ( 
.A(n_1437),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1442),
.Y(n_1462)
);

CKINVDCx16_ASAP7_75t_R g1463 ( 
.A(n_1434),
.Y(n_1463)
);

INVxp67_ASAP7_75t_SL g1464 ( 
.A(n_1450),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1441),
.B(n_1407),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1421),
.A2(n_1418),
.B(n_1437),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1441),
.B(n_1407),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1419),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1447),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1427),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1427),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1429),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1428),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1435),
.B(n_1414),
.Y(n_1474)
);

INVx1_ASAP7_75t_SL g1475 ( 
.A(n_1431),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1428),
.Y(n_1476)
);

INVx4_ASAP7_75t_SL g1477 ( 
.A(n_1446),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1423),
.B(n_1408),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_1446),
.Y(n_1479)
);

BUFx2_ASAP7_75t_L g1480 ( 
.A(n_1421),
.Y(n_1480)
);

OR2x6_ASAP7_75t_L g1481 ( 
.A(n_1445),
.B(n_1380),
.Y(n_1481)
);

INVx4_ASAP7_75t_SL g1482 ( 
.A(n_1446),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1429),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1443),
.B(n_1407),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1449),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1475),
.B(n_1374),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1458),
.B(n_1422),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1464),
.B(n_1424),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1455),
.B(n_1443),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1462),
.Y(n_1490)
);

NOR2x1_ASAP7_75t_L g1491 ( 
.A(n_1485),
.B(n_1444),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1474),
.B(n_1438),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1459),
.B(n_1460),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1473),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1455),
.B(n_1453),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1478),
.B(n_1423),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1455),
.B(n_1454),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1456),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1456),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1478),
.B(n_1423),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1465),
.B(n_1453),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1463),
.Y(n_1502)
);

NOR2xp67_ASAP7_75t_L g1503 ( 
.A(n_1461),
.B(n_1439),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1468),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1468),
.Y(n_1505)
);

INVx4_ASAP7_75t_L g1506 ( 
.A(n_1455),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1470),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1455),
.B(n_1449),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1467),
.B(n_1484),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1470),
.B(n_1423),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1471),
.B(n_1430),
.Y(n_1511)
);

INVxp67_ASAP7_75t_L g1512 ( 
.A(n_1485),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1457),
.B(n_1449),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1457),
.B(n_1437),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1473),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1471),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1476),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1472),
.B(n_1430),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1472),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1479),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1463),
.B(n_1302),
.Y(n_1521)
);

NAND3xp33_ASAP7_75t_L g1522 ( 
.A(n_1481),
.B(n_1433),
.C(n_1436),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1467),
.B(n_1383),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1457),
.B(n_1477),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1483),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1457),
.B(n_1451),
.Y(n_1526)
);

INVxp67_ASAP7_75t_L g1527 ( 
.A(n_1485),
.Y(n_1527)
);

O2A1O1Ixp33_ASAP7_75t_SL g1528 ( 
.A1(n_1502),
.A2(n_1444),
.B(n_1439),
.C(n_1448),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1524),
.B(n_1457),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1498),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1498),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1487),
.B(n_1452),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1510),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1524),
.B(n_1477),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1499),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1497),
.B(n_1477),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1490),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1509),
.B(n_1430),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1492),
.B(n_1484),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1499),
.Y(n_1540)
);

INVxp33_ASAP7_75t_L g1541 ( 
.A(n_1491),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1493),
.B(n_1430),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1504),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1512),
.B(n_1479),
.Y(n_1544)
);

OR2x6_ASAP7_75t_L g1545 ( 
.A(n_1506),
.B(n_1497),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1510),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1506),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1505),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_SL g1549 ( 
.A(n_1497),
.B(n_1477),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1527),
.B(n_1488),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1523),
.B(n_1483),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1507),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1520),
.B(n_1391),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1486),
.B(n_1391),
.Y(n_1554)
);

INVxp67_ASAP7_75t_SL g1555 ( 
.A(n_1503),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1511),
.Y(n_1556)
);

NAND2x1p5_ASAP7_75t_L g1557 ( 
.A(n_1506),
.B(n_1480),
.Y(n_1557)
);

NOR2x1p5_ASAP7_75t_SL g1558 ( 
.A(n_1496),
.B(n_1469),
.Y(n_1558)
);

INVx1_ASAP7_75t_SL g1559 ( 
.A(n_1508),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1516),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1522),
.A2(n_1425),
.B(n_1481),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1519),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1525),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1537),
.B(n_1496),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1529),
.B(n_1508),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1557),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1557),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1547),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1530),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1541),
.B(n_1513),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1541),
.B(n_1513),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1531),
.Y(n_1572)
);

CKINVDCx16_ASAP7_75t_R g1573 ( 
.A(n_1545),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1545),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1559),
.B(n_1521),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1535),
.Y(n_1576)
);

AND3x1_ASAP7_75t_L g1577 ( 
.A(n_1529),
.B(n_1534),
.C(n_1561),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1554),
.B(n_1321),
.Y(n_1578)
);

NOR2x1_ASAP7_75t_L g1579 ( 
.A(n_1545),
.B(n_1526),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1532),
.B(n_1500),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1540),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1539),
.B(n_1477),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1534),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1536),
.B(n_1526),
.Y(n_1584)
);

BUFx3_ASAP7_75t_L g1585 ( 
.A(n_1545),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1543),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1536),
.B(n_1489),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1550),
.B(n_1501),
.Y(n_1588)
);

OAI21xp33_ASAP7_75t_L g1589 ( 
.A1(n_1583),
.A2(n_1544),
.B(n_1549),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1577),
.A2(n_1549),
.B1(n_1528),
.B2(n_1555),
.Y(n_1590)
);

O2A1O1Ixp33_ASAP7_75t_L g1591 ( 
.A1(n_1570),
.A2(n_1528),
.B(n_1481),
.C(n_1560),
.Y(n_1591)
);

OAI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1575),
.A2(n_1425),
.B1(n_1481),
.B2(n_1562),
.C(n_1548),
.Y(n_1592)
);

AO21x1_ASAP7_75t_L g1593 ( 
.A1(n_1574),
.A2(n_1500),
.B(n_1552),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1569),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1573),
.A2(n_1579),
.B1(n_1481),
.B2(n_1571),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1569),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1568),
.B(n_1563),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1572),
.Y(n_1598)
);

AOI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1565),
.A2(n_1389),
.B1(n_1489),
.B2(n_1495),
.Y(n_1599)
);

AOI31xp33_ASAP7_75t_L g1600 ( 
.A1(n_1579),
.A2(n_1514),
.A3(n_1448),
.B(n_1495),
.Y(n_1600)
);

AOI21xp33_ASAP7_75t_L g1601 ( 
.A1(n_1585),
.A2(n_1542),
.B(n_1551),
.Y(n_1601)
);

AOI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1568),
.A2(n_1542),
.B1(n_1432),
.B2(n_1538),
.C(n_1533),
.Y(n_1602)
);

INVxp67_ASAP7_75t_SL g1603 ( 
.A(n_1565),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1574),
.B(n_1553),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1585),
.B(n_1482),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1572),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_SL g1607 ( 
.A1(n_1573),
.A2(n_1389),
.B1(n_1432),
.B2(n_1395),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1603),
.B(n_1584),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1605),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1593),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1589),
.B(n_1584),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1597),
.B(n_1578),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1590),
.B(n_1587),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1604),
.B(n_1587),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1607),
.A2(n_1582),
.B1(n_1395),
.B2(n_1588),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1605),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1595),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1592),
.B(n_1566),
.Y(n_1618)
);

AOI211xp5_ASAP7_75t_L g1619 ( 
.A1(n_1610),
.A2(n_1591),
.B(n_1602),
.C(n_1601),
.Y(n_1619)
);

NOR2xp67_ASAP7_75t_L g1620 ( 
.A(n_1610),
.B(n_1566),
.Y(n_1620)
);

NOR3xp33_ASAP7_75t_L g1621 ( 
.A(n_1617),
.B(n_1600),
.C(n_1596),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1613),
.A2(n_1611),
.B(n_1612),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1614),
.A2(n_1567),
.B(n_1594),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1608),
.Y(n_1624)
);

AOI211xp5_ASAP7_75t_L g1625 ( 
.A1(n_1618),
.A2(n_1567),
.B(n_1606),
.C(n_1598),
.Y(n_1625)
);

AOI222xp33_ASAP7_75t_L g1626 ( 
.A1(n_1615),
.A2(n_1558),
.B1(n_1586),
.B2(n_1576),
.C1(n_1581),
.C2(n_1556),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1609),
.B(n_1580),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1616),
.B(n_1586),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1624),
.B(n_1599),
.Y(n_1629)
);

OAI211xp5_ASAP7_75t_SL g1630 ( 
.A1(n_1619),
.A2(n_1581),
.B(n_1576),
.C(n_1564),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1627),
.Y(n_1631)
);

NOR2x1_ASAP7_75t_L g1632 ( 
.A(n_1620),
.B(n_1564),
.Y(n_1632)
);

A2O1A1Ixp33_ASAP7_75t_L g1633 ( 
.A1(n_1622),
.A2(n_1580),
.B(n_1514),
.C(n_1538),
.Y(n_1633)
);

OAI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1621),
.A2(n_1623),
.B(n_1626),
.Y(n_1634)
);

INVxp67_ASAP7_75t_L g1635 ( 
.A(n_1632),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1631),
.B(n_1625),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1629),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1634),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1630),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1633),
.B(n_1628),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1631),
.B(n_1551),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1635),
.B(n_1533),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1641),
.B(n_1546),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1638),
.A2(n_1482),
.B1(n_1546),
.B2(n_1556),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1636),
.A2(n_1326),
.B(n_1494),
.Y(n_1645)
);

AOI221xp5_ASAP7_75t_L g1646 ( 
.A1(n_1639),
.A2(n_1480),
.B1(n_1517),
.B2(n_1515),
.C(n_1494),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1645),
.B(n_1637),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1643),
.B(n_1636),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1644),
.A2(n_1640),
.B1(n_1482),
.B2(n_1382),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1647),
.Y(n_1650)
);

AOI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1650),
.A2(n_1648),
.B1(n_1649),
.B2(n_1646),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1651),
.Y(n_1652)
);

OAI22x1_ASAP7_75t_L g1653 ( 
.A1(n_1651),
.A2(n_1642),
.B1(n_1461),
.B2(n_1515),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1652),
.A2(n_1326),
.B(n_1517),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1653),
.A2(n_1482),
.B1(n_1382),
.B2(n_1461),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1654),
.B(n_1511),
.Y(n_1656)
);

INVxp33_ASAP7_75t_L g1657 ( 
.A(n_1655),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1657),
.B(n_1461),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1658),
.A2(n_1656),
.B(n_1518),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1659),
.B(n_1518),
.Y(n_1660)
);

INVxp67_ASAP7_75t_L g1661 ( 
.A(n_1660),
.Y(n_1661)
);

AOI31xp33_ASAP7_75t_L g1662 ( 
.A1(n_1661),
.A2(n_1382),
.A3(n_1420),
.B(n_1388),
.Y(n_1662)
);

AOI211xp5_ASAP7_75t_L g1663 ( 
.A1(n_1662),
.A2(n_1294),
.B(n_1362),
.C(n_1466),
.Y(n_1663)
);


endmodule