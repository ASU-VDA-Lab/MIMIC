module fake_jpeg_26355_n_47 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_47);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_47;

wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_7),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_30),
.B(n_29),
.Y(n_34)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_3),
.B1(n_5),
.B2(n_10),
.Y(n_32)
);

AOI22x1_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_37)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_27),
.B(n_16),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_27),
.Y(n_41)
);

OR2x2_ASAP7_75t_SL g35 ( 
.A(n_30),
.B(n_23),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_37),
.B(n_38),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_41),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_43),
.B(n_15),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_17),
.B(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_19),
.Y(n_46)
);

AOI32xp33_ASAP7_75t_SL g47 ( 
.A1(n_46),
.A2(n_20),
.A3(n_21),
.B1(n_40),
.B2(n_36),
.Y(n_47)
);


endmodule