module fake_jpeg_11332_n_283 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_283);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_283;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_41),
.Y(n_79)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_44),
.Y(n_91)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_8),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_50),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_0),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

NAND2x1_ASAP7_75t_SL g55 ( 
.A(n_24),
.B(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_19),
.Y(n_70)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_17),
.B(n_7),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_23),
.B(n_7),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_40),
.B1(n_29),
.B2(n_37),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_67),
.A2(n_76),
.B1(n_100),
.B2(n_105),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_48),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_22),
.B1(n_33),
.B2(n_32),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_88),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_32),
.B1(n_62),
.B2(n_59),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_40),
.B1(n_29),
.B2(n_34),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_62),
.B1(n_44),
.B2(n_64),
.Y(n_78)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_28),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_90),
.Y(n_129)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_46),
.A2(n_34),
.B1(n_37),
.B2(n_54),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_30),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_46),
.A2(n_23),
.B1(n_30),
.B2(n_28),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_95),
.B1(n_97),
.B2(n_3),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_51),
.A2(n_27),
.B1(n_21),
.B2(n_20),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_21),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_48),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_51),
.A2(n_18),
.B1(n_35),
.B2(n_19),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_47),
.A2(n_18),
.B1(n_35),
.B2(n_36),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_35),
.B1(n_36),
.B2(n_2),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_41),
.B(n_35),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_102),
.B(n_103),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_45),
.B(n_9),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_47),
.A2(n_36),
.B1(n_0),
.B2(n_2),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_48),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_106),
.A2(n_4),
.B1(n_9),
.B2(n_11),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_110),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_65),
.A2(n_54),
.B1(n_56),
.B2(n_43),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_109),
.A2(n_132),
.B1(n_140),
.B2(n_122),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_1),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_136),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_79),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

AO221x1_ASAP7_75t_L g165 ( 
.A1(n_113),
.A2(n_124),
.B1(n_83),
.B2(n_98),
.C(n_119),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_66),
.B(n_58),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_114),
.B(n_128),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_116),
.B(n_115),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_117),
.A2(n_127),
.B(n_133),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_71),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_70),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_13),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_65),
.B(n_13),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_130),
.B(n_137),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_87),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_80),
.A2(n_91),
.B1(n_82),
.B2(n_84),
.Y(n_133)
);

AO22x1_ASAP7_75t_SL g134 ( 
.A1(n_68),
.A2(n_15),
.B1(n_85),
.B2(n_97),
.Y(n_134)
);

AO22x1_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_89),
.B1(n_72),
.B2(n_107),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_68),
.B(n_92),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_72),
.B(n_69),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_73),
.B(n_79),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_139),
.B(n_89),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_82),
.A2(n_84),
.B1(n_69),
.B2(n_104),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_91),
.A2(n_98),
.B1(n_104),
.B2(n_94),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_91),
.B1(n_79),
.B2(n_71),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_145),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_113),
.B1(n_126),
.B2(n_131),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_150),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_155),
.A2(n_124),
.B(n_134),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_157),
.B(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_108),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_160),
.B(n_166),
.Y(n_201)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

FAx1_ASAP7_75t_SL g164 ( 
.A(n_111),
.B(n_107),
.CI(n_73),
.CON(n_164),
.SN(n_164)
);

NOR3xp33_ASAP7_75t_SL g200 ( 
.A(n_164),
.B(n_154),
.C(n_149),
.Y(n_200)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_129),
.B(n_83),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_108),
.B(n_110),
.C(n_135),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_127),
.Y(n_174)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_141),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_171),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_129),
.B1(n_173),
.B2(n_161),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_173),
.A2(n_134),
.B1(n_116),
.B2(n_115),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_192),
.C(n_196),
.Y(n_204)
);

HAxp5_ASAP7_75t_SL g176 ( 
.A(n_164),
.B(n_146),
.CON(n_176),
.SN(n_176)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_176),
.A2(n_184),
.B1(n_182),
.B2(n_197),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_177),
.A2(n_144),
.B1(n_155),
.B2(n_147),
.Y(n_202)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_180),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_182),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_112),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_183),
.A2(n_187),
.B1(n_191),
.B2(n_143),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_117),
.B1(n_138),
.B2(n_134),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_123),
.B(n_121),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_194),
.B1(n_195),
.B2(n_197),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_172),
.A2(n_138),
.B1(n_126),
.B2(n_131),
.Y(n_191)
);

OR2x6_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_146),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_146),
.A2(n_167),
.B(n_155),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_181),
.Y(n_222)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_200),
.B(n_156),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_220),
.B1(n_179),
.B2(n_185),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_142),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_203),
.B(n_207),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_206),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_222),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_162),
.C(n_169),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_201),
.B(n_152),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_221),
.Y(n_227)
);

AOI322xp5_ASAP7_75t_SL g211 ( 
.A1(n_200),
.A2(n_144),
.A3(n_152),
.B1(n_163),
.B2(n_150),
.C1(n_148),
.C2(n_168),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_211),
.B(n_214),
.Y(n_238)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_195),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_168),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_186),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_217),
.Y(n_235)
);

A2O1A1O1Ixp25_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_223),
.B(n_195),
.C(n_190),
.D(n_185),
.Y(n_228)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_188),
.A2(n_143),
.B1(n_151),
.B2(n_156),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_151),
.C(n_176),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_191),
.C(n_189),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_208),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_239),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_195),
.B(n_190),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_225),
.A2(n_228),
.B(n_205),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_229),
.A2(n_233),
.B1(n_225),
.B2(n_226),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_219),
.B1(n_215),
.B2(n_209),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_179),
.Y(n_231)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_231),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_198),
.B1(n_199),
.B2(n_193),
.Y(n_233)
);

AO21x1_ASAP7_75t_L g234 ( 
.A1(n_205),
.A2(n_193),
.B(n_180),
.Y(n_234)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

AOI322xp5_ASAP7_75t_L g241 ( 
.A1(n_238),
.A2(n_205),
.A3(n_210),
.B1(n_204),
.B2(n_221),
.C1(n_206),
.C2(n_222),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_251),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_232),
.B(n_228),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_248),
.B1(n_239),
.B2(n_244),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_216),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_250),
.C(n_252),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_216),
.B1(n_233),
.B2(n_231),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_216),
.Y(n_249)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_249),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_227),
.C(n_232),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_232),
.C(n_229),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_240),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_255),
.A2(n_258),
.B1(n_259),
.B2(n_245),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_244),
.A2(n_235),
.B1(n_226),
.B2(n_236),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_257),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_236),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_248),
.A2(n_251),
.B1(n_249),
.B2(n_243),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_267),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_259),
.A2(n_245),
.B1(n_242),
.B2(n_252),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_264),
.A2(n_266),
.B1(n_267),
.B2(n_254),
.Y(n_271)
);

AO21x1_ASAP7_75t_L g266 ( 
.A1(n_260),
.A2(n_247),
.B(n_246),
.Y(n_266)
);

INVx11_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

AOI21xp33_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_253),
.B(n_257),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_268),
.B(n_258),
.Y(n_269)
);

AO21x1_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_271),
.B(n_267),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_254),
.C(n_265),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_266),
.C(n_262),
.Y(n_277)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_272),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_265),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_273),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_277),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_270),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_274),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_280),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_281),
.A2(n_278),
.B(n_266),
.Y(n_282)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_282),
.Y(n_283)
);


endmodule