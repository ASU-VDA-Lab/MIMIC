module fake_jpeg_27244_n_298 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_38),
.Y(n_39)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_28),
.B1(n_25),
.B2(n_15),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_38),
.B1(n_33),
.B2(n_34),
.Y(n_64)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_16),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_15),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_35),
.Y(n_68)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_25),
.Y(n_49)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_36),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_38),
.B1(n_28),
.B2(n_33),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_66),
.B1(n_69),
.B2(n_34),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_59),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_16),
.B(n_26),
.C(n_20),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_78),
.B1(n_32),
.B2(n_52),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_68),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_23),
.B(n_34),
.C(n_32),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_38),
.B1(n_33),
.B2(n_31),
.Y(n_69)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_71),
.Y(n_96)
);

FAx1_ASAP7_75t_SL g72 ( 
.A(n_42),
.B(n_31),
.CI(n_34),
.CON(n_72),
.SN(n_72)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_38),
.B1(n_31),
.B2(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

BUFx2_ASAP7_75t_SL g130 ( 
.A(n_82),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_92),
.B1(n_99),
.B2(n_55),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_35),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_107),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_70),
.A2(n_31),
.B1(n_34),
.B2(n_32),
.Y(n_92)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_97),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_69),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_102),
.Y(n_124)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVxp33_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_44),
.B1(n_32),
.B2(n_72),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_109),
.A2(n_112),
.B1(n_135),
.B2(n_36),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_110),
.B(n_123),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_125),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_68),
.B1(n_73),
.B2(n_67),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_103),
.A2(n_57),
.B(n_76),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_113),
.A2(n_129),
.B(n_131),
.Y(n_157)
);

BUFx24_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_17),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_101),
.A2(n_102),
.B1(n_96),
.B2(n_100),
.Y(n_115)
);

BUFx8_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_32),
.B1(n_79),
.B2(n_60),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_117),
.A2(n_86),
.B1(n_87),
.B2(n_104),
.Y(n_142)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_121),
.B(n_122),
.Y(n_144)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_35),
.Y(n_123)
);

BUFx24_ASAP7_75t_SL g125 ( 
.A(n_93),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_126),
.B(n_127),
.Y(n_146)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_91),
.B(n_61),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_132),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_96),
.A2(n_44),
.B1(n_63),
.B2(n_75),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_96),
.A2(n_26),
.B1(n_22),
.B2(n_24),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_106),
.B(n_27),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_81),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_106),
.Y(n_134)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_82),
.A2(n_36),
.B1(n_35),
.B2(n_30),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_138),
.Y(n_176)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_84),
.C(n_94),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_141),
.C(n_158),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_140),
.B(n_143),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_86),
.C(n_95),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_142),
.A2(n_23),
.B1(n_17),
.B2(n_2),
.Y(n_186)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_20),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_145),
.B(n_150),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_87),
.B1(n_104),
.B2(n_18),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_148),
.A2(n_154),
.B1(n_164),
.B2(n_0),
.Y(n_195)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_19),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_20),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_20),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_132),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_30),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_153),
.B(n_165),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_30),
.B1(n_18),
.B2(n_29),
.Y(n_154)
);

FAx1_ASAP7_75t_SL g155 ( 
.A(n_119),
.B(n_36),
.CI(n_29),
.CON(n_155),
.SN(n_155)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_109),
.B(n_37),
.C(n_36),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_114),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_0),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_162),
.B1(n_23),
.B2(n_17),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_127),
.A2(n_36),
.B1(n_30),
.B2(n_18),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_18),
.B1(n_29),
.B2(n_19),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_27),
.Y(n_165)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_167),
.B(n_168),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_118),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_157),
.A2(n_118),
.B(n_120),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_171),
.A2(n_151),
.B(n_155),
.Y(n_204)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_172),
.B(n_175),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_120),
.C(n_135),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_178),
.C(n_180),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_144),
.B(n_114),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_161),
.A2(n_22),
.B1(n_27),
.B2(n_24),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_177),
.A2(n_194),
.B(n_11),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_114),
.C(n_24),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_183),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_22),
.Y(n_180)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_24),
.C(n_19),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_196),
.C(n_6),
.Y(n_205)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_190),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_186),
.A2(n_162),
.B1(n_155),
.B2(n_154),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_149),
.A2(n_146),
.B1(n_157),
.B2(n_148),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_187),
.A2(n_188),
.B1(n_192),
.B2(n_164),
.Y(n_202)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

OAI22x1_ASAP7_75t_L g192 ( 
.A1(n_151),
.A2(n_23),
.B1(n_1),
.B2(n_2),
.Y(n_192)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_151),
.A2(n_14),
.B1(n_7),
.B2(n_9),
.Y(n_194)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_150),
.B(n_9),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_181),
.A2(n_160),
.B1(n_158),
.B2(n_137),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_197),
.A2(n_202),
.B1(n_207),
.B2(n_215),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_173),
.B1(n_185),
.B2(n_182),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_196),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_189),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_209),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_171),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_10),
.C(n_13),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_214),
.Y(n_224)
);

XNOR2x1_ASAP7_75t_SL g212 ( 
.A(n_191),
.B(n_10),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_180),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_174),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_188),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_216),
.B(n_215),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_170),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_217)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_233),
.Y(n_237)
);

OAI22x1_ASAP7_75t_L g221 ( 
.A1(n_212),
.A2(n_192),
.B1(n_177),
.B2(n_194),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_221),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_223),
.B(n_205),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_203),
.Y(n_225)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_227),
.Y(n_242)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_209),
.B(n_169),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_228),
.B(n_232),
.Y(n_245)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_168),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_167),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_191),
.Y(n_244)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_235),
.B(n_199),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_241),
.C(n_219),
.Y(n_259)
);

BUFx24_ASAP7_75t_SL g239 ( 
.A(n_224),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_247),
.Y(n_252)
);

MAJx2_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_211),
.C(n_233),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_248),
.Y(n_254)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_216),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_200),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_238),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_220),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_250),
.B(n_217),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_207),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_231),
.B1(n_218),
.B2(n_222),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_262),
.B1(n_240),
.B2(n_199),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_203),
.Y(n_257)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_259),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_197),
.C(n_231),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_263),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_243),
.B(n_210),
.Y(n_261)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_218),
.B1(n_198),
.B2(n_236),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_258),
.B(n_236),
.Y(n_264)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g279 ( 
.A1(n_264),
.A2(n_11),
.B(n_12),
.C(n_13),
.D(n_14),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_265),
.A2(n_178),
.B1(n_195),
.B2(n_4),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_269),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_237),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_241),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_273),
.B(n_252),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_254),
.C(n_249),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_280),
.Y(n_288)
);

NAND2xp33_ASAP7_75t_SL g275 ( 
.A(n_266),
.B(n_204),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_275),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_277),
.A2(n_279),
.B(n_4),
.Y(n_287)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_278),
.Y(n_283)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_11),
.C(n_12),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_271),
.B(n_267),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_13),
.B1(n_4),
.B2(n_5),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_284),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_287),
.A2(n_276),
.B(n_275),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_289),
.B(n_291),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_274),
.C(n_276),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_281),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_292),
.A2(n_283),
.B(n_286),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_294),
.A2(n_293),
.B(n_285),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_268),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_296),
.B(n_280),
.Y(n_297)
);

NOR3xp33_ASAP7_75t_SL g298 ( 
.A(n_297),
.B(n_278),
.C(n_5),
.Y(n_298)
);


endmodule