module real_jpeg_6789_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_400;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_0),
.Y(n_191)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_0),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_0),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_0),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_1),
.Y(n_129)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_1),
.Y(n_140)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_1),
.Y(n_361)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_1),
.Y(n_407)
);

BUFx5_ASAP7_75t_L g458 ( 
.A(n_1),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_2),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_2),
.A2(n_49),
.B1(n_228),
.B2(n_311),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_2),
.A2(n_49),
.B1(n_288),
.B2(n_388),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g401 ( 
.A1(n_2),
.A2(n_49),
.B1(n_402),
.B2(n_403),
.Y(n_401)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_3),
.Y(n_330)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_3),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_4),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_4),
.A2(n_56),
.B1(n_346),
.B2(n_348),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_4),
.A2(n_56),
.B1(n_391),
.B2(n_393),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_4),
.A2(n_56),
.B1(n_438),
.B2(n_440),
.Y(n_437)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_5),
.Y(n_534)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_6),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_6),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_6),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_6),
.Y(n_174)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_8),
.A2(n_113),
.B1(n_275),
.B2(n_278),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_8),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_8),
.A2(n_253),
.B1(n_278),
.B2(n_371),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_8),
.A2(n_278),
.B1(n_399),
.B2(n_400),
.Y(n_398)
);

OAI22xp33_ASAP7_75t_L g454 ( 
.A1(n_8),
.A2(n_278),
.B1(n_455),
.B2(n_457),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_9),
.Y(n_114)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_9),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_9),
.Y(n_194)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_11),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_12),
.A2(n_82),
.B1(n_84),
.B2(n_87),
.Y(n_81)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_12),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_12),
.A2(n_87),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_12),
.A2(n_87),
.B1(n_201),
.B2(n_220),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_12),
.A2(n_87),
.B1(n_285),
.B2(n_412),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_13),
.A2(n_160),
.B1(n_164),
.B2(n_165),
.Y(n_159)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_13),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_13),
.A2(n_164),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_13),
.A2(n_39),
.B1(n_164),
.B2(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_13),
.A2(n_164),
.B1(n_360),
.B2(n_362),
.Y(n_359)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_14),
.A2(n_179),
.B1(n_185),
.B2(n_186),
.Y(n_178)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_14),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_14),
.A2(n_120),
.B1(n_185),
.B2(n_252),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_14),
.A2(n_185),
.B1(n_366),
.B2(n_368),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_14),
.A2(n_53),
.B1(n_185),
.B2(n_406),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_15),
.A2(n_206),
.B1(n_208),
.B2(n_209),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_15),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_15),
.A2(n_179),
.B1(n_208),
.B2(n_228),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_15),
.A2(n_65),
.B1(n_208),
.B2(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_15),
.A2(n_54),
.B1(n_128),
.B2(n_208),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_16),
.A2(n_90),
.B1(n_92),
.B2(n_94),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_16),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_16),
.A2(n_94),
.B1(n_120),
.B2(n_123),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_16),
.A2(n_94),
.B1(n_126),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_16),
.A2(n_94),
.B1(n_115),
.B2(n_220),
.Y(n_385)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_18),
.A2(n_123),
.B1(n_154),
.B2(n_157),
.Y(n_153)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_18),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_18),
.B(n_172),
.C(n_175),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_18),
.B(n_73),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_18),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_18),
.B(n_118),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_18),
.B(n_266),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_533),
.B(n_535),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_143),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_141),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_133),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_23),
.B(n_133),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_124),
.C(n_130),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_24),
.A2(n_25),
.B1(n_529),
.B2(n_530),
.Y(n_528)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_57),
.C(n_95),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g520 ( 
.A(n_26),
.B(n_521),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_43),
.B1(n_50),
.B2(n_52),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_27),
.A2(n_50),
.B1(n_52),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_27),
.A2(n_50),
.B1(n_125),
.B2(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_27),
.A2(n_358),
.B(n_405),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_27),
.A2(n_50),
.B1(n_405),
.B2(n_426),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_27),
.A2(n_43),
.B1(n_50),
.B2(n_506),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_28),
.A2(n_356),
.B(n_357),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_28),
.B(n_359),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_36),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_37),
.B1(n_39),
.B2(n_42),
.Y(n_36)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_38),
.Y(n_263)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_38),
.Y(n_270)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_40),
.Y(n_400)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_48),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_50),
.B(n_157),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_50),
.A2(n_426),
.B(n_459),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_51),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_51),
.B(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_57),
.A2(n_95),
.B1(n_96),
.B2(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_57),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_81),
.B1(n_88),
.B2(n_89),
.Y(n_57)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_58),
.A2(n_88),
.B1(n_302),
.B2(n_365),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_58),
.A2(n_88),
.B1(n_398),
.B2(n_401),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_58),
.A2(n_81),
.B1(n_88),
.B2(n_510),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_73),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_65),
.B1(n_68),
.B2(n_70),
.Y(n_59)
);

AOI32xp33_ASAP7_75t_L g281 ( 
.A1(n_60),
.A2(n_265),
.A3(n_282),
.B1(n_285),
.B2(n_287),
.Y(n_281)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_65),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_67),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_69),
.Y(n_291)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx6_ASAP7_75t_L g442 ( 
.A(n_72),
.Y(n_442)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_73),
.A2(n_131),
.B(n_132),
.Y(n_130)
);

AOI22x1_ASAP7_75t_L g427 ( 
.A1(n_73),
.A2(n_131),
.B1(n_306),
.B2(n_428),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_73),
.A2(n_131),
.B1(n_436),
.B2(n_437),
.Y(n_435)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_78),
.B2(n_80),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_77),
.Y(n_211)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_77),
.Y(n_256)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_82),
.Y(n_368)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_88),
.B(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_88),
.A2(n_302),
.B(n_305),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_95),
.A2(n_96),
.B1(n_508),
.B2(n_509),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_95),
.B(n_505),
.C(n_508),
.Y(n_516)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_117),
.B(n_119),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_97),
.A2(n_153),
.B(n_158),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_97),
.A2(n_117),
.B1(n_205),
.B2(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_97),
.A2(n_158),
.B(n_251),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_97),
.A2(n_117),
.B1(n_370),
.B2(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_98),
.B(n_159),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_98),
.A2(n_118),
.B1(n_387),
.B2(n_390),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_98),
.A2(n_118),
.B1(n_390),
.B2(n_411),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_98),
.A2(n_118),
.B1(n_411),
.B2(n_445),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_110),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_105),
.B2(n_107),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_109),
.Y(n_289)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_110),
.A2(n_205),
.B(n_212),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_110)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_114),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_117),
.A2(n_212),
.B(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_118),
.B(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_119),
.Y(n_445)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_122),
.Y(n_371)
);

INVx6_ASAP7_75t_L g395 ( 
.A(n_122),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_124),
.B(n_130),
.Y(n_530)
);

OAI21xp33_ASAP7_75t_SL g356 ( 
.A1(n_127),
.A2(n_157),
.B(n_337),
.Y(n_356)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_131),
.A2(n_259),
.B(n_267),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_131),
.B(n_306),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_131),
.A2(n_267),
.B(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_140),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_527),
.B(n_532),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_498),
.B(n_524),
.Y(n_144)
);

OAI311xp33_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_374),
.A3(n_474),
.B1(n_492),
.C1(n_493),
.Y(n_145)
);

AOI21x1_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_316),
.B(n_373),
.Y(n_146)
);

AO21x1_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_293),
.B(n_315),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_245),
.B(n_292),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_215),
.B(n_244),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_176),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_151),
.B(n_176),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_167),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_152),
.A2(n_167),
.B1(n_168),
.B2(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_152),
.Y(n_242)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_155),
.Y(n_207)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_156),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_157),
.A2(n_189),
.B(n_195),
.Y(n_224)
);

OAI21xp33_ASAP7_75t_SL g259 ( 
.A1(n_157),
.A2(n_260),
.B(n_264),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_157),
.B(n_328),
.Y(n_337)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_163),
.Y(n_170)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_163),
.Y(n_414)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_202),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_177),
.B(n_203),
.C(n_214),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_189),
.B(n_195),
.Y(n_177)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_178),
.Y(n_240)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_183),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_184),
.Y(n_231)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_188),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_189),
.A2(n_340),
.B1(n_341),
.B2(n_344),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_189),
.A2(n_380),
.B1(n_381),
.B2(n_385),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_189),
.A2(n_383),
.B(n_385),
.Y(n_415)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_199),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_190),
.A2(n_233),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_190),
.A2(n_274),
.B1(n_310),
.B2(n_312),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_190),
.A2(n_345),
.B1(n_422),
.B2(n_423),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx8_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_198),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_198),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_213),
.B2(n_214),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_237),
.B(n_243),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_225),
.B(n_236),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_224),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_221),
.Y(n_349)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_223),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_235),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_235),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_232),
.B(n_234),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_227),
.Y(n_239)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_230),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_234),
.A2(n_273),
.B(n_279),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_241),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_246),
.B(n_247),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_271),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_257),
.B2(n_258),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_250),
.B(n_257),
.C(n_271),
.Y(n_294)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx5_ASAP7_75t_SL g253 ( 
.A(n_254),
.Y(n_253)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_255),
.Y(n_389)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_260),
.Y(n_402)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_263),
.Y(n_304)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_263),
.Y(n_325)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_263),
.Y(n_336)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_268),
.Y(n_306)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_281),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_281),
.Y(n_299)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_SL g279 ( 
.A(n_280),
.Y(n_279)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

NAND2xp33_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

INVx4_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_294),
.B(n_295),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_300),
.B2(n_314),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_299),
.C(n_314),
.Y(n_317)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_307),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_301),
.B(n_308),
.C(n_309),
.Y(n_350)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_310),
.Y(n_340)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_317),
.B(n_318),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_353),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_350),
.B1(n_351),
.B2(n_352),
.Y(n_319)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_320),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_338),
.B2(n_339),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_322),
.B(n_338),
.Y(n_470)
);

OAI32xp33_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_326),
.A3(n_329),
.B1(n_331),
.B2(n_337),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_328),
.Y(n_362)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_335),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_343),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_350),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_350),
.B(n_351),
.C(n_353),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_355),
.B1(n_363),
.B2(n_372),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_354),
.B(n_364),
.C(n_369),
.Y(n_483)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx6_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_363),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_369),
.Y(n_363)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_365),
.Y(n_472)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_366),
.Y(n_403)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx5_ASAP7_75t_L g439 ( 
.A(n_367),
.Y(n_439)
);

INVx11_ASAP7_75t_L g392 ( 
.A(n_371),
.Y(n_392)
);

NAND2xp33_ASAP7_75t_SL g374 ( 
.A(n_375),
.B(n_460),
.Y(n_374)
);

A2O1A1Ixp33_ASAP7_75t_SL g493 ( 
.A1(n_375),
.A2(n_460),
.B(n_494),
.C(n_497),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_429),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_376),
.B(n_429),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_408),
.C(n_417),
.Y(n_376)
);

FAx1_ASAP7_75t_SL g473 ( 
.A(n_377),
.B(n_408),
.CI(n_417),
.CON(n_473),
.SN(n_473)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_396),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_378),
.B(n_397),
.C(n_404),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_386),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_379),
.B(n_386),
.Y(n_466)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_380),
.Y(n_422)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx8_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_387),
.Y(n_420)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx3_ASAP7_75t_SL g393 ( 
.A(n_394),
.Y(n_393)
);

INVx8_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_404),
.Y(n_396)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_398),
.Y(n_428)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_401),
.Y(n_436)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_406),
.Y(n_456)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_409),
.A2(n_410),
.B1(n_415),
.B2(n_416),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_410),
.B(n_415),
.Y(n_449)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_415),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_415),
.A2(n_416),
.B1(n_451),
.B2(n_452),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_415),
.A2(n_449),
.B(n_452),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_424),
.C(n_427),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_418),
.B(n_464),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_419),
.B(n_421),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_419),
.B(n_421),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_424),
.A2(n_425),
.B1(n_427),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_427),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_430),
.B(n_433),
.C(n_447),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_433),
.B1(n_447),
.B2(n_448),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_434),
.A2(n_443),
.B(n_446),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_435),
.B(n_444),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_437),
.Y(n_510)
);

INVx4_ASAP7_75t_SL g438 ( 
.A(n_439),
.Y(n_438)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_446),
.B(n_503),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_446),
.B(n_501),
.C(n_503),
.Y(n_523)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_459),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_454),
.Y(n_506)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_473),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_461),
.B(n_473),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_466),
.C(n_467),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_462),
.A2(n_463),
.B1(n_466),
.B2(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_466),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_467),
.B(n_485),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_470),
.C(n_471),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_468),
.A2(n_469),
.B1(n_471),
.B2(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_470),
.B(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_471),
.Y(n_480)
);

BUFx24_ASAP7_75t_SL g540 ( 
.A(n_473),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_487),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_476),
.A2(n_495),
.B(n_496),
.Y(n_494)
);

NOR2x1_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_484),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_477),
.B(n_484),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_481),
.C(n_483),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_478),
.B(n_490),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_481),
.A2(n_482),
.B1(n_483),
.B2(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_483),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_488),
.B(n_489),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_513),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_500),
.B(n_512),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_500),
.B(n_512),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_502),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_504),
.A2(n_505),
.B1(n_507),
.B2(n_511),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_504),
.A2(n_505),
.B1(n_519),
.B2(n_520),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_504),
.B(n_515),
.C(n_519),
.Y(n_531)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_507),
.Y(n_511)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_513),
.A2(n_525),
.B(n_526),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_514),
.B(n_523),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_514),
.B(n_523),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_515),
.A2(n_516),
.B1(n_517),
.B2(n_518),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_531),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_528),
.B(n_531),
.Y(n_532)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx8_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx13_ASAP7_75t_L g537 ( 
.A(n_534),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_536),
.B(n_538),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);


endmodule