module fake_jpeg_900_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_SL g8 ( 
.A(n_3),
.B(n_1),
.Y(n_8)
);

INVxp67_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_21),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_0),
.C(n_1),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_23),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g19 ( 
.A(n_10),
.B(n_11),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_19),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_5),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_4),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_8),
.B(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_22),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_3),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_17),
.A2(n_14),
.B1(n_11),
.B2(n_12),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_SL g37 ( 
.A1(n_24),
.A2(n_15),
.B(n_13),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_4),
.Y(n_39)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_12),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_14),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_40),
.B1(n_24),
.B2(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_39),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_15),
.B(n_31),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_46),
.B1(n_40),
.B2(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_38),
.B1(n_26),
.B2(n_25),
.Y(n_48)
);

XNOR2x1_ASAP7_75t_SL g50 ( 
.A(n_48),
.B(n_26),
.Y(n_50)
);

AOI322xp5_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_42),
.A3(n_27),
.B1(n_32),
.B2(n_45),
.C1(n_44),
.C2(n_35),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_42),
.B(n_49),
.Y(n_52)
);

NOR3xp33_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_32),
.C(n_34),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_41),
.Y(n_54)
);


endmodule