module fake_jpeg_8447_n_95 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_95);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_95;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx5_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx6_ASAP7_75t_SL g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_12),
.B(n_0),
.Y(n_23)
);

OR2x4_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_1),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_17),
.B1(n_12),
.B2(n_15),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

MAJx2_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_13),
.C(n_17),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

AO22x1_ASAP7_75t_SL g29 ( 
.A1(n_22),
.A2(n_13),
.B1(n_17),
.B2(n_3),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_12),
.B1(n_15),
.B2(n_19),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_20),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_SL g55 ( 
.A1(n_35),
.A2(n_36),
.B(n_14),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_24),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_42),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_27),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_51),
.B(n_54),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_19),
.B(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_52),
.B(n_14),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_22),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_22),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_19),
.B(n_16),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_55),
.B(n_14),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_57),
.B(n_62),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_61),
.C(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_63),
.Y(n_71)
);

MAJx2_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_53),
.C(n_51),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_18),
.Y(n_63)
);

OA21x2_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_33),
.B(n_17),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_64),
.A2(n_25),
.B1(n_21),
.B2(n_32),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_47),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_68),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_64),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_72),
.Y(n_73)
);

AO21x1_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_17),
.B(n_26),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_21),
.B1(n_25),
.B2(n_49),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_70),
.A2(n_11),
.B1(n_56),
.B2(n_26),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_64),
.Y(n_72)
);

MAJx2_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_61),
.C(n_68),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_72),
.C(n_67),
.Y(n_83)
);

AO221x1_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_17),
.B1(n_2),
.B2(n_4),
.C(n_1),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_18),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_77),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_69),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_56),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_80),
.A2(n_84),
.B(n_74),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_78),
.B(n_77),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_86),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_82),
.B(n_9),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_82),
.A2(n_6),
.B(n_8),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_9),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_91),
.B(n_1),
.Y(n_92)
);

OAI21x1_ASAP7_75t_SL g94 ( 
.A1(n_92),
.A2(n_93),
.B(n_4),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_90),
.A2(n_2),
.B1(n_4),
.B2(n_26),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_26),
.Y(n_95)
);


endmodule