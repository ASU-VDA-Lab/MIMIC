module real_aes_7037_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_363;
wire n_754;
wire n_182;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_0), .B(n_109), .C(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g128 ( .A(n_0), .Y(n_128) );
INVx1_ASAP7_75t_L g518 ( .A(n_1), .Y(n_518) );
INVx1_ASAP7_75t_L g159 ( .A(n_2), .Y(n_159) );
OAI22xp5_ASAP7_75t_SL g741 ( .A1(n_3), .A2(n_742), .B1(n_745), .B2(n_746), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_3), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g129 ( .A1(n_4), .A2(n_130), .B1(n_131), .B2(n_454), .Y(n_129) );
INVx1_ASAP7_75t_L g454 ( .A(n_4), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_5), .A2(n_40), .B1(n_184), .B2(n_474), .Y(n_503) );
AOI21xp33_ASAP7_75t_L g203 ( .A1(n_6), .A2(n_175), .B(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_7), .B(n_173), .Y(n_529) );
AND2x6_ASAP7_75t_L g152 ( .A(n_8), .B(n_153), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_9), .A2(n_257), .B(n_258), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_10), .B(n_41), .Y(n_114) );
INVx1_ASAP7_75t_L g209 ( .A(n_11), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_12), .B(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g144 ( .A(n_13), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_14), .B(n_165), .Y(n_482) );
INVx1_ASAP7_75t_L g263 ( .A(n_15), .Y(n_263) );
INVx1_ASAP7_75t_L g512 ( .A(n_16), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_17), .B(n_140), .Y(n_534) );
AO32x2_ASAP7_75t_L g501 ( .A1(n_18), .A2(n_139), .A3(n_173), .B1(n_476), .B2(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_19), .B(n_184), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_20), .B(n_180), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_21), .B(n_140), .Y(n_520) );
OAI22xp5_ASAP7_75t_SL g450 ( .A1(n_22), .A2(n_33), .B1(n_451), .B2(n_452), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_22), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_23), .A2(n_52), .B1(n_184), .B2(n_474), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_24), .B(n_175), .Y(n_220) );
AOI22xp33_ASAP7_75t_SL g475 ( .A1(n_25), .A2(n_79), .B1(n_165), .B2(n_184), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_26), .B(n_184), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_27), .B(n_187), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_28), .A2(n_261), .B(n_262), .C(n_264), .Y(n_260) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_29), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_30), .B(n_170), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_31), .B(n_163), .Y(n_162) );
AOI222xp33_ASAP7_75t_L g459 ( .A1(n_32), .A2(n_460), .B1(n_741), .B2(n_747), .C1(n_750), .C2(n_751), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_33), .Y(n_452) );
INVx1_ASAP7_75t_L g198 ( .A(n_34), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_35), .B(n_170), .Y(n_499) );
INVx2_ASAP7_75t_L g150 ( .A(n_36), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_37), .B(n_184), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_38), .B(n_170), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_39), .A2(n_152), .B(n_155), .C(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g196 ( .A(n_42), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_43), .B(n_163), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_44), .B(n_184), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_45), .B(n_456), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_46), .A2(n_89), .B1(n_227), .B2(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_47), .B(n_184), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_48), .B(n_184), .Y(n_513) );
CKINVDCx16_ASAP7_75t_R g199 ( .A(n_49), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_50), .B(n_517), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_51), .B(n_175), .Y(n_240) );
AOI22xp33_ASAP7_75t_SL g538 ( .A1(n_53), .A2(n_62), .B1(n_165), .B2(n_184), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_54), .A2(n_155), .B1(n_165), .B2(n_194), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_55), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_56), .B(n_184), .Y(n_481) );
CKINVDCx16_ASAP7_75t_R g146 ( .A(n_57), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_58), .B(n_184), .Y(n_552) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_59), .A2(n_183), .B(n_207), .C(n_208), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_60), .Y(n_254) );
INVx1_ASAP7_75t_L g205 ( .A(n_61), .Y(n_205) );
INVx1_ASAP7_75t_L g153 ( .A(n_63), .Y(n_153) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_64), .A2(n_104), .B1(n_115), .B2(n_754), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_65), .B(n_184), .Y(n_519) );
INVx1_ASAP7_75t_L g143 ( .A(n_66), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_67), .Y(n_120) );
AO32x2_ASAP7_75t_L g471 ( .A1(n_68), .A2(n_173), .A3(n_232), .B1(n_472), .B2(n_476), .Y(n_471) );
INVx1_ASAP7_75t_L g551 ( .A(n_69), .Y(n_551) );
INVx1_ASAP7_75t_L g494 ( .A(n_70), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_71), .A2(n_78), .B1(n_743), .B2(n_744), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_71), .Y(n_744) );
A2O1A1Ixp33_ASAP7_75t_SL g179 ( .A1(n_72), .A2(n_180), .B(n_181), .C(n_183), .Y(n_179) );
INVxp67_ASAP7_75t_L g182 ( .A(n_73), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_74), .B(n_165), .Y(n_495) );
INVx1_ASAP7_75t_L g112 ( .A(n_75), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_76), .Y(n_201) );
INVx1_ASAP7_75t_L g247 ( .A(n_77), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_78), .Y(n_743) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_80), .A2(n_152), .B(n_155), .C(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_81), .B(n_474), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_82), .B(n_165), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_83), .B(n_160), .Y(n_223) );
INVx2_ASAP7_75t_L g141 ( .A(n_84), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_85), .B(n_180), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_86), .B(n_165), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_87), .A2(n_152), .B(n_155), .C(n_158), .Y(n_154) );
INVx2_ASAP7_75t_L g109 ( .A(n_88), .Y(n_109) );
OR2x2_ASAP7_75t_L g125 ( .A(n_88), .B(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g463 ( .A(n_88), .B(n_127), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_90), .A2(n_102), .B1(n_165), .B2(n_166), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_91), .B(n_170), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_92), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_93), .A2(n_152), .B(n_155), .C(n_235), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_94), .Y(n_242) );
INVx1_ASAP7_75t_L g178 ( .A(n_95), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_96), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_97), .B(n_160), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_98), .B(n_165), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_99), .B(n_173), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_100), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_101), .A2(n_175), .B(n_176), .Y(n_174) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_107), .Y(n_755) );
OR2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_113), .Y(n_107) );
OR2x2_ASAP7_75t_L g740 ( .A(n_109), .B(n_127), .Y(n_740) );
NOR2x2_ASAP7_75t_L g753 ( .A(n_109), .B(n_126), .Y(n_753) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVxp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g127 ( .A(n_114), .B(n_128), .Y(n_127) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_458), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
NAND3xp33_ASAP7_75t_L g458 ( .A(n_117), .B(n_455), .C(n_459), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_129), .B(n_455), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_125), .Y(n_457) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_449), .B1(n_450), .B2(n_453), .Y(n_131) );
INVx2_ASAP7_75t_L g453 ( .A(n_132), .Y(n_453) );
OAI22xp5_ASAP7_75t_SL g460 ( .A1(n_132), .A2(n_461), .B1(n_464), .B2(n_738), .Y(n_460) );
OR4x1_ASAP7_75t_L g132 ( .A(n_133), .B(n_338), .C(n_398), .D(n_425), .Y(n_132) );
NAND4xp25_ASAP7_75t_SL g133 ( .A(n_134), .B(n_286), .C(n_317), .D(n_334), .Y(n_133) );
O2A1O1Ixp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_211), .B(n_213), .C(n_266), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_189), .Y(n_135) );
INVx1_ASAP7_75t_L g328 ( .A(n_136), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_136), .A2(n_369), .B1(n_417), .B2(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_171), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_137), .B(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g279 ( .A(n_137), .B(n_191), .Y(n_279) );
AND2x2_ASAP7_75t_L g321 ( .A(n_137), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_137), .B(n_212), .Y(n_333) );
INVx1_ASAP7_75t_L g373 ( .A(n_137), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_137), .B(n_427), .Y(n_426) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g301 ( .A(n_138), .B(n_191), .Y(n_301) );
INVx3_ASAP7_75t_L g305 ( .A(n_138), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_138), .B(n_363), .Y(n_362) );
AO21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_145), .B(n_167), .Y(n_138) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_139), .A2(n_192), .B(n_200), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_139), .B(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g228 ( .A(n_139), .Y(n_228) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_140), .Y(n_173) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_SL g170 ( .A(n_141), .B(n_142), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
OAI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_154), .Y(n_145) );
OAI22xp33_ASAP7_75t_L g192 ( .A1(n_147), .A2(n_185), .B1(n_193), .B2(n_199), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g246 ( .A1(n_147), .A2(n_247), .B(n_248), .Y(n_246) );
NAND2x1p5_ASAP7_75t_L g147 ( .A(n_148), .B(n_152), .Y(n_147) );
AND2x4_ASAP7_75t_L g175 ( .A(n_148), .B(n_152), .Y(n_175) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx1_ASAP7_75t_L g517 ( .A(n_149), .Y(n_517) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
INVx1_ASAP7_75t_L g166 ( .A(n_150), .Y(n_166) );
INVx1_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
INVx3_ASAP7_75t_L g161 ( .A(n_151), .Y(n_161) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_151), .Y(n_163) );
INVx1_ASAP7_75t_L g180 ( .A(n_151), .Y(n_180) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_151), .Y(n_195) );
INVx4_ASAP7_75t_SL g185 ( .A(n_152), .Y(n_185) );
BUFx3_ASAP7_75t_L g476 ( .A(n_152), .Y(n_476) );
OAI21xp5_ASAP7_75t_L g479 ( .A1(n_152), .A2(n_480), .B(n_484), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_152), .A2(n_493), .B(n_496), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_152), .A2(n_511), .B(n_515), .Y(n_510) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_152), .A2(n_523), .B(n_526), .Y(n_522) );
INVx5_ASAP7_75t_L g177 ( .A(n_155), .Y(n_177) );
AND2x6_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_156), .Y(n_184) );
BUFx3_ASAP7_75t_L g227 ( .A(n_156), .Y(n_227) );
INVx1_ASAP7_75t_L g474 ( .A(n_156), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_162), .C(n_164), .Y(n_158) );
O2A1O1Ixp5_ASAP7_75t_SL g493 ( .A1(n_160), .A2(n_183), .B(n_494), .C(n_495), .Y(n_493) );
INVx2_ASAP7_75t_L g504 ( .A(n_160), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_160), .A2(n_524), .B(n_525), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_160), .A2(n_548), .B(n_549), .Y(n_547) );
INVx5_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_161), .B(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_161), .B(n_209), .Y(n_208) );
OAI22xp5_ASAP7_75t_SL g472 ( .A1(n_161), .A2(n_163), .B1(n_473), .B2(n_475), .Y(n_472) );
INVx2_ASAP7_75t_L g207 ( .A(n_163), .Y(n_207) );
INVx4_ASAP7_75t_L g238 ( .A(n_163), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_163), .A2(n_503), .B1(n_504), .B2(n_505), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_163), .A2(n_504), .B1(n_537), .B2(n_538), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_164), .A2(n_512), .B(n_513), .C(n_514), .Y(n_511) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_169), .B(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_169), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g232 ( .A(n_170), .Y(n_232) );
OA21x2_ASAP7_75t_L g255 ( .A1(n_170), .A2(n_256), .B(n_265), .Y(n_255) );
OA21x2_ASAP7_75t_L g478 ( .A1(n_170), .A2(n_479), .B(n_487), .Y(n_478) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_170), .A2(n_492), .B(n_499), .Y(n_491) );
AND2x2_ASAP7_75t_L g392 ( .A(n_171), .B(n_202), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_171), .B(n_305), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_171), .B(n_420), .Y(n_419) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g212 ( .A(n_172), .B(n_191), .Y(n_212) );
INVx1_ASAP7_75t_L g274 ( .A(n_172), .Y(n_274) );
BUFx2_ASAP7_75t_L g278 ( .A(n_172), .Y(n_278) );
AND2x2_ASAP7_75t_L g322 ( .A(n_172), .B(n_190), .Y(n_322) );
OR2x2_ASAP7_75t_L g361 ( .A(n_172), .B(n_190), .Y(n_361) );
AND2x2_ASAP7_75t_L g386 ( .A(n_172), .B(n_202), .Y(n_386) );
AND2x2_ASAP7_75t_L g445 ( .A(n_172), .B(n_275), .Y(n_445) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_186), .Y(n_172) );
INVx4_ASAP7_75t_L g188 ( .A(n_173), .Y(n_188) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_173), .A2(n_522), .B(n_529), .Y(n_521) );
BUFx2_ASAP7_75t_L g257 ( .A(n_175), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_179), .C(n_185), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g204 ( .A1(n_177), .A2(n_185), .B(n_205), .C(n_206), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_177), .A2(n_185), .B(n_259), .C(n_260), .Y(n_258) );
INVx1_ASAP7_75t_L g483 ( .A(n_180), .Y(n_483) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_184), .Y(n_239) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_187), .A2(n_203), .B(n_210), .Y(n_202) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_SL g229 ( .A(n_188), .B(n_230), .Y(n_229) );
NAND3xp33_ASAP7_75t_L g535 ( .A(n_188), .B(n_476), .C(n_536), .Y(n_535) );
AO21x1_ASAP7_75t_L g582 ( .A1(n_188), .A2(n_536), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g420 ( .A(n_189), .Y(n_420) );
OR2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_202), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_190), .B(n_202), .Y(n_306) );
AND2x2_ASAP7_75t_L g316 ( .A(n_190), .B(n_305), .Y(n_316) );
BUFx2_ASAP7_75t_L g327 ( .A(n_190), .Y(n_327) );
INVx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g349 ( .A(n_191), .B(n_202), .Y(n_349) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_191), .Y(n_404) );
OAI22xp5_ASAP7_75t_SL g194 ( .A1(n_195), .A2(n_196), .B1(n_197), .B2(n_198), .Y(n_194) );
INVx2_ASAP7_75t_L g197 ( .A(n_195), .Y(n_197) );
INVx4_ASAP7_75t_L g261 ( .A(n_195), .Y(n_261) );
AND2x2_ASAP7_75t_SL g211 ( .A(n_202), .B(n_212), .Y(n_211) );
INVx1_ASAP7_75t_SL g275 ( .A(n_202), .Y(n_275) );
BUFx2_ASAP7_75t_L g300 ( .A(n_202), .Y(n_300) );
INVx2_ASAP7_75t_L g319 ( .A(n_202), .Y(n_319) );
AND2x2_ASAP7_75t_L g381 ( .A(n_202), .B(n_305), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_207), .A2(n_485), .B(n_486), .Y(n_484) );
O2A1O1Ixp5_ASAP7_75t_L g550 ( .A1(n_207), .A2(n_516), .B(n_551), .C(n_552), .Y(n_550) );
AOI321xp33_ASAP7_75t_L g400 ( .A1(n_211), .A2(n_401), .A3(n_402), .B1(n_403), .B2(n_405), .C(n_406), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_212), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_212), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g394 ( .A(n_212), .B(n_373), .Y(n_394) );
AND2x2_ASAP7_75t_L g427 ( .A(n_212), .B(n_319), .Y(n_427) );
INVx1_ASAP7_75t_SL g213 ( .A(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_243), .Y(n_214) );
OR2x2_ASAP7_75t_L g329 ( .A(n_215), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_231), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx3_ASAP7_75t_L g281 ( .A(n_218), .Y(n_281) );
AND2x2_ASAP7_75t_L g291 ( .A(n_218), .B(n_245), .Y(n_291) );
AND2x2_ASAP7_75t_L g296 ( .A(n_218), .B(n_271), .Y(n_296) );
INVx1_ASAP7_75t_L g313 ( .A(n_218), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_218), .B(n_294), .Y(n_332) );
AND2x2_ASAP7_75t_L g337 ( .A(n_218), .B(n_270), .Y(n_337) );
OR2x2_ASAP7_75t_L g369 ( .A(n_218), .B(n_358), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_218), .B(n_282), .Y(n_408) );
AND2x2_ASAP7_75t_L g442 ( .A(n_218), .B(n_268), .Y(n_442) );
OR2x6_ASAP7_75t_L g218 ( .A(n_219), .B(n_229), .Y(n_218) );
AOI21xp5_ASAP7_75t_SL g219 ( .A1(n_220), .A2(n_221), .B(n_228), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_225), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_225), .A2(n_250), .B(n_251), .Y(n_249) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g264 ( .A(n_227), .Y(n_264) );
INVx1_ASAP7_75t_L g252 ( .A(n_228), .Y(n_252) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_228), .A2(n_510), .B(n_520), .Y(n_509) );
OA21x2_ASAP7_75t_L g545 ( .A1(n_228), .A2(n_546), .B(n_553), .Y(n_545) );
INVx1_ASAP7_75t_L g269 ( .A(n_231), .Y(n_269) );
INVx2_ASAP7_75t_L g284 ( .A(n_231), .Y(n_284) );
AND2x2_ASAP7_75t_L g324 ( .A(n_231), .B(n_295), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_231), .B(n_271), .Y(n_346) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_241), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_240), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_239), .Y(n_235) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g430 ( .A(n_244), .B(n_281), .Y(n_430) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_255), .Y(n_244) );
INVx2_ASAP7_75t_L g271 ( .A(n_245), .Y(n_271) );
AND2x2_ASAP7_75t_L g424 ( .A(n_245), .B(n_284), .Y(n_424) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_252), .B(n_253), .Y(n_245) );
AND2x2_ASAP7_75t_L g270 ( .A(n_255), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g285 ( .A(n_255), .Y(n_285) );
INVx1_ASAP7_75t_L g295 ( .A(n_255), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_261), .B(n_263), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_261), .A2(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g514 ( .A(n_261), .Y(n_514) );
OAI22xp33_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_272), .B1(n_276), .B2(n_280), .Y(n_266) );
OAI22xp33_ASAP7_75t_L g421 ( .A1(n_267), .A2(n_385), .B1(n_422), .B2(n_423), .Y(n_421) );
INVx1_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx1_ASAP7_75t_L g336 ( .A(n_269), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_270), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g331 ( .A(n_271), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_271), .B(n_284), .Y(n_358) );
INVx1_ASAP7_75t_L g374 ( .A(n_271), .Y(n_374) );
AND2x2_ASAP7_75t_L g315 ( .A(n_273), .B(n_316), .Y(n_315) );
INVx3_ASAP7_75t_SL g354 ( .A(n_273), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_273), .B(n_279), .Y(n_431) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx1_ASAP7_75t_L g440 ( .A(n_276), .Y(n_440) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_277), .B(n_373), .Y(n_415) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx3_ASAP7_75t_SL g320 ( .A(n_279), .Y(n_320) );
NAND2x1_ASAP7_75t_SL g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AND2x2_ASAP7_75t_L g341 ( .A(n_281), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g348 ( .A(n_281), .B(n_285), .Y(n_348) );
AND2x2_ASAP7_75t_L g353 ( .A(n_281), .B(n_294), .Y(n_353) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_281), .Y(n_402) );
OAI311xp33_ASAP7_75t_L g425 ( .A1(n_282), .A2(n_426), .A3(n_428), .B1(n_429), .C1(n_439), .Y(n_425) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g438 ( .A(n_283), .B(n_311), .Y(n_438) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x2_ASAP7_75t_L g294 ( .A(n_284), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g342 ( .A(n_284), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g397 ( .A(n_284), .Y(n_397) );
INVx1_ASAP7_75t_L g290 ( .A(n_285), .Y(n_290) );
INVx1_ASAP7_75t_L g310 ( .A(n_285), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_285), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g343 ( .A(n_285), .Y(n_343) );
AOI221xp5_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_289), .B1(n_297), .B2(n_302), .C(n_307), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_292), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx4_ASAP7_75t_L g311 ( .A(n_291), .Y(n_311) );
AND2x2_ASAP7_75t_L g405 ( .A(n_291), .B(n_324), .Y(n_405) );
AND2x2_ASAP7_75t_L g412 ( .A(n_291), .B(n_294), .Y(n_412) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_294), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g323 ( .A(n_296), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_299), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g448 ( .A(n_301), .B(n_392), .Y(n_448) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g433 ( .A(n_305), .B(n_361), .Y(n_433) );
OAI211xp5_ASAP7_75t_L g398 ( .A1(n_306), .A2(n_399), .B(n_400), .C(n_413), .Y(n_398) );
AOI21xp33_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_312), .B(n_314), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NOR2xp67_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g377 ( .A(n_311), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g406 ( .A1(n_312), .A2(n_407), .B1(n_408), .B2(n_409), .C(n_410), .Y(n_406) );
AND2x2_ASAP7_75t_L g383 ( .A(n_313), .B(n_324), .Y(n_383) );
AND2x2_ASAP7_75t_L g436 ( .A(n_313), .B(n_331), .Y(n_436) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_316), .B(n_354), .Y(n_378) );
O2A1O1Ixp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_321), .B(n_323), .C(n_325), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g364 ( .A(n_319), .B(n_322), .Y(n_364) );
OR2x2_ASAP7_75t_L g407 ( .A(n_319), .B(n_361), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_320), .B(n_386), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_320), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g351 ( .A(n_321), .Y(n_351) );
INVx1_ASAP7_75t_L g417 ( .A(n_324), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_329), .B1(n_332), .B2(n_333), .Y(n_325) );
INVx1_ASAP7_75t_L g340 ( .A(n_326), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_327), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g403 ( .A(n_328), .B(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g389 ( .A(n_330), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_331), .B(n_417), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g390 ( .A1(n_332), .A2(n_391), .B1(n_393), .B2(n_395), .Y(n_390) );
INVx1_ASAP7_75t_L g399 ( .A(n_335), .Y(n_399) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
AND2x2_ASAP7_75t_L g441 ( .A(n_336), .B(n_436), .Y(n_441) );
AOI222xp33_ASAP7_75t_L g370 ( .A1(n_337), .A2(n_371), .B1(n_374), .B2(n_375), .C1(n_378), .C2(n_379), .Y(n_370) );
NAND4xp25_ASAP7_75t_SL g338 ( .A(n_339), .B(n_359), .C(n_370), .D(n_382), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B1(n_344), .B2(n_349), .C(n_350), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_342), .B(n_377), .Y(n_376) );
INVxp67_ASAP7_75t_L g368 ( .A(n_343), .Y(n_368) );
AOI221xp5_ASAP7_75t_L g413 ( .A1(n_344), .A2(n_414), .B1(n_416), .B2(n_418), .C(n_421), .Y(n_413) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g356 ( .A(n_348), .B(n_357), .Y(n_356) );
OAI21xp33_ASAP7_75t_L g410 ( .A1(n_349), .A2(n_411), .B(n_412), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_352), .B1(n_354), .B2(n_355), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI21xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_362), .B(n_365), .Y(n_359) );
INVxp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g401 ( .A(n_372), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_373), .B(n_392), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_373), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_377), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_SL g409 ( .A(n_381), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B1(n_387), .B2(n_389), .C(n_390), .Y(n_382) );
INVxp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI222xp33_ASAP7_75t_L g429 ( .A1(n_392), .A2(n_430), .B1(n_431), .B2(n_432), .C1(n_434), .C2(n_437), .Y(n_429) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_396), .B(n_436), .Y(n_435) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g428 ( .A(n_402), .Y(n_428) );
INVxp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVxp33_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B1(n_442), .B2(n_443), .C(n_446), .Y(n_439) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVxp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_453), .A2(n_461), .B1(n_748), .B2(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g749 ( .A(n_464), .Y(n_749) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND3x1_ASAP7_75t_L g465 ( .A(n_466), .B(n_658), .C(n_706), .Y(n_465) );
NOR4xp25_ASAP7_75t_L g466 ( .A(n_467), .B(n_586), .C(n_631), .D(n_645), .Y(n_466) );
OAI311xp33_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_506), .A3(n_530), .B1(n_539), .C1(n_554), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_477), .Y(n_468) );
OAI21xp33_ASAP7_75t_L g539 ( .A1(n_469), .A2(n_540), .B(n_542), .Y(n_539) );
AND2x2_ASAP7_75t_L g647 ( .A(n_469), .B(n_574), .Y(n_647) );
AND2x2_ASAP7_75t_L g704 ( .A(n_469), .B(n_590), .Y(n_704) );
BUFx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g597 ( .A(n_470), .B(n_500), .Y(n_597) );
AND2x2_ASAP7_75t_L g654 ( .A(n_470), .B(n_602), .Y(n_654) );
INVx1_ASAP7_75t_L g695 ( .A(n_470), .Y(n_695) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_471), .Y(n_563) );
AND2x2_ASAP7_75t_L g604 ( .A(n_471), .B(n_500), .Y(n_604) );
AND2x2_ASAP7_75t_L g608 ( .A(n_471), .B(n_501), .Y(n_608) );
INVx1_ASAP7_75t_L g620 ( .A(n_471), .Y(n_620) );
OAI21xp5_ASAP7_75t_L g546 ( .A1(n_476), .A2(n_547), .B(n_550), .Y(n_546) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_488), .Y(n_477) );
AND2x2_ASAP7_75t_L g541 ( .A(n_478), .B(n_500), .Y(n_541) );
INVx2_ASAP7_75t_L g575 ( .A(n_478), .Y(n_575) );
AND2x2_ASAP7_75t_L g590 ( .A(n_478), .B(n_501), .Y(n_590) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_478), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_478), .B(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g610 ( .A(n_478), .B(n_573), .Y(n_610) );
INVx1_ASAP7_75t_L g622 ( .A(n_478), .Y(n_622) );
INVx1_ASAP7_75t_L g663 ( .A(n_478), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_478), .B(n_563), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B(n_483), .Y(n_480) );
NOR2xp67_ASAP7_75t_L g488 ( .A(n_489), .B(n_500), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g540 ( .A(n_490), .B(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_490), .Y(n_568) );
AND2x2_ASAP7_75t_SL g621 ( .A(n_490), .B(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g625 ( .A(n_490), .B(n_500), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_490), .B(n_620), .Y(n_683) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g573 ( .A(n_491), .Y(n_573) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_491), .Y(n_589) );
OR2x2_ASAP7_75t_L g662 ( .A(n_491), .B(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx2_ASAP7_75t_L g569 ( .A(n_501), .Y(n_569) );
AND2x2_ASAP7_75t_L g574 ( .A(n_501), .B(n_575), .Y(n_574) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_504), .A2(n_516), .B(n_518), .C(n_519), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_504), .A2(n_527), .B(n_528), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_506), .B(n_557), .Y(n_720) );
INVx1_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
OR2x2_ASAP7_75t_L g690 ( .A(n_507), .B(n_532), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_521), .Y(n_507) );
AND2x2_ASAP7_75t_L g566 ( .A(n_508), .B(n_557), .Y(n_566) );
INVx2_ASAP7_75t_L g578 ( .A(n_508), .Y(n_578) );
AND2x2_ASAP7_75t_L g612 ( .A(n_508), .B(n_560), .Y(n_612) );
AND2x2_ASAP7_75t_L g679 ( .A(n_508), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_509), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g559 ( .A(n_509), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g599 ( .A(n_509), .B(n_521), .Y(n_599) );
AND2x2_ASAP7_75t_L g616 ( .A(n_509), .B(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g542 ( .A(n_521), .B(n_543), .Y(n_542) );
INVx3_ASAP7_75t_L g560 ( .A(n_521), .Y(n_560) );
AND2x2_ASAP7_75t_L g565 ( .A(n_521), .B(n_545), .Y(n_565) );
AND2x2_ASAP7_75t_L g638 ( .A(n_521), .B(n_617), .Y(n_638) );
AND2x2_ASAP7_75t_L g703 ( .A(n_521), .B(n_693), .Y(n_703) );
OAI311xp33_ASAP7_75t_L g586 ( .A1(n_530), .A2(n_587), .A3(n_591), .B1(n_593), .C1(n_613), .Y(n_586) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g598 ( .A(n_531), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g657 ( .A(n_531), .B(n_565), .Y(n_657) );
AND2x2_ASAP7_75t_L g731 ( .A(n_531), .B(n_612), .Y(n_731) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_532), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g666 ( .A(n_532), .Y(n_666) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx3_ASAP7_75t_L g557 ( .A(n_533), .Y(n_557) );
NOR2x1_ASAP7_75t_L g629 ( .A(n_533), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g686 ( .A(n_533), .B(n_560), .Y(n_686) );
AND2x4_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g583 ( .A(n_534), .Y(n_583) );
AND2x2_ASAP7_75t_L g561 ( .A(n_541), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g614 ( .A(n_541), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g694 ( .A(n_541), .B(n_695), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g593 ( .A1(n_542), .A2(n_574), .B1(n_594), .B2(n_598), .C(n_600), .Y(n_593) );
INVx1_ASAP7_75t_L g718 ( .A(n_543), .Y(n_718) );
OR2x2_ASAP7_75t_L g684 ( .A(n_544), .B(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g579 ( .A(n_545), .B(n_560), .Y(n_579) );
OR2x2_ASAP7_75t_L g581 ( .A(n_545), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g606 ( .A(n_545), .Y(n_606) );
INVx2_ASAP7_75t_L g617 ( .A(n_545), .Y(n_617) );
AND2x2_ASAP7_75t_L g644 ( .A(n_545), .B(n_582), .Y(n_644) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_545), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_561), .B1(n_564), .B2(n_567), .C(n_570), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
AND2x2_ASAP7_75t_L g655 ( .A(n_557), .B(n_565), .Y(n_655) );
AND2x2_ASAP7_75t_L g705 ( .A(n_557), .B(n_559), .Y(n_705) );
INVx2_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g592 ( .A(n_559), .B(n_563), .Y(n_592) );
AND2x2_ASAP7_75t_L g671 ( .A(n_559), .B(n_644), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_560), .B(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g630 ( .A(n_560), .Y(n_630) );
OAI21xp33_ASAP7_75t_L g640 ( .A1(n_561), .A2(n_641), .B(n_643), .Y(n_640) );
OR2x2_ASAP7_75t_L g584 ( .A(n_562), .B(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g650 ( .A(n_562), .B(n_610), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_562), .B(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g627 ( .A(n_563), .B(n_596), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_563), .B(n_710), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_564), .B(n_590), .Y(n_700) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
AND2x2_ASAP7_75t_L g623 ( .A(n_565), .B(n_578), .Y(n_623) );
INVx1_ASAP7_75t_L g639 ( .A(n_566), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_576), .B1(n_580), .B2(n_584), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx2_ASAP7_75t_L g602 ( .A(n_573), .Y(n_602) );
INVx1_ASAP7_75t_L g615 ( .A(n_573), .Y(n_615) );
INVx1_ASAP7_75t_L g585 ( .A(n_574), .Y(n_585) );
AND2x2_ASAP7_75t_L g656 ( .A(n_574), .B(n_602), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_574), .B(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
OR2x2_ASAP7_75t_L g580 ( .A(n_577), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_577), .B(n_693), .Y(n_692) );
NOR2xp67_ASAP7_75t_L g724 ( .A(n_577), .B(n_725), .Y(n_724) );
INVx3_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g727 ( .A(n_579), .B(n_679), .Y(n_727) );
INVx1_ASAP7_75t_SL g693 ( .A(n_581), .Y(n_693) );
AND2x2_ASAP7_75t_L g633 ( .A(n_582), .B(n_617), .Y(n_633) );
INVx1_ASAP7_75t_L g680 ( .A(n_582), .Y(n_680) );
OAI222xp33_ASAP7_75t_L g721 ( .A1(n_587), .A2(n_677), .B1(n_722), .B2(n_723), .C1(n_726), .C2(n_728), .Y(n_721) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g642 ( .A(n_589), .Y(n_642) );
AND2x2_ASAP7_75t_L g653 ( .A(n_590), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_590), .B(n_695), .Y(n_722) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_592), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g697 ( .A(n_594), .Y(n_697) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_SL g635 ( .A(n_597), .Y(n_635) );
AND2x2_ASAP7_75t_L g714 ( .A(n_597), .B(n_675), .Y(n_714) );
AND2x2_ASAP7_75t_L g737 ( .A(n_597), .B(n_621), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_599), .B(n_633), .Y(n_632) );
OAI32xp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_603), .A3(n_605), .B1(n_607), .B2(n_611), .Y(n_600) );
BUFx2_ASAP7_75t_L g675 ( .A(n_602), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_603), .B(n_621), .Y(n_702) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g641 ( .A(n_604), .B(n_642), .Y(n_641) );
AND2x4_ASAP7_75t_L g709 ( .A(n_604), .B(n_710), .Y(n_709) );
OR2x2_ASAP7_75t_L g698 ( .A(n_605), .B(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
AND2x2_ASAP7_75t_L g669 ( .A(n_608), .B(n_642), .Y(n_669) );
INVx2_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
OAI221xp5_ASAP7_75t_SL g631 ( .A1(n_610), .A2(n_632), .B1(n_634), .B2(n_636), .C(n_640), .Y(n_631) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g643 ( .A(n_612), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g649 ( .A(n_612), .B(n_633), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_616), .B1(n_618), .B2(n_623), .C(n_624), .Y(n_613) );
INVx1_ASAP7_75t_L g732 ( .A(n_614), .Y(n_732) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_615), .B(n_709), .Y(n_708) );
NAND2x1p5_ASAP7_75t_L g628 ( .A(n_616), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_621), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g687 ( .A(n_621), .Y(n_687) );
BUFx3_ASAP7_75t_L g710 ( .A(n_622), .Y(n_710) );
INVx1_ASAP7_75t_SL g651 ( .A(n_623), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_623), .B(n_665), .Y(n_664) );
AOI21xp33_ASAP7_75t_SL g624 ( .A1(n_625), .A2(n_626), .B(n_628), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g729 ( .A1(n_625), .A2(n_726), .B1(n_730), .B2(n_732), .C(n_733), .Y(n_729) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g672 ( .A(n_630), .B(n_633), .Y(n_672) );
INVx1_ASAP7_75t_L g736 ( .A(n_630), .Y(n_736) );
INVx2_ASAP7_75t_L g725 ( .A(n_633), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_633), .B(n_736), .Y(n_735) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g678 ( .A(n_638), .B(n_679), .Y(n_678) );
OAI221xp5_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_648), .B1(n_650), .B2(n_651), .C(n_652), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_655), .B1(n_656), .B2(n_657), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_654), .A2(n_716), .B1(n_717), .B2(n_719), .Y(n_715) );
OAI21xp5_ASAP7_75t_L g733 ( .A1(n_657), .A2(n_734), .B(n_737), .Y(n_733) );
NOR4xp25_ASAP7_75t_SL g658 ( .A(n_659), .B(n_667), .C(n_676), .D(n_696), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_664), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_670), .B1(n_673), .B2(n_674), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
INVx1_ASAP7_75t_L g712 ( .A(n_672), .Y(n_712) );
OAI221xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_681), .B1(n_684), .B2(n_687), .C(n_688), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g699 ( .A(n_679), .Y(n_699) );
INVx1_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OAI21xp5_ASAP7_75t_SL g688 ( .A1(n_689), .A2(n_691), .B(n_694), .Y(n_688) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI211xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_698), .B(n_700), .C(n_701), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B1(n_704), .B2(n_705), .Y(n_701) );
CKINVDCx14_ASAP7_75t_R g711 ( .A(n_705), .Y(n_711) );
NOR3xp33_ASAP7_75t_L g706 ( .A(n_707), .B(n_721), .C(n_729), .Y(n_706) );
OAI221xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_711), .B1(n_712), .B2(n_713), .C(n_715), .Y(n_707) );
INVxp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
CKINVDCx16_ASAP7_75t_R g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g748 ( .A(n_739), .Y(n_748) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
CKINVDCx16_ASAP7_75t_R g750 ( .A(n_741), .Y(n_750) );
INVx1_ASAP7_75t_L g745 ( .A(n_742), .Y(n_745) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
INVx3_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_755), .Y(n_754) );
endmodule