module fake_jpeg_3332_n_339 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_3),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_52),
.Y(n_136)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_53),
.Y(n_135)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_23),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_56),
.B(n_61),
.Y(n_133)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_65),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_0),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_26),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_66),
.B(n_70),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_37),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_72),
.B(n_80),
.Y(n_142)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_73),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_37),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

BUFx4f_ASAP7_75t_SL g75 ( 
.A(n_26),
.Y(n_75)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_38),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_81),
.B(n_87),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_94),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_38),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_88),
.B(n_89),
.Y(n_149)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_1),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_90),
.B(n_96),
.Y(n_152)
);

BUFx16f_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_91),
.Y(n_129)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_92),
.B(n_30),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_44),
.B(n_2),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_93),
.B(n_99),
.Y(n_157)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_2),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_98),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_28),
.B(n_2),
.Y(n_96)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_97),
.A2(n_33),
.B1(n_34),
.B2(n_42),
.Y(n_103)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_100),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_24),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_102),
.Y(n_145)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g188 ( 
.A(n_103),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_67),
.A2(n_31),
.B1(n_42),
.B2(n_40),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_106),
.A2(n_113),
.B1(n_137),
.B2(n_139),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_64),
.A2(n_49),
.B1(n_41),
.B2(n_39),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_108),
.A2(n_130),
.B1(n_105),
.B2(n_115),
.Y(n_193)
);

NAND3xp33_ASAP7_75t_L g195 ( 
.A(n_111),
.B(n_146),
.C(n_120),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_69),
.A2(n_78),
.B1(n_74),
.B2(n_91),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_54),
.A2(n_30),
.B1(n_40),
.B2(n_35),
.Y(n_121)
);

AO22x1_ASAP7_75t_SL g198 ( 
.A1(n_121),
.A2(n_105),
.B1(n_115),
.B2(n_126),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_68),
.A2(n_35),
.B1(n_32),
.B2(n_31),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_123),
.A2(n_58),
.B1(n_60),
.B2(n_102),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_79),
.A2(n_41),
.B1(n_39),
.B2(n_28),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_138),
.B1(n_140),
.B2(n_143),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_69),
.A2(n_32),
.B1(n_46),
.B2(n_5),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_96),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_77),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_99),
.A2(n_4),
.B1(n_7),
.B2(n_10),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_99),
.A2(n_7),
.B1(n_12),
.B2(n_15),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_90),
.B(n_66),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_71),
.A2(n_89),
.B1(n_101),
.B2(n_100),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_125),
.B1(n_104),
.B2(n_118),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_75),
.B(n_82),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_71),
.Y(n_163)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_158),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_160),
.A2(n_178),
.B1(n_190),
.B2(n_195),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_151),
.B1(n_134),
.B2(n_123),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_181),
.B1(n_193),
.B2(n_198),
.Y(n_200)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_163),
.B(n_168),
.Y(n_221)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

INVx13_ASAP7_75t_L g213 ( 
.A(n_164),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_157),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_142),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_166),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_107),
.B(n_133),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_167),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_132),
.Y(n_168)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_171),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_129),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_172),
.B(n_175),
.Y(n_228)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_180),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_121),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_176),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_122),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_121),
.B(n_109),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_177),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_121),
.B(n_109),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_185),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_122),
.B(n_120),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_117),
.A2(n_148),
.B1(n_116),
.B2(n_153),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_187),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_117),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_183),
.Y(n_227)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_184),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_116),
.B(n_114),
.Y(n_185)
);

INVx13_ASAP7_75t_L g186 ( 
.A(n_124),
.Y(n_186)
);

BUFx12_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_110),
.Y(n_187)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_191),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_148),
.A2(n_127),
.B1(n_130),
.B2(n_153),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_155),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_155),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_192),
.Y(n_209)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_194),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_154),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_196),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_154),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_197),
.B(n_110),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_126),
.B1(n_119),
.B2(n_125),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_202),
.A2(n_219),
.B1(n_200),
.B2(n_220),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_182),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_176),
.B(n_119),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_206),
.B(n_218),
.Y(n_242)
);

AND2x6_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_104),
.Y(n_208)
);

A2O1A1O1Ixp25_ASAP7_75t_L g240 ( 
.A1(n_208),
.A2(n_206),
.B(n_224),
.C(n_228),
.D(n_221),
.Y(n_240)
);

OAI22x1_ASAP7_75t_SL g214 ( 
.A1(n_198),
.A2(n_179),
.B1(n_161),
.B2(n_188),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_214),
.A2(n_220),
.B1(n_190),
.B2(n_188),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_185),
.B(n_171),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_169),
.A2(n_159),
.B1(n_198),
.B2(n_160),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_197),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_230),
.B(n_231),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_212),
.B(n_194),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_232),
.Y(n_272)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_234),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_235),
.A2(n_237),
.B1(n_244),
.B2(n_245),
.Y(n_275)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_236),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_224),
.A2(n_189),
.B1(n_162),
.B2(n_183),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_239),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_192),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_191),
.C(n_187),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_248),
.C(n_253),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_177),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_243),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_200),
.A2(n_170),
.B1(n_173),
.B2(n_184),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_214),
.A2(n_158),
.B1(n_164),
.B2(n_186),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_211),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_246),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_225),
.B(n_201),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_247),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_207),
.B(n_226),
.C(n_204),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_207),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_249),
.Y(n_273)
);

AND2x2_ASAP7_75t_SL g250 ( 
.A(n_208),
.B(n_222),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_250),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_229),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_223),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_209),
.A2(n_199),
.B(n_203),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_210),
.C(n_203),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_227),
.A2(n_223),
.B1(n_217),
.B2(n_205),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_210),
.B(n_217),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_255),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_251),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_234),
.A2(n_205),
.B1(n_213),
.B2(n_216),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_261),
.A2(n_271),
.B1(n_252),
.B2(n_233),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_235),
.A2(n_250),
.B1(n_239),
.B2(n_231),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_267),
.A2(n_270),
.B1(n_232),
.B2(n_254),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_250),
.A2(n_205),
.B1(n_213),
.B2(n_216),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_213),
.B1(n_216),
.B2(n_237),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_246),
.Y(n_276)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_276),
.Y(n_294)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

NAND3xp33_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_247),
.C(n_230),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_279),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_281),
.Y(n_305)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_271),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_282),
.Y(n_297)
);

NAND3xp33_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_242),
.C(n_248),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_265),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_238),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_250),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_289),
.B1(n_291),
.B2(n_292),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_242),
.B(n_240),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_260),
.Y(n_303)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_241),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_272),
.C(n_258),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_266),
.B(n_243),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_290),
.B(n_264),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_302),
.C(n_286),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_282),
.A2(n_274),
.B1(n_267),
.B2(n_268),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_300),
.A2(n_301),
.B1(n_292),
.B2(n_257),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_287),
.A2(n_274),
.B1(n_258),
.B2(n_261),
.Y(n_301)
);

OAI21x1_ASAP7_75t_L g310 ( 
.A1(n_303),
.A2(n_260),
.B(n_272),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_312),
.C(n_313),
.Y(n_321)
);

A2O1A1Ixp33_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_288),
.B(n_280),
.C(n_266),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_305),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_259),
.Y(n_308)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_308),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_309),
.A2(n_293),
.B1(n_297),
.B2(n_305),
.Y(n_316)
);

AO21x1_ASAP7_75t_L g315 ( 
.A1(n_310),
.A2(n_296),
.B(n_300),
.Y(n_315)
);

FAx1_ASAP7_75t_SL g311 ( 
.A(n_302),
.B(n_270),
.CI(n_232),
.CON(n_311),
.SN(n_311)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_298),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_277),
.C(n_281),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_279),
.C(n_289),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_259),
.Y(n_314)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_314),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_315),
.A2(n_319),
.B(n_307),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_318),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_323),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_319),
.A2(n_312),
.B(n_306),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_314),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_325),
.B(n_317),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_313),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_315),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_329),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_320),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_236),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_331),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_298),
.C(n_304),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_333),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_332),
.B(n_329),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_334),
.C(n_304),
.Y(n_337)
);

OAI31xp33_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_311),
.A3(n_216),
.B(n_275),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_311),
.Y(n_339)
);


endmodule