module real_aes_8714_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_504;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g112 ( .A(n_0), .Y(n_112) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_1), .A2(n_129), .B(n_132), .C(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g195 ( .A(n_2), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_3), .A2(n_124), .B(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_4), .B(n_205), .Y(n_519) );
AOI21xp33_ASAP7_75t_L g206 ( .A1(n_5), .A2(n_124), .B(n_207), .Y(n_206) );
AND2x6_ASAP7_75t_L g129 ( .A(n_6), .B(n_130), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_7), .A2(n_175), .B(n_176), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_8), .B(n_41), .Y(n_113) );
INVx1_ASAP7_75t_L g454 ( .A(n_9), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_10), .B(n_165), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_11), .B(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g212 ( .A(n_12), .Y(n_212) );
AOI222xp33_ASAP7_75t_L g114 ( .A1(n_13), .A2(n_19), .B1(n_115), .B2(n_712), .C1(n_713), .C2(n_716), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_13), .Y(n_712) );
INVx1_ASAP7_75t_L g150 ( .A(n_14), .Y(n_150) );
INVx1_ASAP7_75t_L g183 ( .A(n_15), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g462 ( .A1(n_16), .A2(n_138), .B(n_184), .C(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_17), .B(n_205), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_18), .B(n_140), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g123 ( .A(n_20), .B(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_21), .B(n_555), .Y(n_554) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_22), .A2(n_164), .B(n_198), .C(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_23), .B(n_205), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_24), .B(n_165), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_25), .A2(n_180), .B(n_182), .C(n_184), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_26), .B(n_165), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g504 ( .A(n_27), .Y(n_504) );
INVx1_ASAP7_75t_L g493 ( .A(n_28), .Y(n_493) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_29), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_30), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_31), .B(n_165), .Y(n_196) );
INVx1_ASAP7_75t_L g551 ( .A(n_32), .Y(n_551) );
INVx1_ASAP7_75t_L g222 ( .A(n_33), .Y(n_222) );
INVx2_ASAP7_75t_L g127 ( .A(n_34), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_35), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_36), .A2(n_164), .B(n_213), .C(n_517), .Y(n_516) );
INVxp67_ASAP7_75t_L g552 ( .A(n_37), .Y(n_552) );
A2O1A1Ixp33_ASAP7_75t_L g131 ( .A1(n_38), .A2(n_129), .B(n_132), .C(n_135), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_39), .A2(n_132), .B(n_492), .C(n_497), .Y(n_491) );
CKINVDCx14_ASAP7_75t_R g515 ( .A(n_40), .Y(n_515) );
INVx1_ASAP7_75t_L g220 ( .A(n_42), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g452 ( .A1(n_43), .A2(n_142), .B(n_210), .C(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_44), .B(n_165), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_45), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_46), .Y(n_548) );
INVx1_ASAP7_75t_L g482 ( .A(n_47), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g223 ( .A(n_48), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_49), .B(n_124), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_50), .A2(n_132), .B1(n_198), .B2(n_219), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_51), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g191 ( .A(n_52), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_53), .A2(n_210), .B(n_211), .C(n_213), .Y(n_209) );
CKINVDCx14_ASAP7_75t_R g451 ( .A(n_54), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_55), .Y(n_260) );
INVx1_ASAP7_75t_L g208 ( .A(n_56), .Y(n_208) );
INVx1_ASAP7_75t_L g130 ( .A(n_57), .Y(n_130) );
INVx1_ASAP7_75t_L g149 ( .A(n_58), .Y(n_149) );
INVx1_ASAP7_75t_SL g518 ( .A(n_59), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_60), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_61), .B(n_205), .Y(n_486) );
INVx1_ASAP7_75t_L g507 ( .A(n_62), .Y(n_507) );
AOI22xp33_ASAP7_75t_SL g99 ( .A1(n_63), .A2(n_100), .B1(n_727), .B2(n_731), .Y(n_99) );
A2O1A1Ixp33_ASAP7_75t_SL g230 ( .A1(n_64), .A2(n_140), .B(n_213), .C(n_231), .Y(n_230) );
INVxp67_ASAP7_75t_L g232 ( .A(n_65), .Y(n_232) );
INVx1_ASAP7_75t_L g730 ( .A(n_66), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_67), .A2(n_124), .B(n_450), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_68), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_69), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_70), .A2(n_124), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g253 ( .A(n_71), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_72), .A2(n_175), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g461 ( .A(n_73), .Y(n_461) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_74), .Y(n_490) );
OAI22xp5_ASAP7_75t_SL g723 ( .A1(n_75), .A2(n_442), .B1(n_724), .B2(n_725), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_75), .Y(n_725) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_76), .A2(n_129), .B(n_132), .C(n_255), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_77), .A2(n_124), .B(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g464 ( .A(n_78), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_79), .B(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g147 ( .A(n_80), .Y(n_147) );
INVx1_ASAP7_75t_L g473 ( .A(n_81), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_82), .B(n_140), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_83), .A2(n_129), .B(n_132), .C(n_194), .Y(n_193) );
OR2x2_ASAP7_75t_L g109 ( .A(n_84), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g441 ( .A(n_84), .Y(n_441) );
OR2x2_ASAP7_75t_L g711 ( .A(n_84), .B(n_111), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_85), .A2(n_132), .B(n_506), .C(n_509), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_86), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_87), .B(n_158), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_88), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g160 ( .A1(n_89), .A2(n_129), .B(n_132), .C(n_161), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_90), .Y(n_170) );
INVx1_ASAP7_75t_L g229 ( .A(n_91), .Y(n_229) );
CKINVDCx16_ASAP7_75t_R g177 ( .A(n_92), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_93), .B(n_137), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_94), .B(n_154), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_95), .B(n_154), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_96), .A2(n_124), .B(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g485 ( .A(n_97), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_98), .B(n_730), .Y(n_729) );
AOI22x1_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_114), .B1(n_720), .B2(n_722), .Y(n_100) );
NOR2xp33_ASAP7_75t_L g101 ( .A(n_102), .B(n_105), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
BUFx2_ASAP7_75t_L g721 ( .A(n_103), .Y(n_721) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_105), .A2(n_723), .B(n_726), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g726 ( .A(n_108), .Y(n_726) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NOR2x2_ASAP7_75t_L g715 ( .A(n_110), .B(n_441), .Y(n_715) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g440 ( .A(n_111), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
OAI22xp5_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_440), .B1(n_442), .B2(n_711), .Y(n_115) );
INVx2_ASAP7_75t_L g717 ( .A(n_116), .Y(n_717) );
AND2x2_ASAP7_75t_SL g116 ( .A(n_117), .B(n_409), .Y(n_116) );
NOR3xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_302), .C(n_375), .Y(n_117) );
OAI211xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_187), .B(n_234), .C(n_286), .Y(n_118) );
INVxp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_155), .Y(n_120) );
AND2x2_ASAP7_75t_L g250 ( .A(n_121), .B(n_251), .Y(n_250) );
INVx3_ASAP7_75t_L g269 ( .A(n_121), .Y(n_269) );
INVx2_ASAP7_75t_L g284 ( .A(n_121), .Y(n_284) );
INVx1_ASAP7_75t_L g314 ( .A(n_121), .Y(n_314) );
AND2x2_ASAP7_75t_L g364 ( .A(n_121), .B(n_285), .Y(n_364) );
AOI32xp33_ASAP7_75t_L g391 ( .A1(n_121), .A2(n_319), .A3(n_392), .B1(n_394), .B2(n_395), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_121), .B(n_240), .Y(n_397) );
AND2x2_ASAP7_75t_L g424 ( .A(n_121), .B(n_267), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_121), .B(n_433), .Y(n_432) );
OR2x6_ASAP7_75t_L g121 ( .A(n_122), .B(n_151), .Y(n_121) );
AOI21xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_131), .B(n_144), .Y(n_122) );
BUFx2_ASAP7_75t_L g175 ( .A(n_124), .Y(n_175) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_129), .Y(n_124) );
NAND2x1p5_ASAP7_75t_L g192 ( .A(n_125), .B(n_129), .Y(n_192) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_128), .Y(n_125) );
INVx1_ASAP7_75t_L g496 ( .A(n_126), .Y(n_496) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g133 ( .A(n_127), .Y(n_133) );
INVx1_ASAP7_75t_L g199 ( .A(n_127), .Y(n_199) );
INVx1_ASAP7_75t_L g134 ( .A(n_128), .Y(n_134) );
INVx3_ASAP7_75t_L g138 ( .A(n_128), .Y(n_138) );
INVx1_ASAP7_75t_L g140 ( .A(n_128), .Y(n_140) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_128), .Y(n_165) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_128), .Y(n_181) );
INVx4_ASAP7_75t_SL g185 ( .A(n_129), .Y(n_185) );
BUFx3_ASAP7_75t_L g497 ( .A(n_129), .Y(n_497) );
INVx5_ASAP7_75t_L g178 ( .A(n_132), .Y(n_178) );
AND2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
BUFx3_ASAP7_75t_L g143 ( .A(n_133), .Y(n_143) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_133), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_139), .B(n_141), .Y(n_135) );
O2A1O1Ixp33_ASAP7_75t_L g194 ( .A1(n_137), .A2(n_195), .B(n_196), .C(n_197), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_137), .A2(n_493), .B(n_494), .C(n_495), .Y(n_492) );
OAI22xp33_ASAP7_75t_L g550 ( .A1(n_137), .A2(n_180), .B1(n_551), .B2(n_552), .Y(n_550) );
INVx5_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_138), .B(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_138), .B(n_232), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_138), .B(n_454), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_141), .A2(n_256), .B(n_257), .Y(n_255) );
O2A1O1Ixp5_ASAP7_75t_L g472 ( .A1(n_141), .A2(n_473), .B(n_474), .C(n_475), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g506 ( .A1(n_141), .A2(n_474), .B(n_507), .C(n_508), .Y(n_506) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g184 ( .A(n_143), .Y(n_184) );
INVx1_ASAP7_75t_L g258 ( .A(n_144), .Y(n_258) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_145), .A2(n_190), .B(n_200), .Y(n_189) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_145), .A2(n_217), .B(n_224), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_145), .B(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_147), .B(n_148), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
NOR2xp33_ASAP7_75t_SL g151 ( .A(n_152), .B(n_153), .Y(n_151) );
INVx3_ASAP7_75t_L g205 ( .A(n_153), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_153), .B(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_153), .B(n_499), .Y(n_498) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_153), .A2(n_503), .B(n_510), .Y(n_502) );
INVx4_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_154), .A2(n_227), .B(n_233), .Y(n_226) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_154), .Y(n_458) );
AND2x2_ASAP7_75t_L g313 ( .A(n_155), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g335 ( .A(n_155), .Y(n_335) );
AND2x2_ASAP7_75t_L g420 ( .A(n_155), .B(n_250), .Y(n_420) );
AND2x2_ASAP7_75t_L g423 ( .A(n_155), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g155 ( .A(n_156), .B(n_172), .Y(n_155) );
INVx2_ASAP7_75t_L g242 ( .A(n_156), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_156), .B(n_267), .Y(n_273) );
AND2x2_ASAP7_75t_L g283 ( .A(n_156), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g319 ( .A(n_156), .Y(n_319) );
AO21x2_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .B(n_169), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_157), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g555 ( .A(n_157), .Y(n_555) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g171 ( .A(n_158), .Y(n_171) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_158), .A2(n_174), .B(n_186), .Y(n_173) );
OA21x2_ASAP7_75t_L g448 ( .A1(n_158), .A2(n_449), .B(n_455), .Y(n_448) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_158), .A2(n_192), .B(n_490), .C(n_491), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_168), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_166), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_164), .B(n_518), .Y(n_517) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g210 ( .A(n_165), .Y(n_210) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx3_ASAP7_75t_L g213 ( .A(n_167), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_171), .B(n_201), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_171), .B(n_260), .Y(n_259) );
AO21x2_ASAP7_75t_L g468 ( .A1(n_171), .A2(n_469), .B(n_476), .Y(n_468) );
AND2x2_ASAP7_75t_L g261 ( .A(n_172), .B(n_242), .Y(n_261) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g243 ( .A(n_173), .Y(n_243) );
AND2x2_ASAP7_75t_L g285 ( .A(n_173), .B(n_267), .Y(n_285) );
AND2x2_ASAP7_75t_L g354 ( .A(n_173), .B(n_251), .Y(n_354) );
O2A1O1Ixp33_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_179), .C(n_185), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_178), .A2(n_185), .B(n_208), .C(n_209), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_178), .A2(n_185), .B(n_229), .C(n_230), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_SL g450 ( .A1(n_178), .A2(n_185), .B(n_451), .C(n_452), .Y(n_450) );
O2A1O1Ixp33_ASAP7_75t_SL g460 ( .A1(n_178), .A2(n_185), .B(n_461), .C(n_462), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_SL g481 ( .A1(n_178), .A2(n_185), .B(n_482), .C(n_483), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_178), .A2(n_185), .B(n_515), .C(n_516), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_SL g547 ( .A1(n_178), .A2(n_185), .B(n_548), .C(n_549), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_180), .B(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_180), .B(n_464), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_180), .B(n_485), .Y(n_484) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
OAI22xp5_ASAP7_75t_SL g219 ( .A1(n_181), .A2(n_220), .B1(n_221), .B2(n_222), .Y(n_219) );
INVx2_ASAP7_75t_L g221 ( .A(n_181), .Y(n_221) );
OAI22xp33_ASAP7_75t_L g217 ( .A1(n_185), .A2(n_192), .B1(n_218), .B2(n_223), .Y(n_217) );
INVx1_ASAP7_75t_L g509 ( .A(n_185), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_188), .B(n_202), .Y(n_187) );
OR2x2_ASAP7_75t_L g248 ( .A(n_188), .B(n_216), .Y(n_248) );
INVx1_ASAP7_75t_L g327 ( .A(n_188), .Y(n_327) );
AND2x2_ASAP7_75t_L g341 ( .A(n_188), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_188), .B(n_215), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_188), .B(n_339), .Y(n_393) );
AND2x2_ASAP7_75t_L g401 ( .A(n_188), .B(n_402), .Y(n_401) );
INVx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx3_ASAP7_75t_L g238 ( .A(n_189), .Y(n_238) );
AND2x2_ASAP7_75t_L g308 ( .A(n_189), .B(n_216), .Y(n_308) );
OAI21xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_193), .Y(n_190) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_192), .A2(n_253), .B(n_254), .Y(n_252) );
OAI21xp5_ASAP7_75t_L g469 ( .A1(n_192), .A2(n_470), .B(n_471), .Y(n_469) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_192), .A2(n_504), .B(n_505), .Y(n_503) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_202), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g435 ( .A(n_202), .Y(n_435) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_215), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_203), .B(n_279), .Y(n_301) );
OR2x2_ASAP7_75t_L g330 ( .A(n_203), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g362 ( .A(n_203), .B(n_342), .Y(n_362) );
INVx1_ASAP7_75t_SL g382 ( .A(n_203), .Y(n_382) );
AND2x2_ASAP7_75t_L g386 ( .A(n_203), .B(n_247), .Y(n_386) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_SL g239 ( .A(n_204), .B(n_215), .Y(n_239) );
AND2x2_ASAP7_75t_L g246 ( .A(n_204), .B(n_226), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_204), .B(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g289 ( .A(n_204), .B(n_271), .Y(n_289) );
INVx1_ASAP7_75t_SL g296 ( .A(n_204), .Y(n_296) );
BUFx2_ASAP7_75t_L g307 ( .A(n_204), .Y(n_307) );
AND2x2_ASAP7_75t_L g323 ( .A(n_204), .B(n_238), .Y(n_323) );
AND2x2_ASAP7_75t_L g338 ( .A(n_204), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g402 ( .A(n_204), .B(n_216), .Y(n_402) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_214), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_215), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g326 ( .A(n_215), .B(n_327), .Y(n_326) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_215), .A2(n_344), .B1(n_347), .B2(n_350), .C(n_355), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_215), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_226), .Y(n_215) );
INVx3_ASAP7_75t_L g271 ( .A(n_216), .Y(n_271) );
INVx2_ASAP7_75t_L g474 ( .A(n_221), .Y(n_474) );
BUFx2_ASAP7_75t_L g281 ( .A(n_226), .Y(n_281) );
AND2x2_ASAP7_75t_L g295 ( .A(n_226), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g312 ( .A(n_226), .Y(n_312) );
OR2x2_ASAP7_75t_L g331 ( .A(n_226), .B(n_271), .Y(n_331) );
INVx3_ASAP7_75t_L g339 ( .A(n_226), .Y(n_339) );
AND2x2_ASAP7_75t_L g342 ( .A(n_226), .B(n_271), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_240), .B1(n_244), .B2(n_249), .C(n_262), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_239), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_237), .B(n_311), .Y(n_436) );
OR2x2_ASAP7_75t_L g439 ( .A(n_237), .B(n_270), .Y(n_439) );
INVx1_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
OAI221xp5_ASAP7_75t_SL g262 ( .A1(n_238), .A2(n_263), .B1(n_270), .B2(n_272), .C(n_275), .Y(n_262) );
AND2x2_ASAP7_75t_L g279 ( .A(n_238), .B(n_271), .Y(n_279) );
AND2x2_ASAP7_75t_L g287 ( .A(n_238), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_238), .B(n_295), .Y(n_294) );
NAND2x1_ASAP7_75t_L g337 ( .A(n_238), .B(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g389 ( .A(n_238), .B(n_331), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_240), .A2(n_349), .B1(n_378), .B2(n_380), .Y(n_377) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AOI322xp5_ASAP7_75t_L g286 ( .A1(n_241), .A2(n_250), .A3(n_287), .B1(n_290), .B2(n_293), .C1(n_297), .C2(n_300), .Y(n_286) );
OR2x2_ASAP7_75t_L g298 ( .A(n_241), .B(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_242), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g277 ( .A(n_242), .B(n_251), .Y(n_277) );
INVx1_ASAP7_75t_L g292 ( .A(n_242), .Y(n_292) );
AND2x2_ASAP7_75t_L g358 ( .A(n_242), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g268 ( .A(n_243), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g359 ( .A(n_243), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_243), .B(n_267), .Y(n_433) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_247), .B(n_382), .Y(n_381) );
INVx3_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g333 ( .A(n_248), .B(n_280), .Y(n_333) );
OR2x2_ASAP7_75t_L g430 ( .A(n_248), .B(n_281), .Y(n_430) );
INVx1_ASAP7_75t_L g411 ( .A(n_249), .Y(n_411) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_261), .Y(n_249) );
INVx4_ASAP7_75t_L g299 ( .A(n_250), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_250), .B(n_318), .Y(n_324) );
INVx2_ASAP7_75t_L g267 ( .A(n_251), .Y(n_267) );
AO21x2_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_258), .B(n_259), .Y(n_251) );
AO21x2_ASAP7_75t_L g544 ( .A1(n_258), .A2(n_545), .B(n_553), .Y(n_544) );
INVx1_ASAP7_75t_L g562 ( .A(n_258), .Y(n_562) );
INVx1_ASAP7_75t_L g349 ( .A(n_261), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_261), .B(n_321), .Y(n_390) );
AOI21xp33_ASAP7_75t_L g336 ( .A1(n_263), .A2(n_337), .B(n_340), .Y(n_336) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_268), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g321 ( .A(n_267), .Y(n_321) );
INVx1_ASAP7_75t_L g348 ( .A(n_267), .Y(n_348) );
INVx1_ASAP7_75t_L g274 ( .A(n_268), .Y(n_274) );
AND2x2_ASAP7_75t_L g276 ( .A(n_268), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g372 ( .A(n_269), .B(n_358), .Y(n_372) );
AND2x2_ASAP7_75t_L g394 ( .A(n_269), .B(n_354), .Y(n_394) );
BUFx2_ASAP7_75t_L g346 ( .A(n_271), .Y(n_346) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
AOI32xp33_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_278), .A3(n_279), .B1(n_280), .B2(n_282), .Y(n_275) );
INVx1_ASAP7_75t_L g356 ( .A(n_276), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_276), .A2(n_404), .B1(n_405), .B2(n_407), .Y(n_403) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_279), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_279), .B(n_338), .Y(n_379) );
AND2x2_ASAP7_75t_L g426 ( .A(n_279), .B(n_311), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_280), .B(n_327), .Y(n_374) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g427 ( .A(n_282), .Y(n_427) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVx1_ASAP7_75t_L g352 ( .A(n_283), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_285), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g399 ( .A(n_285), .B(n_319), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_285), .B(n_314), .Y(n_406) );
INVx1_ASAP7_75t_SL g388 ( .A(n_287), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_288), .B(n_339), .Y(n_366) );
NOR4xp25_ASAP7_75t_L g412 ( .A(n_288), .B(n_311), .C(n_413), .D(n_416), .Y(n_412) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_289), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVxp67_ASAP7_75t_L g369 ( .A(n_292), .Y(n_369) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OAI21xp33_ASAP7_75t_L g419 ( .A1(n_295), .A2(n_386), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g311 ( .A(n_296), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g360 ( .A(n_299), .Y(n_360) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND4xp25_ASAP7_75t_SL g302 ( .A(n_303), .B(n_328), .C(n_343), .D(n_363), .Y(n_302) );
O2A1O1Ixp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_309), .B(n_313), .C(n_315), .Y(n_303) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g395 ( .A(n_308), .B(n_338), .Y(n_395) );
AND2x2_ASAP7_75t_L g404 ( .A(n_308), .B(n_382), .Y(n_404) );
INVx3_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_311), .B(n_346), .Y(n_408) );
AND2x2_ASAP7_75t_L g320 ( .A(n_314), .B(n_321), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_322), .B1(n_324), .B2(n_325), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
AND2x2_ASAP7_75t_L g418 ( .A(n_318), .B(n_364), .Y(n_418) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_320), .B(n_369), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_321), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_332), .B(n_334), .C(n_336), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_329), .A2(n_364), .B1(n_365), .B2(n_367), .C(n_370), .Y(n_363) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OAI221xp5_ASAP7_75t_L g421 ( .A1(n_337), .A2(n_422), .B1(n_425), .B2(n_427), .C(n_428), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_338), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_346), .B(n_415), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx1_ASAP7_75t_L g376 ( .A(n_348), .Y(n_376) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_351), .A2(n_371), .B1(n_373), .B2(n_374), .Y(n_370) );
OR2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AOI21xp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_357), .B(n_361), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_360), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g434 ( .A1(n_371), .A2(n_397), .B1(n_435), .B2(n_436), .C(n_437), .Y(n_434) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g416 ( .A(n_373), .Y(n_416) );
OAI211xp5_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_377), .B(n_383), .C(n_403), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI211xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_386), .B(n_387), .C(n_396), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
A2O1A1Ixp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B(n_390), .C(n_391), .Y(n_387) );
INVx1_ASAP7_75t_L g415 ( .A(n_393), .Y(n_415) );
OAI21xp5_ASAP7_75t_SL g437 ( .A1(n_394), .A2(n_420), .B(n_438), .Y(n_437) );
AOI21xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B(n_400), .Y(n_396) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI21xp5_ASAP7_75t_SL g429 ( .A1(n_406), .A2(n_430), .B(n_431), .Y(n_429) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NOR3xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_421), .C(n_434), .Y(n_409) );
OAI211xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B(n_417), .C(n_419), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
CKINVDCx14_ASAP7_75t_R g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g719 ( .A(n_440), .Y(n_719) );
INVx1_ASAP7_75t_L g724 ( .A(n_442), .Y(n_724) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI22xp5_ASAP7_75t_SL g716 ( .A1(n_443), .A2(n_711), .B1(n_717), .B2(n_718), .Y(n_716) );
OR2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_641), .Y(n_443) );
NAND5xp2_ASAP7_75t_L g444 ( .A(n_445), .B(n_556), .C(n_588), .D(n_605), .E(n_628), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_487), .B1(n_520), .B2(n_524), .C(n_528), .Y(n_445) );
INVx1_ASAP7_75t_L g668 ( .A(n_446), .Y(n_668) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_466), .Y(n_446) );
AND3x2_ASAP7_75t_L g643 ( .A(n_447), .B(n_468), .C(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_456), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_448), .B(n_526), .Y(n_525) );
BUFx3_ASAP7_75t_L g535 ( .A(n_448), .Y(n_535) );
AND2x2_ASAP7_75t_L g539 ( .A(n_448), .B(n_478), .Y(n_539) );
INVx2_ASAP7_75t_L g565 ( .A(n_448), .Y(n_565) );
OR2x2_ASAP7_75t_L g576 ( .A(n_448), .B(n_479), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_448), .B(n_467), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_448), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g655 ( .A(n_448), .B(n_479), .Y(n_655) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_456), .Y(n_538) );
AND2x2_ASAP7_75t_L g596 ( .A(n_456), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_456), .B(n_467), .Y(n_615) );
INVx1_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g527 ( .A(n_457), .B(n_467), .Y(n_527) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_457), .Y(n_534) );
AND2x2_ASAP7_75t_L g582 ( .A(n_457), .B(n_479), .Y(n_582) );
NAND3xp33_ASAP7_75t_L g607 ( .A(n_457), .B(n_466), .C(n_565), .Y(n_607) );
AND2x2_ASAP7_75t_L g672 ( .A(n_457), .B(n_468), .Y(n_672) );
AND2x2_ASAP7_75t_L g706 ( .A(n_457), .B(n_467), .Y(n_706) );
OA21x2_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_459), .B(n_465), .Y(n_457) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_458), .A2(n_480), .B(n_486), .Y(n_479) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_458), .A2(n_513), .B(n_519), .Y(n_512) );
INVxp67_ASAP7_75t_L g536 ( .A(n_466), .Y(n_536) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_478), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_467), .B(n_565), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_467), .B(n_596), .Y(n_604) );
AND2x2_ASAP7_75t_L g654 ( .A(n_467), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g682 ( .A(n_467), .Y(n_682) );
INVx4_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g589 ( .A(n_468), .B(n_582), .Y(n_589) );
BUFx3_ASAP7_75t_L g621 ( .A(n_468), .Y(n_621) );
INVx2_ASAP7_75t_L g597 ( .A(n_478), .Y(n_597) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_479), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_487), .A2(n_657), .B1(n_659), .B2(n_660), .Y(n_656) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_500), .Y(n_487) );
AND2x2_ASAP7_75t_L g520 ( .A(n_488), .B(n_521), .Y(n_520) );
INVx3_ASAP7_75t_SL g531 ( .A(n_488), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_488), .B(n_560), .Y(n_592) );
OR2x2_ASAP7_75t_L g611 ( .A(n_488), .B(n_501), .Y(n_611) );
AND2x2_ASAP7_75t_L g616 ( .A(n_488), .B(n_568), .Y(n_616) );
AND2x2_ASAP7_75t_L g619 ( .A(n_488), .B(n_561), .Y(n_619) );
AND2x2_ASAP7_75t_L g631 ( .A(n_488), .B(n_512), .Y(n_631) );
AND2x2_ASAP7_75t_L g647 ( .A(n_488), .B(n_502), .Y(n_647) );
AND2x4_ASAP7_75t_L g650 ( .A(n_488), .B(n_522), .Y(n_650) );
OR2x2_ASAP7_75t_L g667 ( .A(n_488), .B(n_603), .Y(n_667) );
OR2x2_ASAP7_75t_L g698 ( .A(n_488), .B(n_544), .Y(n_698) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_488), .B(n_626), .Y(n_700) );
OR2x6_ASAP7_75t_L g488 ( .A(n_489), .B(n_498), .Y(n_488) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_496), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g574 ( .A(n_500), .B(n_542), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_500), .B(n_561), .Y(n_693) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_512), .Y(n_500) );
AND2x2_ASAP7_75t_L g530 ( .A(n_501), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g560 ( .A(n_501), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g568 ( .A(n_501), .B(n_544), .Y(n_568) );
AND2x2_ASAP7_75t_L g586 ( .A(n_501), .B(n_522), .Y(n_586) );
OR2x2_ASAP7_75t_L g603 ( .A(n_501), .B(n_561), .Y(n_603) );
INVx2_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
BUFx2_ASAP7_75t_L g523 ( .A(n_502), .Y(n_523) );
AND2x2_ASAP7_75t_L g626 ( .A(n_502), .B(n_512), .Y(n_626) );
INVx2_ASAP7_75t_L g522 ( .A(n_512), .Y(n_522) );
INVx1_ASAP7_75t_L g638 ( .A(n_512), .Y(n_638) );
AND2x2_ASAP7_75t_L g688 ( .A(n_512), .B(n_531), .Y(n_688) );
AND2x2_ASAP7_75t_L g541 ( .A(n_521), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g572 ( .A(n_521), .B(n_531), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_521), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
AND2x2_ASAP7_75t_L g559 ( .A(n_522), .B(n_531), .Y(n_559) );
OR2x2_ASAP7_75t_L g675 ( .A(n_523), .B(n_649), .Y(n_675) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_526), .B(n_655), .Y(n_661) );
INVx2_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
OAI32xp33_ASAP7_75t_L g617 ( .A1(n_527), .A2(n_618), .A3(n_620), .B1(n_622), .B2(n_623), .Y(n_617) );
OR2x2_ASAP7_75t_L g634 ( .A(n_527), .B(n_576), .Y(n_634) );
OAI21xp33_ASAP7_75t_SL g659 ( .A1(n_527), .A2(n_537), .B(n_564), .Y(n_659) );
OAI22xp33_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_532), .B1(n_537), .B2(n_540), .Y(n_528) );
INVxp33_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_530), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_531), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g585 ( .A(n_531), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g685 ( .A(n_531), .B(n_626), .Y(n_685) );
OR2x2_ASAP7_75t_L g709 ( .A(n_531), .B(n_603), .Y(n_709) );
AOI21xp33_ASAP7_75t_L g692 ( .A1(n_532), .A2(n_591), .B(n_693), .Y(n_692) );
OR2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_536), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g569 ( .A(n_534), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_534), .B(n_539), .Y(n_587) );
AND2x2_ASAP7_75t_L g609 ( .A(n_535), .B(n_582), .Y(n_609) );
INVx1_ASAP7_75t_L g622 ( .A(n_535), .Y(n_622) );
OR2x2_ASAP7_75t_L g627 ( .A(n_535), .B(n_561), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_538), .B(n_576), .Y(n_575) );
OAI22xp33_ASAP7_75t_L g557 ( .A1(n_539), .A2(n_558), .B1(n_563), .B2(n_567), .Y(n_557) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_542), .A2(n_600), .B1(n_607), .B2(n_608), .Y(n_606) );
AND2x2_ASAP7_75t_L g684 ( .A(n_542), .B(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_544), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g703 ( .A(n_544), .B(n_586), .Y(n_703) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OA21x2_ASAP7_75t_L g561 ( .A1(n_546), .A2(n_554), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AOI221xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_569), .B1(n_570), .B2(n_575), .C(n_577), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_559), .B(n_561), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_559), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g578 ( .A(n_560), .Y(n_578) );
O2A1O1Ixp33_ASAP7_75t_L g665 ( .A1(n_560), .A2(n_666), .B(n_667), .C(n_668), .Y(n_665) );
AND2x2_ASAP7_75t_L g670 ( .A(n_560), .B(n_650), .Y(n_670) );
O2A1O1Ixp33_ASAP7_75t_SL g708 ( .A1(n_560), .A2(n_649), .B(n_709), .C(n_710), .Y(n_708) );
BUFx3_ASAP7_75t_L g600 ( .A(n_561), .Y(n_600) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_564), .B(n_621), .Y(n_664) );
AOI211xp5_ASAP7_75t_L g683 ( .A1(n_564), .A2(n_684), .B(n_686), .C(n_692), .Y(n_683) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
INVxp67_ASAP7_75t_L g644 ( .A(n_566), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_568), .B(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_571), .B(n_573), .Y(n_570) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
AOI211xp5_ASAP7_75t_L g588 ( .A1(n_572), .A2(n_589), .B(n_590), .C(n_598), .Y(n_588) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g673 ( .A(n_576), .Y(n_673) );
OR2x2_ASAP7_75t_L g690 ( .A(n_576), .B(n_620), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_579), .B1(n_584), .B2(n_587), .Y(n_577) );
OAI22xp33_ASAP7_75t_L g590 ( .A1(n_579), .A2(n_591), .B1(n_592), .B2(n_593), .Y(n_590) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
OR2x2_ASAP7_75t_L g677 ( .A(n_581), .B(n_621), .Y(n_677) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g632 ( .A(n_582), .B(n_622), .Y(n_632) );
INVx1_ASAP7_75t_L g640 ( .A(n_583), .Y(n_640) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_586), .B(n_600), .Y(n_648) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_596), .B(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g705 ( .A(n_597), .Y(n_705) );
AOI21xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_601), .B(n_604), .Y(n_598) );
INVx1_ASAP7_75t_L g635 ( .A(n_599), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_600), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_600), .B(n_631), .Y(n_630) );
NAND2x1p5_ASAP7_75t_L g651 ( .A(n_600), .B(n_626), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_600), .B(n_647), .Y(n_658) );
OAI211xp5_ASAP7_75t_L g662 ( .A1(n_600), .A2(n_610), .B(n_650), .C(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
AOI221xp5_ASAP7_75t_SL g605 ( .A1(n_606), .A2(n_610), .B1(n_612), .B2(n_616), .C(n_617), .Y(n_605) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVxp67_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_614), .B(n_622), .Y(n_696) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_L g707 ( .A1(n_616), .A2(n_631), .B(n_633), .C(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_619), .B(n_626), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_620), .B(n_673), .Y(n_710) );
CKINVDCx16_ASAP7_75t_R g620 ( .A(n_621), .Y(n_620) );
INVxp33_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
AOI21xp33_ASAP7_75t_SL g636 ( .A1(n_625), .A2(n_637), .B(n_639), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_625), .B(n_698), .Y(n_697) );
INVx2_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_626), .B(n_680), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_632), .B1(n_633), .B2(n_635), .C(n_636), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_632), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g666 ( .A(n_638), .Y(n_666) );
NAND5xp2_ASAP7_75t_L g641 ( .A(n_642), .B(n_669), .C(n_683), .D(n_694), .E(n_707), .Y(n_641) );
AOI211xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B(n_652), .C(n_665), .Y(n_642) );
INVx2_ASAP7_75t_SL g689 ( .A(n_643), .Y(n_689) );
NAND4xp25_ASAP7_75t_SL g645 ( .A(n_646), .B(n_648), .C(n_649), .D(n_651), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx3_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI211xp5_ASAP7_75t_SL g652 ( .A1(n_651), .A2(n_653), .B(n_656), .C(n_662), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_654), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_654), .A2(n_695), .B1(n_697), .B2(n_699), .C(n_701), .Y(n_694) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AOI221xp5_ASAP7_75t_SL g669 ( .A1(n_670), .A2(n_671), .B1(n_674), .B2(n_676), .C(n_678), .Y(n_669) );
AND2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_677), .A2(n_700), .B1(n_702), .B2(n_704), .Y(n_701) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .B1(n_690), .B2(n_691), .Y(n_686) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g728 ( .A(n_714), .B(n_729), .Y(n_728) );
INVx3_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g732 ( .A(n_728), .Y(n_732) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
endmodule