module fake_jpeg_5667_n_302 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_247;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_273;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_35),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_41),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_15),
.B1(n_30),
.B2(n_22),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_42),
.A2(n_43),
.B1(n_45),
.B2(n_47),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_15),
.B(n_26),
.Y(n_43)
);

OA22x2_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_15),
.B1(n_30),
.B2(n_26),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_48),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_30),
.B1(n_19),
.B2(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_32),
.A2(n_25),
.B1(n_18),
.B2(n_21),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_33),
.B1(n_38),
.B2(n_41),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_32),
.A2(n_19),
.B1(n_18),
.B2(n_27),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_59),
.B1(n_42),
.B2(n_45),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_33),
.A2(n_27),
.B1(n_28),
.B2(n_26),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_28),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_63),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_14),
.B(n_13),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_67),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_26),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_68),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_69),
.B(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_40),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_72),
.A2(n_81),
.B1(n_58),
.B2(n_49),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_73),
.B(n_84),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

CKINVDCx6p67_ASAP7_75t_R g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx4f_ASAP7_75t_SL g86 ( 
.A(n_76),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_80),
.B1(n_58),
.B2(n_49),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_0),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_78),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_38),
.B1(n_33),
.B2(n_41),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

AND2x4_ASAP7_75t_SL g85 ( 
.A(n_67),
.B(n_45),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_85),
.A2(n_89),
.B(n_95),
.Y(n_125)
);

CKINVDCx9p33_ASAP7_75t_R g87 ( 
.A(n_76),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_100),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_45),
.C(n_56),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_103),
.C(n_80),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_53),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_72),
.A2(n_58),
.B1(n_60),
.B2(n_46),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_98),
.B1(n_81),
.B2(n_77),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_57),
.B(n_56),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_81),
.B1(n_65),
.B2(n_82),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_55),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_79),
.A2(n_51),
.B(n_52),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_101),
.B(n_80),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_46),
.C(n_62),
.Y(n_103)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_54),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_49),
.B1(n_82),
.B2(n_76),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_74),
.B1(n_96),
.B2(n_105),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_108),
.B(n_85),
.Y(n_134)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_112),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_103),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_88),
.C(n_103),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_115),
.A2(n_118),
.B(n_119),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_98),
.B1(n_93),
.B2(n_101),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_95),
.B(n_96),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_77),
.C(n_65),
.Y(n_118)
);

AO22x1_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_76),
.B1(n_36),
.B2(n_62),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_120),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_69),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_122),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_86),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_123),
.B(n_130),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_71),
.Y(n_124)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_102),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_126),
.Y(n_144)
);

MAJx2_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_74),
.C(n_70),
.Y(n_127)
);

XOR2x2_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_100),
.Y(n_149)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_70),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_109),
.B(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_91),
.C(n_36),
.Y(n_181)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_130),
.A2(n_85),
.B1(n_101),
.B2(n_89),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_119),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_139),
.A2(n_152),
.B1(n_92),
.B2(n_128),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_140),
.A2(n_145),
.B(n_146),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_125),
.B(n_121),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_124),
.B(n_108),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_129),
.Y(n_161)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_150),
.B(n_153),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_119),
.A2(n_113),
.B1(n_107),
.B2(n_118),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_108),
.A2(n_105),
.B(n_100),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_155),
.B(n_86),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_115),
.C(n_111),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_158),
.C(n_160),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_150),
.A2(n_118),
.B1(n_119),
.B2(n_115),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_157),
.A2(n_173),
.B1(n_137),
.B2(n_142),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_159),
.A2(n_163),
.B(n_155),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_127),
.C(n_126),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_176),
.Y(n_185)
);

OA21x2_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_86),
.B(n_123),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_78),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_165),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_112),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_166),
.B(n_153),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_102),
.C(n_86),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_181),
.C(n_36),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_104),
.Y(n_169)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_144),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_172),
.Y(n_197)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_149),
.A2(n_75),
.B1(n_82),
.B2(n_86),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_179),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_104),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_175),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_131),
.B(n_114),
.Y(n_176)
);

BUFx12_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_178),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_83),
.B1(n_68),
.B2(n_37),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_167),
.A2(n_132),
.B1(n_139),
.B2(n_140),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_183),
.A2(n_192),
.B1(n_194),
.B2(n_196),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_145),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_188),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_154),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_136),
.B(n_143),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_173),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_152),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_191),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_135),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_143),
.B(n_133),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_177),
.A2(n_141),
.B1(n_148),
.B2(n_137),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_SL g198 ( 
.A(n_164),
.B(n_148),
.C(n_142),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_204),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_205),
.C(n_181),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_166),
.A2(n_122),
.B1(n_83),
.B2(n_68),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_157),
.B(n_62),
.C(n_37),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_206),
.A2(n_210),
.B(n_211),
.Y(n_230)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_193),
.Y(n_209)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_170),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_170),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_165),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_217),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_192),
.A2(n_163),
.B1(n_178),
.B2(n_168),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_219),
.B(n_221),
.Y(n_237)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_176),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_163),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_222),
.A2(n_225),
.B(n_226),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_191),
.A2(n_205),
.B1(n_188),
.B2(n_200),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_223),
.A2(n_214),
.B1(n_220),
.B2(n_224),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_195),
.C(n_202),
.Y(n_231)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

A2O1A1O1Ixp25_ASAP7_75t_L g226 ( 
.A1(n_185),
.A2(n_178),
.B(n_37),
.C(n_87),
.D(n_26),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_187),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_233),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_232),
.C(n_235),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_195),
.C(n_17),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_23),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_236),
.C(n_240),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_17),
.C(n_23),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_23),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_220),
.A2(n_17),
.B1(n_13),
.B2(n_2),
.Y(n_238)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_1),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_23),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_17),
.C(n_23),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_232),
.C(n_235),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_207),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_242)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_218),
.Y(n_248)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_242),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_249),
.A2(n_253),
.B(n_259),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_250),
.A2(n_257),
.B(n_3),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_0),
.Y(n_251)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_0),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_252),
.B(n_2),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_1),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_256),
.A2(n_260),
.B(n_261),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_16),
.C(n_3),
.Y(n_257)
);

NOR2x1p5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_16),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_236),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_262),
.A2(n_270),
.B(n_272),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_10),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_254),
.A2(n_231),
.B1(n_229),
.B2(n_234),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_275),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_227),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_273),
.Y(n_280)
);

NOR2x1_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_3),
.Y(n_269)
);

FAx1_ASAP7_75t_SL g278 ( 
.A(n_269),
.B(n_257),
.CI(n_247),
.CON(n_278),
.SN(n_278)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_258),
.B(n_16),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_246),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_246),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_274),
.B(n_4),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_250),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_269),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_278),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

AOI322xp5_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_264),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_6),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_5),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_283),
.A2(n_284),
.B(n_285),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_5),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_266),
.B(n_5),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_6),
.C(n_7),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_275),
.C(n_266),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_277),
.A2(n_267),
.B(n_273),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_291),
.C(n_292),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_285),
.B(n_280),
.Y(n_292)
);

AOI21x1_ASAP7_75t_L g295 ( 
.A1(n_293),
.A2(n_6),
.B(n_7),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_289),
.A2(n_278),
.B1(n_7),
.B2(n_9),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_295),
.Y(n_299)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

AO21x1_ASAP7_75t_L g300 ( 
.A1(n_296),
.A2(n_298),
.B(n_9),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_290),
.A2(n_9),
.B(n_287),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_297),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_299),
.Y(n_302)
);


endmodule