module real_jpeg_27857_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_191;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

INVx5_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_0),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_1),
.A2(n_79),
.B1(n_84),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_1),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_1),
.A2(n_49),
.B1(n_50),
.B2(n_134),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_1),
.A2(n_27),
.B1(n_30),
.B2(n_134),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_1),
.A2(n_33),
.B1(n_36),
.B2(n_134),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_2),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_2),
.B(n_82),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_2),
.B(n_49),
.Y(n_190)
);

AOI21xp33_ASAP7_75t_L g194 ( 
.A1(n_2),
.A2(n_49),
.B(n_190),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_152),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_2),
.A2(n_33),
.B(n_37),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_2),
.B(n_100),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_2),
.A2(n_63),
.B1(n_66),
.B2(n_238),
.Y(n_241)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_4),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_4),
.A2(n_27),
.B1(n_30),
.B2(n_58),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_4),
.A2(n_33),
.B1(n_36),
.B2(n_58),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_6),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_7),
.A2(n_27),
.B1(n_30),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_7),
.A2(n_43),
.B1(n_79),
.B2(n_84),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_7),
.A2(n_33),
.B1(n_36),
.B2(n_43),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_7),
.A2(n_43),
.B1(n_49),
.B2(n_50),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_8),
.A2(n_79),
.B1(n_84),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_8),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_8),
.A2(n_49),
.B1(n_50),
.B2(n_107),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_8),
.A2(n_27),
.B1(n_30),
.B2(n_107),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_8),
.A2(n_33),
.B1(n_36),
.B2(n_107),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_9),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_9),
.A2(n_29),
.B1(n_33),
.B2(n_36),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_9),
.A2(n_29),
.B1(n_79),
.B2(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_9),
.A2(n_29),
.B1(n_49),
.B2(n_50),
.Y(n_129)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_11),
.A2(n_49),
.B1(n_50),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_11),
.A2(n_27),
.B1(n_30),
.B2(n_56),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_11),
.A2(n_33),
.B1(n_36),
.B2(n_56),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_12),
.A2(n_79),
.B1(n_84),
.B2(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_12),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_154),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_12),
.A2(n_27),
.B1(n_30),
.B2(n_154),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_12),
.A2(n_33),
.B1(n_36),
.B2(n_154),
.Y(n_238)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_14),
.A2(n_27),
.B1(n_30),
.B2(n_53),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_15),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_136),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_135),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_110),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_20),
.B(n_110),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_89),
.B2(n_109),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_60),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_44),
.B(n_59),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_25),
.A2(n_40),
.B(n_198),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_26),
.Y(n_145)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_27),
.A2(n_30),
.B1(n_35),
.B2(n_37),
.Y(n_41)
);

NAND2xp33_ASAP7_75t_SL g191 ( 
.A(n_27),
.B(n_47),
.Y(n_191)
);

A2O1A1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_27),
.A2(n_35),
.B(n_152),
.C(n_217),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g189 ( 
.A1(n_30),
.A2(n_50),
.A3(n_53),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_31),
.B(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_32),
.A2(n_40),
.B1(n_71),
.B2(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_32),
.A2(n_38),
.B(n_98),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_32),
.A2(n_40),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_32),
.A2(n_40),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_32),
.A2(n_40),
.B1(n_197),
.B2(n_215),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_32),
.B(n_152),
.Y(n_236)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_33),
.Y(n_36)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_36),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_40),
.A2(n_71),
.B(n_72),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_40),
.A2(n_72),
.B(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_52),
.B1(n_54),
.B2(n_57),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_45),
.B(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_45),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_45),
.A2(n_52),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_45),
.A2(n_52),
.B1(n_148),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_45),
.A2(n_52),
.B1(n_177),
.B2(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_46)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_50),
.B1(n_77),
.B2(n_78),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_49),
.B(n_77),
.Y(n_166)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_50),
.A2(n_81),
.B1(n_151),
.B2(n_166),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_52),
.B(n_102),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_52),
.B(n_129),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_55),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_73),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_70),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_62),
.A2(n_74),
.B1(n_75),
.B2(n_88),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_62),
.A2(n_70),
.B1(n_88),
.B2(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_67),
.B(n_68),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_63),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_63),
.A2(n_66),
.B1(n_120),
.B2(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_63),
.A2(n_95),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_63),
.A2(n_230),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_64),
.A2(n_69),
.B(n_122),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_64),
.A2(n_96),
.B1(n_229),
.B2(n_231),
.Y(n_228)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_67),
.A2(n_92),
.B(n_168),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_67),
.B(n_152),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_70),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_83),
.B(n_85),
.Y(n_75)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_76),
.A2(n_82),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_79),
.B(n_81),
.C(n_82),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_79),
.Y(n_81)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

HAxp5_ASAP7_75t_SL g151 ( 
.A(n_79),
.B(n_152),
.CON(n_151),
.SN(n_151)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_82),
.B(n_83),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_86),
.A2(n_105),
.B1(n_106),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_86),
.A2(n_105),
.B1(n_133),
.B2(n_159),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_99),
.C(n_103),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_91),
.B(n_97),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_123),
.Y(n_122)
);

INVx11_ASAP7_75t_L g239 ( 
.A(n_96),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_99),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B(n_108),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.C(n_117),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_115),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_117),
.B(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_126),
.C(n_131),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_118),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_125),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_125),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_126),
.A2(n_131),
.B1(n_132),
.B2(n_272),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_126),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B(n_130),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_127),
.A2(n_162),
.B(n_163),
.Y(n_161)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_276),
.B(n_281),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_181),
.B(n_262),
.C(n_275),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_169),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_139),
.B(n_169),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_155),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_141),
.B(n_142),
.C(n_155),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.C(n_150),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_150),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_164),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_160),
.B2(n_161),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_157),
.B(n_161),
.C(n_164),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_167),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.C(n_175),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_170),
.A2(n_171),
.B1(n_257),
.B2(n_259),
.Y(n_256)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_175),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_180),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_180),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_261),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_254),
.B(n_260),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_208),
.B(n_253),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_199),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_185),
.B(n_199),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_192),
.C(n_195),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_186),
.A2(n_187),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_189),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_192),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_204),
.B2(n_205),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_200),
.B(n_206),
.C(n_207),
.Y(n_255)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_247),
.B(n_252),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_226),
.B(n_246),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_218),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_211),
.B(n_218),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_216),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_212),
.A2(n_213),
.B1(n_216),
.B2(n_233),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_224),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_223),
.C(n_224),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_225),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_234),
.B(n_245),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_232),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_228),
.B(n_232),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_240),
.B(n_244),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_236),
.B(n_237),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_248),
.B(n_249),
.Y(n_252)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_255),
.B(n_256),
.Y(n_260)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_257),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_263),
.B(n_264),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_273),
.B2(n_274),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_270),
.C(n_274),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_273),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_277),
.B(n_278),
.Y(n_281)
);


endmodule