module fake_jpeg_25129_n_272 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_38;
wire n_26;
wire n_28;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx11_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_33),
.Y(n_52)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_44),
.Y(n_60)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_33),
.B1(n_19),
.B2(n_26),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_63),
.B1(n_66),
.B2(n_35),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_19),
.B1(n_33),
.B2(n_26),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_61),
.B1(n_64),
.B2(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_27),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_56),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_24),
.Y(n_56)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_17),
.B1(n_21),
.B2(n_32),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_38),
.A2(n_27),
.B1(n_25),
.B2(n_21),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_22),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_17),
.B1(n_21),
.B2(n_31),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_69),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_31),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_71),
.Y(n_89)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_41),
.B1(n_38),
.B2(n_17),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_72),
.A2(n_75),
.B1(n_81),
.B2(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_52),
.B(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_83),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_18),
.B(n_29),
.Y(n_100)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_78),
.Y(n_108)
);

NOR2x1_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_35),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_93),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_46),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_87),
.C(n_45),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_38),
.B1(n_41),
.B2(n_20),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_84),
.B(n_85),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_55),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_51),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_86),
.B(n_91),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_42),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_36),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_94),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_51),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_62),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_39),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_55),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_68),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_58),
.B(n_18),
.C(n_29),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_112),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_67),
.B1(n_71),
.B2(n_41),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_78),
.B1(n_93),
.B2(n_86),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_79),
.B1(n_80),
.B2(n_73),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_101),
.B1(n_110),
.B2(n_120),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_87),
.B1(n_78),
.B2(n_91),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_58),
.B1(n_70),
.B2(n_57),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_102),
.B(n_117),
.Y(n_139)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_116),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_106),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_76),
.A2(n_57),
.B1(n_48),
.B2(n_42),
.Y(n_110)
);

BUFx12_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_111),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_46),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_46),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_87),
.C(n_82),
.Y(n_121)
);

AO22x1_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_45),
.B1(n_62),
.B2(n_48),
.Y(n_114)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_13),
.Y(n_117)
);

XNOR2x1_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_45),
.Y(n_132)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_119),
.B(n_82),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_80),
.A2(n_62),
.B1(n_20),
.B2(n_32),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_112),
.Y(n_155)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_115),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_125),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_136),
.B1(n_141),
.B2(n_144),
.Y(n_152)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_131),
.Y(n_147)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_113),
.Y(n_148)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_99),
.A2(n_84),
.B1(n_92),
.B2(n_74),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_106),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_137),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_88),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_143),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_98),
.A2(n_74),
.B1(n_88),
.B2(n_85),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_105),
.A2(n_88),
.B1(n_95),
.B2(n_20),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_120),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_109),
.C(n_117),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_146),
.B(n_150),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_159),
.Y(n_190)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_164),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_125),
.A2(n_103),
.B1(n_116),
.B2(n_105),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_168),
.C(n_142),
.Y(n_179)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_156),
.B(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_165),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_104),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_96),
.B(n_118),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_138),
.B(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_171),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_111),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_170),
.Y(n_194)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

NOR4xp25_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_111),
.C(n_30),
.D(n_22),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_172),
.B(n_1),
.Y(n_212)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_175),
.Y(n_197)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_169),
.A2(n_131),
.B1(n_126),
.B2(n_135),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_180),
.B1(n_181),
.B2(n_187),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_159),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_152),
.A2(n_134),
.B1(n_126),
.B2(n_128),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_186),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_143),
.C(n_130),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_179),
.C(n_190),
.Y(n_205)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_152),
.A2(n_108),
.B1(n_127),
.B2(n_20),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_163),
.B1(n_166),
.B2(n_162),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_28),
.B1(n_68),
.B2(n_3),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_0),
.B(n_1),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_189),
.B(n_0),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_22),
.Y(n_192)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_32),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_193),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_205),
.Y(n_217)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_149),
.C(n_168),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_198),
.B(n_203),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_199),
.A2(n_201),
.B1(n_208),
.B2(n_189),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_194),
.A2(n_148),
.B1(n_32),
.B2(n_28),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_200),
.A2(n_209),
.B1(n_214),
.B2(n_187),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_177),
.A2(n_28),
.B1(n_30),
.B2(n_3),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_192),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_172),
.B(n_10),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_204),
.B(n_212),
.Y(n_227)
);

OA21x2_ASAP7_75t_SL g207 ( 
.A1(n_191),
.A2(n_30),
.B(n_28),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_208),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_194),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_176),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_210),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_15),
.C(n_5),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_188),
.C(n_193),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_183),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_221),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_176),
.Y(n_218)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_184),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_211),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_202),
.A2(n_185),
.B1(n_183),
.B2(n_182),
.Y(n_220)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_224),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_196),
.Y(n_224)
);

INVx11_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_230),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_229),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_186),
.C(n_175),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_206),
.C(n_195),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g229 ( 
.A1(n_197),
.A2(n_174),
.B(n_178),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_202),
.A2(n_181),
.B1(n_180),
.B2(n_9),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_236),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_206),
.B1(n_209),
.B2(n_211),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_236),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_242),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_197),
.Y(n_239)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_239),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_212),
.C(n_213),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_222),
.C(n_227),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_219),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_250),
.C(n_240),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_228),
.C(n_216),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_232),
.C(n_12),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_226),
.Y(n_247)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_247),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_237),
.A2(n_225),
.B(n_227),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_248),
.A2(n_8),
.B(n_12),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_231),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_7),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_235),
.B1(n_241),
.B2(n_233),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_254),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_237),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_255),
.B(n_245),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_257),
.C(n_250),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_244),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_259),
.B(n_262),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_243),
.C(n_249),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_263),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_262),
.A2(n_253),
.B1(n_245),
.B2(n_13),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_265),
.Y(n_268)
);

A2O1A1O1Ixp25_ASAP7_75t_L g267 ( 
.A1(n_260),
.A2(n_8),
.B(n_12),
.C(n_13),
.D(n_14),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_14),
.C(n_15),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_264),
.C(n_266),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_268),
.C(n_14),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_15),
.Y(n_272)
);


endmodule