module real_aes_4470_n_249 (n_17, n_28, n_226, n_76, n_202, n_926, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_925, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_926;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_925;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_905;
wire n_503;
wire n_673;
wire n_386;
wire n_635;
wire n_518;
wire n_254;
wire n_792;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_909;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_898;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_526;
wire n_637;
wire n_653;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_922;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_259;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_0), .A2(n_45), .B1(n_687), .B2(n_690), .Y(n_695) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_1), .Y(n_645) );
AND2x4_ASAP7_75t_L g660 ( .A(n_1), .B(n_661), .Y(n_660) );
AND2x4_ASAP7_75t_L g670 ( .A(n_1), .B(n_243), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_2), .A2(n_98), .B1(n_304), .B2(n_305), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_3), .A2(n_135), .B1(n_294), .B2(n_416), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_4), .A2(n_55), .B1(n_294), .B2(n_301), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_5), .A2(n_162), .B1(n_261), .B2(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_6), .B(n_467), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_7), .A2(n_84), .B1(n_466), .B2(n_467), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_8), .A2(n_187), .B1(n_459), .B2(n_622), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_9), .A2(n_231), .B1(n_372), .B2(n_373), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_10), .A2(n_200), .B1(n_312), .B2(n_428), .Y(n_427) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_11), .A2(n_540), .B(n_541), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_12), .A2(n_214), .B1(n_369), .B2(n_370), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_13), .A2(n_78), .B1(n_680), .B2(n_694), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_14), .A2(n_27), .B1(n_301), .B2(n_532), .Y(n_531) );
AO22x1_ASAP7_75t_L g403 ( .A1(n_15), .A2(n_143), .B1(n_404), .B2(n_405), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_16), .A2(n_114), .B1(n_435), .B2(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g667 ( .A(n_17), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_18), .A2(n_51), .B1(n_334), .B2(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_19), .A2(n_155), .B1(n_318), .B2(n_321), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_20), .A2(n_219), .B1(n_545), .B2(n_546), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_21), .A2(n_178), .B1(n_415), .B2(n_416), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_22), .A2(n_109), .B1(n_321), .B2(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_23), .A2(n_145), .B1(n_428), .B2(n_527), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_24), .A2(n_190), .B1(n_418), .B2(n_456), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_25), .A2(n_76), .B1(n_673), .B2(n_703), .Y(n_753) );
INVx1_ASAP7_75t_SL g736 ( .A(n_26), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_26), .A2(n_899), .B1(n_901), .B2(n_920), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_28), .A2(n_97), .B1(n_363), .B2(n_364), .Y(n_602) );
INVx1_ASAP7_75t_L g907 ( .A(n_29), .Y(n_907) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_30), .A2(n_364), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g280 ( .A(n_31), .Y(n_280) );
INVxp67_ASAP7_75t_L g329 ( .A(n_31), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_31), .B(n_189), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_32), .A2(n_86), .B1(n_657), .B2(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_33), .A2(n_195), .B1(n_318), .B2(n_431), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_34), .A2(n_117), .B1(n_416), .B2(n_532), .Y(n_914) );
CKINVDCx5p33_ASAP7_75t_R g566 ( .A(n_35), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_36), .A2(n_90), .B1(n_589), .B2(n_590), .Y(n_588) );
AOI21xp33_ASAP7_75t_SL g511 ( .A1(n_37), .A2(n_512), .B(n_513), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_38), .A2(n_140), .B1(n_415), .B2(n_481), .Y(n_480) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_39), .A2(n_66), .B1(n_363), .B2(n_364), .C(n_365), .Y(n_362) );
AO22x1_ASAP7_75t_L g398 ( .A1(n_40), .A2(n_136), .B1(n_304), .B2(n_305), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_41), .B(n_337), .Y(n_336) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_42), .A2(n_102), .B1(n_261), .B2(n_283), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_43), .B(n_265), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_44), .A2(n_242), .B1(n_519), .B2(n_520), .Y(n_626) );
OAI21x1_ASAP7_75t_L g354 ( .A1(n_45), .A2(n_355), .B(n_378), .Y(n_354) );
NAND4xp25_ASAP7_75t_L g378 ( .A(n_45), .B(n_356), .C(n_361), .D(n_374), .Y(n_378) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_46), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_47), .A2(n_248), .B1(n_669), .B2(n_704), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_48), .A2(n_71), .B1(n_622), .B2(n_623), .C(n_624), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g306 ( .A1(n_49), .A2(n_170), .B1(n_307), .B2(n_312), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_50), .A2(n_175), .B1(n_312), .B2(n_358), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_52), .A2(n_83), .B1(n_372), .B2(n_373), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_53), .A2(n_225), .B1(n_492), .B2(n_545), .Y(n_627) );
INVxp67_ASAP7_75t_R g671 ( .A(n_54), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_56), .A2(n_246), .B1(n_420), .B2(n_564), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_57), .A2(n_157), .B1(n_534), .B2(n_916), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_58), .A2(n_105), .B1(n_545), .B2(n_546), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_59), .B(n_363), .Y(n_387) );
INVx2_ASAP7_75t_L g643 ( .A(n_60), .Y(n_643) );
AOI21xp33_ASAP7_75t_L g340 ( .A1(n_61), .A2(n_341), .B(n_343), .Y(n_340) );
XNOR2x1_ASAP7_75t_L g469 ( .A(n_62), .B(n_470), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_63), .A2(n_197), .B1(n_519), .B2(n_520), .Y(n_518) );
INVx1_ASAP7_75t_L g659 ( .A(n_64), .Y(n_659) );
AND2x4_ASAP7_75t_L g664 ( .A(n_64), .B(n_643), .Y(n_664) );
INVx1_ASAP7_75t_SL g681 ( .A(n_64), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_65), .A2(n_194), .B1(n_404), .B2(n_405), .Y(n_610) );
XNOR2x1_ASAP7_75t_L g536 ( .A(n_67), .B(n_537), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_68), .A2(n_69), .B1(n_428), .B2(n_454), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g904 ( .A1(n_70), .A2(n_905), .B(n_906), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_72), .A2(n_180), .B1(n_680), .B2(n_694), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_73), .A2(n_152), .B1(n_294), .B2(n_376), .Y(n_375) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_74), .Y(n_265) );
AOI22xp33_ASAP7_75t_SL g604 ( .A1(n_75), .A2(n_148), .B1(n_369), .B2(n_370), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_77), .A2(n_176), .B1(n_372), .B2(n_373), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_79), .A2(n_171), .B1(n_369), .B2(n_370), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_80), .A2(n_234), .B1(n_261), .B2(n_360), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_81), .A2(n_205), .B1(n_376), .B2(n_415), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_82), .A2(n_217), .B1(n_283), .B2(n_425), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_85), .A2(n_128), .B1(n_473), .B2(n_474), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_87), .A2(n_119), .B1(n_495), .B2(n_497), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g665 ( .A(n_88), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_89), .A2(n_159), .B1(n_657), .B2(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g266 ( .A(n_91), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_91), .B(n_188), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_92), .A2(n_230), .B1(n_442), .B2(n_893), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_93), .A2(n_160), .B1(n_451), .B2(n_478), .Y(n_549) );
INVx1_ASAP7_75t_L g366 ( .A(n_94), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_95), .A2(n_99), .B1(n_418), .B2(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g344 ( .A(n_96), .Y(n_344) );
INVx1_ASAP7_75t_L g682 ( .A(n_100), .Y(n_682) );
INVx1_ASAP7_75t_L g392 ( .A(n_101), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_103), .A2(n_161), .B1(n_703), .B2(n_704), .Y(n_702) );
INVx1_ASAP7_75t_L g886 ( .A(n_104), .Y(n_886) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_106), .A2(n_172), .B1(n_428), .B2(n_454), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_107), .A2(n_241), .B1(n_261), .B2(n_304), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_108), .B(n_489), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_110), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g330 ( .A1(n_111), .A2(n_196), .B1(n_331), .B2(n_334), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_112), .A2(n_222), .B1(n_478), .B2(n_534), .Y(n_875) );
INVx1_ASAP7_75t_L g440 ( .A(n_113), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_115), .A2(n_123), .B1(n_575), .B2(n_576), .Y(n_574) );
XNOR2x1_ASAP7_75t_L g411 ( .A(n_116), .B(n_412), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_118), .A2(n_122), .B1(n_526), .B2(n_527), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_120), .A2(n_164), .B1(n_669), .B2(n_673), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_121), .A2(n_240), .B1(n_418), .B2(n_481), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_124), .A2(n_133), .B1(n_526), .B2(n_527), .Y(n_525) );
AO22x1_ASAP7_75t_L g399 ( .A1(n_125), .A2(n_237), .B1(n_400), .B2(n_401), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_126), .A2(n_174), .B1(n_454), .B2(n_526), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_127), .A2(n_146), .B1(n_358), .B2(n_562), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_129), .A2(n_198), .B1(n_397), .B2(n_401), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_130), .A2(n_215), .B1(n_305), .B2(n_400), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_131), .A2(n_207), .B1(n_415), .B2(n_416), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_132), .A2(n_211), .B1(n_474), .B2(n_632), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_134), .A2(n_218), .B1(n_418), .B2(n_481), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_137), .A2(n_144), .B1(n_522), .B2(n_523), .Y(n_521) );
INVx1_ASAP7_75t_L g468 ( .A(n_138), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_139), .A2(n_201), .B1(n_304), .B2(n_305), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_141), .A2(n_244), .B1(n_585), .B2(n_587), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_142), .A2(n_156), .B1(n_450), .B2(n_451), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_147), .Y(n_569) );
INVx1_ASAP7_75t_L g685 ( .A(n_149), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_150), .A2(n_226), .B1(n_687), .B2(n_690), .Y(n_699) );
INVx1_ASAP7_75t_L g683 ( .A(n_151), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_153), .B(n_508), .Y(n_507) );
CKINVDCx14_ASAP7_75t_R g598 ( .A(n_154), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_158), .A2(n_224), .B1(n_476), .B2(n_478), .Y(n_475) );
XNOR2x2_ASAP7_75t_L g384 ( .A(n_161), .B(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_163), .B(n_442), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_165), .A2(n_221), .B1(n_418), .B2(n_420), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g434 ( .A1(n_166), .A2(n_202), .B1(n_435), .B2(n_437), .C(n_439), .Y(n_434) );
INVx1_ASAP7_75t_L g486 ( .A(n_167), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_168), .B(n_467), .Y(n_543) );
OA22x2_ASAP7_75t_L g270 ( .A1(n_169), .A2(n_189), .B1(n_265), .B2(n_269), .Y(n_270) );
INVx1_ASAP7_75t_L g290 ( .A(n_169), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_173), .A2(n_227), .B1(n_420), .B2(n_564), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_177), .A2(n_191), .B1(n_431), .B2(n_459), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_179), .A2(n_238), .B1(n_428), .B2(n_454), .Y(n_479) );
INVx1_ASAP7_75t_L g514 ( .A(n_181), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_182), .A2(n_199), .B1(n_416), .B2(n_532), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_183), .A2(n_210), .B1(n_478), .B2(n_534), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_184), .A2(n_229), .B1(n_459), .B2(n_495), .Y(n_547) );
CKINVDCx6p67_ASAP7_75t_R g662 ( .A(n_185), .Y(n_662) );
INVx1_ASAP7_75t_L g887 ( .A(n_186), .Y(n_887) );
INVx1_ASAP7_75t_L g282 ( .A(n_188), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_188), .B(n_288), .Y(n_353) );
OAI21xp33_ASAP7_75t_L g291 ( .A1(n_189), .A2(n_206), .B(n_292), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g618 ( .A(n_192), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_193), .A2(n_247), .B1(n_657), .B2(n_706), .Y(n_725) );
INVx1_ASAP7_75t_L g504 ( .A(n_203), .Y(n_504) );
INVx1_ASAP7_75t_L g881 ( .A(n_204), .Y(n_881) );
INVx1_ASAP7_75t_L g268 ( .A(n_206), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_206), .B(n_235), .Y(n_351) );
INVx1_ASAP7_75t_L g883 ( .A(n_208), .Y(n_883) );
CKINVDCx16_ASAP7_75t_R g542 ( .A(n_209), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_212), .A2(n_223), .B1(n_331), .B2(n_334), .Y(n_433) );
INVx1_ASAP7_75t_L g737 ( .A(n_213), .Y(n_737) );
INVx1_ASAP7_75t_L g890 ( .A(n_216), .Y(n_890) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_220), .A2(n_484), .B(n_485), .Y(n_483) );
INVx1_ASAP7_75t_L g257 ( .A(n_226), .Y(n_257) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_228), .A2(n_236), .B1(n_418), .B2(n_456), .Y(n_455) );
XOR2xp5_ASAP7_75t_L g901 ( .A(n_232), .B(n_902), .Y(n_901) );
CKINVDCx20_ASAP7_75t_R g591 ( .A(n_233), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_235), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_239), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g661 ( .A(n_243), .Y(n_661) );
HB1xp67_ASAP7_75t_L g922 ( .A(n_243), .Y(n_922) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_245), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_638), .B(n_646), .Y(n_249) );
XNOR2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_557), .Y(n_250) );
XNOR2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_407), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_380), .B1(n_381), .B2(n_406), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g406 ( .A(n_254), .Y(n_406) );
AO22x2_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B1(n_354), .B2(n_379), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
XNOR2x1_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NOR2x1_ASAP7_75t_L g258 ( .A(n_259), .B(n_316), .Y(n_258) );
NAND4xp25_ASAP7_75t_L g259 ( .A(n_260), .B(n_293), .C(n_303), .D(n_306), .Y(n_259) );
AND2x4_ASAP7_75t_L g261 ( .A(n_262), .B(n_271), .Y(n_261) );
AND2x4_ASAP7_75t_L g304 ( .A(n_262), .B(n_299), .Y(n_304) );
AND2x2_ASAP7_75t_L g333 ( .A(n_262), .B(n_310), .Y(n_333) );
AND2x2_ASAP7_75t_L g339 ( .A(n_262), .B(n_314), .Y(n_339) );
AND2x2_ASAP7_75t_L g363 ( .A(n_262), .B(n_314), .Y(n_363) );
AND2x4_ASAP7_75t_L g369 ( .A(n_262), .B(n_310), .Y(n_369) );
AND2x2_ASAP7_75t_L g419 ( .A(n_262), .B(n_299), .Y(n_419) );
AND2x4_ASAP7_75t_L g426 ( .A(n_262), .B(n_402), .Y(n_426) );
AND2x2_ASAP7_75t_L g477 ( .A(n_262), .B(n_299), .Y(n_477) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_270), .Y(n_262) );
INVx1_ASAP7_75t_L g297 ( .A(n_263), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
NAND2xp33_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g269 ( .A(n_265), .Y(n_269) );
INVx3_ASAP7_75t_L g275 ( .A(n_265), .Y(n_275) );
NAND2xp33_ASAP7_75t_L g281 ( .A(n_265), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g292 ( .A(n_265), .Y(n_292) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_265), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_266), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g328 ( .A1(n_268), .A2(n_292), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g298 ( .A(n_270), .Y(n_298) );
AND2x2_ASAP7_75t_L g320 ( .A(n_270), .B(n_297), .Y(n_320) );
AND2x2_ASAP7_75t_L g327 ( .A(n_270), .B(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g285 ( .A(n_271), .B(n_286), .Y(n_285) );
AND2x4_ASAP7_75t_L g302 ( .A(n_271), .B(n_296), .Y(n_302) );
AND2x4_ASAP7_75t_L g397 ( .A(n_271), .B(n_286), .Y(n_397) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g402 ( .A(n_272), .Y(n_402) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_277), .Y(n_272) );
AND2x4_ASAP7_75t_L g299 ( .A(n_273), .B(n_300), .Y(n_299) );
AND2x4_ASAP7_75t_L g310 ( .A(n_273), .B(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g315 ( .A(n_273), .Y(n_315) );
AND2x2_ASAP7_75t_L g323 ( .A(n_273), .B(n_324), .Y(n_323) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_275), .B(n_280), .Y(n_279) );
INVxp67_ASAP7_75t_L g288 ( .A(n_275), .Y(n_288) );
NAND3xp33_ASAP7_75t_L g352 ( .A(n_276), .B(n_287), .C(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g300 ( .A(n_277), .Y(n_300) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g311 ( .A(n_278), .Y(n_311) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_283), .Y(n_576) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx3_ASAP7_75t_L g360 ( .A(n_284), .Y(n_360) );
INVx5_ASAP7_75t_L g451 ( .A(n_284), .Y(n_451) );
INVx2_ASAP7_75t_L g474 ( .A(n_284), .Y(n_474) );
INVx6_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx12f_ASAP7_75t_L g534 ( .A(n_285), .Y(n_534) );
AND2x4_ASAP7_75t_L g305 ( .A(n_286), .B(n_299), .Y(n_305) );
AND2x4_ASAP7_75t_L g335 ( .A(n_286), .B(n_314), .Y(n_335) );
AND2x4_ASAP7_75t_L g373 ( .A(n_286), .B(n_314), .Y(n_373) );
AND2x4_ASAP7_75t_L g422 ( .A(n_286), .B(n_299), .Y(n_422) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_291), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_294), .Y(n_571) );
BUFx12f_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_295), .Y(n_415) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_295), .Y(n_532) );
AND2x4_ASAP7_75t_L g295 ( .A(n_296), .B(n_299), .Y(n_295) );
AND2x4_ASAP7_75t_L g309 ( .A(n_296), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g313 ( .A(n_296), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g400 ( .A(n_296), .B(n_299), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_296), .B(n_402), .Y(n_401) );
AND2x4_ASAP7_75t_L g404 ( .A(n_296), .B(n_310), .Y(n_404) );
AND2x4_ASAP7_75t_L g405 ( .A(n_296), .B(n_314), .Y(n_405) );
AND2x4_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_302), .Y(n_376) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_302), .Y(n_416) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_302), .Y(n_473) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g358 ( .A(n_308), .Y(n_358) );
INVx3_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx12f_ASAP7_75t_L g428 ( .A(n_309), .Y(n_428) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_309), .Y(n_526) );
AND2x4_ASAP7_75t_L g319 ( .A(n_310), .B(n_320), .Y(n_319) );
AND2x4_ASAP7_75t_L g372 ( .A(n_310), .B(n_320), .Y(n_372) );
AND2x4_ASAP7_75t_L g314 ( .A(n_311), .B(n_315), .Y(n_314) );
BUFx2_ASAP7_75t_L g562 ( .A(n_312), .Y(n_562) );
BUFx3_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_313), .Y(n_454) );
BUFx5_ASAP7_75t_L g527 ( .A(n_313), .Y(n_527) );
AND2x4_ASAP7_75t_L g342 ( .A(n_314), .B(n_320), .Y(n_342) );
AND2x2_ASAP7_75t_L g364 ( .A(n_314), .B(n_320), .Y(n_364) );
NAND4xp25_ASAP7_75t_L g316 ( .A(n_317), .B(n_330), .C(n_336), .D(n_340), .Y(n_316) );
INVx2_ASAP7_75t_L g586 ( .A(n_318), .Y(n_586) );
BUFx3_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx3_ASAP7_75t_L g461 ( .A(n_319), .Y(n_461) );
INVx1_ASAP7_75t_L g496 ( .A(n_319), .Y(n_496) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_319), .Y(n_622) );
BUFx4f_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx5_ASAP7_75t_L g432 ( .A(n_322), .Y(n_432) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_327), .Y(n_322) );
AND2x4_ASAP7_75t_L g370 ( .A(n_323), .B(n_327), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g348 ( .A(n_325), .Y(n_348) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g497 ( .A(n_332), .Y(n_497) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_333), .Y(n_459) );
BUFx3_ASAP7_75t_L g519 ( .A(n_333), .Y(n_519) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx3_ASAP7_75t_L g493 ( .A(n_335), .Y(n_493) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_335), .Y(n_523) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g484 ( .A(n_338), .Y(n_484) );
INVx2_ASAP7_75t_L g623 ( .A(n_338), .Y(n_623) );
INVx3_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx3_ASAP7_75t_L g466 ( .A(n_339), .Y(n_466) );
INVx2_ASAP7_75t_L g510 ( .A(n_339), .Y(n_510) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g436 ( .A(n_342), .Y(n_436) );
INVx2_ASAP7_75t_L g464 ( .A(n_342), .Y(n_464) );
BUFx3_ASAP7_75t_L g545 ( .A(n_342), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_345), .B(n_366), .Y(n_365) );
INVx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx4_ASAP7_75t_L g393 ( .A(n_346), .Y(n_393) );
INVx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_347), .Y(n_443) );
AO21x2_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_349), .B(n_352), .Y(n_347) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_349), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
INVx2_ASAP7_75t_L g379 ( .A(n_354), .Y(n_379) );
AND3x1_ASAP7_75t_L g355 ( .A(n_356), .B(n_361), .C(n_374), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_367), .Y(n_361) );
INVx2_ASAP7_75t_L g438 ( .A(n_363), .Y(n_438) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_371), .Y(n_367) );
INVx4_ASAP7_75t_L g487 ( .A(n_370), .Y(n_487) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx2_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_394), .Y(n_385) );
AND4x1_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .C(n_389), .D(n_390), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx4_ASAP7_75t_L g467 ( .A(n_393), .Y(n_467) );
INVx1_ASAP7_75t_L g582 ( .A(n_393), .Y(n_582) );
NOR4xp25_ASAP7_75t_L g394 ( .A(n_395), .B(n_398), .C(n_399), .D(n_403), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_499), .B1(n_500), .B2(n_556), .Y(n_407) );
INVx2_ASAP7_75t_L g556 ( .A(n_408), .Y(n_556) );
OA22x2_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_444), .B1(n_445), .B2(n_498), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g498 ( .A(n_410), .Y(n_498) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NAND4xp75_ASAP7_75t_L g412 ( .A(n_413), .B(n_423), .C(n_429), .D(n_434), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_417), .Y(n_413) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx8_ASAP7_75t_L g564 ( .A(n_419), .Y(n_564) );
INVx4_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx4_ASAP7_75t_L g456 ( .A(n_421), .Y(n_456) );
INVx4_ASAP7_75t_L g481 ( .A(n_421), .Y(n_481) );
INVx2_ASAP7_75t_L g529 ( .A(n_421), .Y(n_529) );
INVx8_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_427), .Y(n_423) );
BUFx3_ASAP7_75t_L g575 ( .A(n_425), .Y(n_575) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx12f_ASAP7_75t_L g450 ( .A(n_426), .Y(n_450) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_426), .Y(n_478) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_426), .Y(n_632) );
BUFx3_ASAP7_75t_L g916 ( .A(n_426), .Y(n_916) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_433), .Y(n_429) );
INVx2_ASAP7_75t_L g908 ( .A(n_431), .Y(n_908) );
INVx4_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g520 ( .A(n_432), .Y(n_520) );
INVx2_ASAP7_75t_L g893 ( .A(n_432), .Y(n_893) );
INVx2_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_SL g522 ( .A(n_436), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g885 ( .A1(n_436), .A2(n_886), .B1(n_887), .B2(n_888), .Y(n_885) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
INVx2_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_443), .Y(n_490) );
INVx2_ASAP7_75t_L g516 ( .A(n_443), .Y(n_516) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
XNOR2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_469), .Y(n_445) );
XOR2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_468), .Y(n_446) );
NOR2x1_ASAP7_75t_L g447 ( .A(n_448), .B(n_457), .Y(n_447) );
NAND4xp25_ASAP7_75t_L g448 ( .A(n_449), .B(n_452), .C(n_453), .D(n_455), .Y(n_448) );
NAND4xp25_ASAP7_75t_L g457 ( .A(n_458), .B(n_460), .C(n_462), .D(n_465), .Y(n_457) );
BUFx3_ASAP7_75t_L g587 ( .A(n_459), .Y(n_587) );
INVx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g589 ( .A(n_464), .Y(n_589) );
BUFx3_ASAP7_75t_L g580 ( .A(n_466), .Y(n_580) );
OR2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_482), .Y(n_470) );
NAND4xp25_ASAP7_75t_L g471 ( .A(n_472), .B(n_475), .C(n_479), .D(n_480), .Y(n_471) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_473), .Y(n_568) );
BUFx4f_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND3xp33_ASAP7_75t_SL g482 ( .A(n_483), .B(n_491), .C(n_494), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B(n_488), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g541 ( .A1(n_487), .A2(n_542), .B(n_543), .Y(n_541) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_490), .B(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx3_ASAP7_75t_L g546 ( .A(n_493), .Y(n_546) );
INVx2_ASAP7_75t_L g590 ( .A(n_493), .Y(n_590) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g512 ( .A(n_496), .Y(n_512) );
INVx2_ASAP7_75t_L g884 ( .A(n_497), .Y(n_884) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_535), .B1(n_553), .B2(n_555), .Y(n_500) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g554 ( .A(n_503), .Y(n_554) );
XNOR2x1_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
NOR4xp75_ASAP7_75t_L g505 ( .A(n_506), .B(n_517), .C(n_524), .D(n_530), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_511), .Y(n_506) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g540 ( .A(n_509), .Y(n_540) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
INVx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_521), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_525), .B(n_528), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_531), .B(n_533), .Y(n_530) );
INVx1_ASAP7_75t_L g555 ( .A(n_535), .Y(n_555) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_548), .Y(n_537) );
NAND3xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_544), .C(n_547), .Y(n_538) );
INVx1_ASAP7_75t_L g888 ( .A(n_546), .Y(n_888) );
NAND4xp25_ASAP7_75t_SL g548 ( .A(n_549), .B(n_550), .C(n_551), .D(n_552), .Y(n_548) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_594), .B1(n_595), .B2(n_637), .Y(n_557) );
INVx2_ASAP7_75t_L g637 ( .A(n_558), .Y(n_637) );
AO211x2_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_572), .B(n_592), .C(n_593), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_565), .Y(n_559) );
AO22x2_ASAP7_75t_L g593 ( .A1(n_560), .A2(n_573), .B1(n_591), .B2(n_926), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_561), .B(n_563), .Y(n_560) );
AO22x1_ASAP7_75t_L g592 ( .A1(n_565), .A2(n_583), .B1(n_591), .B2(n_925), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_567), .B1(n_569), .B2(n_570), .Y(n_565) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NOR3xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_583), .C(n_591), .Y(n_572) );
NAND2x1_ASAP7_75t_L g573 ( .A(n_574), .B(n_577), .Y(n_573) );
OA21x2_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_579), .B(n_581), .Y(n_577) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_588), .Y(n_583) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
AO22x2_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_614), .B1(n_634), .B2(n_636), .Y(n_595) );
INVx2_ASAP7_75t_L g636 ( .A(n_596), .Y(n_636) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OAI21x1_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B(n_611), .Y(n_597) );
NAND3xp33_ASAP7_75t_SL g611 ( .A(n_598), .B(n_612), .C(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_606), .Y(n_600) );
INVx1_ASAP7_75t_L g613 ( .A(n_601), .Y(n_613) );
NAND4xp25_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .C(n_604), .D(n_605), .Y(n_601) );
INVxp67_ASAP7_75t_L g612 ( .A(n_606), .Y(n_612) );
NAND4xp25_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .C(n_609), .D(n_610), .Y(n_606) );
INVxp67_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVxp67_ASAP7_75t_SL g635 ( .A(n_617), .Y(n_635) );
XNOR2x1_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
OR2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_628), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_626), .C(n_627), .Y(n_620) );
INVx4_ASAP7_75t_L g882 ( .A(n_622), .Y(n_882) );
INVx2_ASAP7_75t_L g891 ( .A(n_623), .Y(n_891) );
NAND4xp25_ASAP7_75t_SL g628 ( .A(n_629), .B(n_630), .C(n_631), .D(n_633), .Y(n_628) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
BUFx4_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
NAND3xp33_ASAP7_75t_L g640 ( .A(n_641), .B(n_644), .C(n_645), .Y(n_640) );
AND2x2_ASAP7_75t_L g895 ( .A(n_641), .B(n_896), .Y(n_895) );
AND2x2_ASAP7_75t_L g900 ( .A(n_641), .B(n_897), .Y(n_900) );
AOI21xp5_ASAP7_75t_L g923 ( .A1(n_641), .A2(n_645), .B(n_681), .Y(n_923) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AO21x1_ASAP7_75t_L g921 ( .A1(n_642), .A2(n_922), .B(n_923), .Y(n_921) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g658 ( .A(n_643), .B(n_659), .Y(n_658) );
AND3x4_ASAP7_75t_L g680 ( .A(n_643), .B(n_660), .C(n_681), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g896 ( .A(n_644), .B(n_897), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_645), .Y(n_897) );
OAI221xp5_ASAP7_75t_SL g646 ( .A1(n_647), .A2(n_867), .B1(n_870), .B2(n_894), .C(n_898), .Y(n_646) );
AND5x1_ASAP7_75t_L g647 ( .A(n_648), .B(n_811), .C(n_828), .D(n_837), .E(n_857), .Y(n_647) );
AOI222xp33_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_734), .B1(n_748), .B2(n_757), .C1(n_790), .C2(n_810), .Y(n_648) );
OAI221xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_728), .B1(n_734), .B2(n_739), .C(n_744), .Y(n_649) );
NOR3xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_707), .C(n_720), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_674), .Y(n_651) );
AND2x2_ASAP7_75t_L g862 ( .A(n_652), .B(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI221xp5_ASAP7_75t_L g707 ( .A1(n_653), .A2(n_708), .B1(n_713), .B2(n_717), .C(n_719), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_653), .B(n_785), .Y(n_784) );
BUFx2_ASAP7_75t_L g807 ( .A(n_653), .Y(n_807) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx3_ASAP7_75t_L g715 ( .A(n_654), .Y(n_715) );
AND2x2_ASAP7_75t_L g731 ( .A(n_654), .B(n_729), .Y(n_731) );
OR2x2_ASAP7_75t_L g765 ( .A(n_654), .B(n_723), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_654), .B(n_677), .Y(n_767) );
AND2x2_ASAP7_75t_L g779 ( .A(n_654), .B(n_723), .Y(n_779) );
OR2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_666), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_662), .B1(n_663), .B2(n_665), .Y(n_655) );
OAI221xp5_ASAP7_75t_L g735 ( .A1(n_656), .A2(n_663), .B1(n_736), .B2(n_737), .C(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g869 ( .A(n_656), .Y(n_869) );
INVx3_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
AND2x4_ASAP7_75t_L g669 ( .A(n_658), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g690 ( .A(n_658), .B(n_670), .Y(n_690) );
AND2x2_ASAP7_75t_L g703 ( .A(n_658), .B(n_670), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_660), .B(n_664), .Y(n_663) );
AND2x4_ASAP7_75t_L g694 ( .A(n_660), .B(n_664), .Y(n_694) );
AND2x4_ASAP7_75t_L g706 ( .A(n_660), .B(n_664), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_663), .A2(n_679), .B1(n_682), .B2(n_683), .Y(n_678) );
AND2x4_ASAP7_75t_L g673 ( .A(n_664), .B(n_670), .Y(n_673) );
AND2x2_ASAP7_75t_L g687 ( .A(n_664), .B(n_670), .Y(n_687) );
AND2x2_ASAP7_75t_L g704 ( .A(n_664), .B(n_670), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B1(n_671), .B2(n_672), .Y(n_666) );
INVx3_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_674), .B(n_773), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_691), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_675), .B(n_710), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_675), .B(n_773), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_675), .B(n_752), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_675), .B(n_709), .Y(n_866) );
INVx3_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
CKINVDCx6p67_ASAP7_75t_R g716 ( .A(n_677), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_677), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g760 ( .A(n_677), .B(n_733), .Y(n_760) );
AND2x2_ASAP7_75t_L g770 ( .A(n_677), .B(n_715), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_677), .B(n_715), .Y(n_798) );
AND2x2_ASAP7_75t_L g817 ( .A(n_677), .B(n_783), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_677), .B(n_712), .Y(n_853) );
OR2x6_ASAP7_75t_SL g677 ( .A(n_678), .B(n_684), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_686), .B1(n_688), .B2(n_689), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g772 ( .A(n_691), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_691), .B(n_709), .Y(n_832) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_696), .Y(n_691) );
CKINVDCx6p67_ASAP7_75t_R g712 ( .A(n_692), .Y(n_712) );
INVx1_ASAP7_75t_L g743 ( .A(n_692), .Y(n_743) );
OR2x2_ASAP7_75t_L g747 ( .A(n_692), .B(n_697), .Y(n_747) );
OAI32xp33_ASAP7_75t_L g763 ( .A1(n_692), .A2(n_747), .A3(n_764), .B1(n_765), .B2(n_766), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_692), .B(n_697), .Y(n_781) );
AND2x2_ASAP7_75t_L g783 ( .A(n_692), .B(n_710), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_692), .B(n_711), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_692), .B(n_733), .Y(n_861) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_695), .Y(n_692) );
INVx2_ASAP7_75t_SL g756 ( .A(n_694), .Y(n_756) );
OR2x2_ASAP7_75t_L g764 ( .A(n_696), .B(n_710), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_696), .B(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g814 ( .A(n_696), .B(n_712), .Y(n_814) );
INVx1_ASAP7_75t_L g852 ( .A(n_696), .Y(n_852) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_700), .Y(n_696) );
CKINVDCx5p33_ASAP7_75t_R g711 ( .A(n_697), .Y(n_711) );
AND2x2_ASAP7_75t_L g803 ( .A(n_697), .B(n_701), .Y(n_803) );
AND2x4_ASAP7_75t_SL g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx1_ASAP7_75t_L g718 ( .A(n_700), .Y(n_718) );
AND2x2_ASAP7_75t_L g727 ( .A(n_700), .B(n_712), .Y(n_727) );
AND2x2_ASAP7_75t_L g733 ( .A(n_700), .B(n_711), .Y(n_733) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g710 ( .A(n_701), .B(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_705), .Y(n_701) );
OAI211xp5_ASAP7_75t_SL g815 ( .A1(n_708), .A2(n_766), .B(n_816), .C(n_818), .Y(n_815) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_SL g709 ( .A(n_710), .B(n_712), .Y(n_709) );
AND2x2_ASAP7_75t_L g775 ( .A(n_710), .B(n_776), .Y(n_775) );
OAI21xp33_ASAP7_75t_L g805 ( .A1(n_710), .A2(n_714), .B(n_727), .Y(n_805) );
AND2x2_ASAP7_75t_L g844 ( .A(n_710), .B(n_820), .Y(n_844) );
OAI222xp33_ASAP7_75t_L g720 ( .A1(n_711), .A2(n_721), .B1(n_726), .B2(n_728), .C1(n_730), .C2(n_732), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_711), .B(n_742), .Y(n_741) );
AOI22xp33_ASAP7_75t_SL g791 ( .A1(n_711), .A2(n_779), .B1(n_792), .B2(n_793), .Y(n_791) );
AND2x2_ASAP7_75t_L g776 ( .A(n_712), .B(n_716), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_712), .B(n_733), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_712), .B(n_803), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_712), .B(n_824), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_712), .B(n_760), .Y(n_839) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_714), .B(n_749), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
AND2x2_ASAP7_75t_L g722 ( .A(n_715), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g745 ( .A(n_715), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_715), .B(n_771), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_715), .B(n_819), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_715), .B(n_844), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_716), .B(n_722), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_716), .B(n_741), .Y(n_740) );
NOR2x1p5_ASAP7_75t_L g746 ( .A(n_716), .B(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_716), .B(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g795 ( .A(n_716), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_716), .B(n_814), .Y(n_813) );
AND2x2_ASAP7_75t_L g820 ( .A(n_716), .B(n_742), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_716), .B(n_731), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_716), .B(n_765), .Y(n_836) );
INVx1_ASAP7_75t_L g797 ( .A(n_717), .Y(n_797) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVxp67_ASAP7_75t_L g858 ( .A(n_721), .Y(n_858) );
INVx1_ASAP7_75t_L g804 ( .A(n_722), .Y(n_804) );
INVx2_ASAP7_75t_L g729 ( .A(n_723), .Y(n_729) );
AND2x2_ASAP7_75t_L g842 ( .A(n_723), .B(n_752), .Y(n_842) );
AND2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g782 ( .A1(n_727), .A2(n_783), .B1(n_784), .B2(n_786), .C(n_787), .Y(n_782) );
AOI211xp5_ASAP7_75t_L g799 ( .A1(n_727), .A2(n_800), .B(n_801), .C(n_808), .Y(n_799) );
OAI211xp5_ASAP7_75t_SL g757 ( .A1(n_728), .A2(n_758), .B(n_761), .C(n_782), .Y(n_757) );
INVx3_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OR2x2_ASAP7_75t_L g771 ( .A(n_729), .B(n_752), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_729), .B(n_751), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_729), .B(n_752), .Y(n_864) );
OAI221xp5_ASAP7_75t_L g845 ( .A1(n_730), .A2(n_846), .B1(n_848), .B2(n_850), .C(n_854), .Y(n_845) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
BUFx3_ASAP7_75t_L g810 ( .A(n_735), .Y(n_810) );
XNOR2x1_ASAP7_75t_L g872 ( .A(n_736), .B(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g759 ( .A(n_742), .B(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
INVx3_ASAP7_75t_L g762 ( .A(n_748), .Y(n_762) );
OAI311xp33_ASAP7_75t_L g801 ( .A1(n_748), .A2(n_802), .A3(n_804), .B1(n_805), .C1(n_806), .Y(n_801) );
INVx3_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx3_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_750), .B(n_809), .Y(n_808) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_751), .B(n_775), .Y(n_774) );
INVx3_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g785 ( .A(n_752), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_752), .B(n_779), .Y(n_789) );
AND2x2_ASAP7_75t_L g826 ( .A(n_752), .B(n_827), .Y(n_826) );
AND2x4_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
AOI211xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_763), .B(n_768), .C(n_777), .Y(n_761) );
INVx1_ASAP7_75t_L g827 ( .A(n_765), .Y(n_827) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
OAI221xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_771), .B1(n_772), .B2(n_773), .C(n_774), .Y(n_768) );
INVx1_ASAP7_75t_L g793 ( .A(n_771), .Y(n_793) );
OAI221xp5_ASAP7_75t_SL g790 ( .A1(n_773), .A2(n_791), .B1(n_794), .B2(n_796), .C(n_799), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_776), .B(n_803), .Y(n_856) );
AOI21xp33_ASAP7_75t_SL g777 ( .A1(n_778), .A2(n_780), .B(n_781), .Y(n_777) );
AOI211xp5_ASAP7_75t_SL g837 ( .A1(n_779), .A2(n_838), .B(n_840), .C(n_845), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_781), .B(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g859 ( .A(n_781), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_783), .B(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g809 ( .A(n_783), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g846 ( .A(n_783), .B(n_847), .Y(n_846) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
INVx1_ASAP7_75t_L g792 ( .A(n_788), .Y(n_792) );
AOI221xp5_ASAP7_75t_L g811 ( .A1(n_793), .A2(n_800), .B1(n_812), .B2(n_815), .C(n_821), .Y(n_811) );
CKINVDCx14_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
AND2x2_ASAP7_75t_L g819 ( .A(n_803), .B(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g824 ( .A(n_803), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_807), .B(n_817), .Y(n_816) );
AOI322xp5_ASAP7_75t_L g857 ( .A1(n_810), .A2(n_842), .A3(n_858), .B1(n_859), .B2(n_860), .C1(n_862), .C2(n_865), .Y(n_857) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_825), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_827), .B(n_849), .Y(n_848) );
OAI21xp33_ASAP7_75t_L g854 ( .A1(n_827), .A2(n_842), .B(n_855), .Y(n_854) );
AOI211xp5_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_831), .B(n_833), .C(n_834), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVxp67_ASAP7_75t_SL g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_841), .B(n_843), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
NOR2xp33_ASAP7_75t_L g851 ( .A(n_852), .B(n_853), .Y(n_851) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
CKINVDCx5p33_ASAP7_75t_R g867 ( .A(n_868), .Y(n_867) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx2_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
AND2x2_ASAP7_75t_L g873 ( .A(n_874), .B(n_879), .Y(n_873) );
AND4x1_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .C(n_877), .D(n_878), .Y(n_874) );
NOR3xp33_ASAP7_75t_L g879 ( .A(n_880), .B(n_885), .C(n_889), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_881), .A2(n_882), .B1(n_883), .B2(n_884), .Y(n_880) );
OAI21xp33_ASAP7_75t_L g889 ( .A1(n_890), .A2(n_891), .B(n_892), .Y(n_889) );
INVx1_ASAP7_75t_L g905 ( .A(n_891), .Y(n_905) );
CKINVDCx20_ASAP7_75t_R g894 ( .A(n_895), .Y(n_894) );
BUFx2_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
HB1xp67_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
NAND4xp75_ASAP7_75t_L g903 ( .A(n_904), .B(n_910), .C(n_913), .D(n_917), .Y(n_903) );
OAI21xp5_ASAP7_75t_L g906 ( .A1(n_907), .A2(n_908), .B(n_909), .Y(n_906) );
AND2x2_ASAP7_75t_L g910 ( .A(n_911), .B(n_912), .Y(n_910) );
AND2x2_ASAP7_75t_L g913 ( .A(n_914), .B(n_915), .Y(n_913) );
AND2x2_ASAP7_75t_L g917 ( .A(n_918), .B(n_919), .Y(n_917) );
BUFx2_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
endmodule