module fake_jpeg_12265_n_383 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_383);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_383;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_38),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_60),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_23),
.A2(n_7),
.B1(n_1),
.B2(n_2),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_19),
.B1(n_29),
.B2(n_28),
.Y(n_86)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_53),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_22),
.A2(n_7),
.B(n_1),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_34),
.C(n_32),
.Y(n_66)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_30),
.B(n_8),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx2_ASAP7_75t_R g62 ( 
.A(n_61),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_66),
.B(n_25),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_36),
.A2(n_20),
.B1(n_32),
.B2(n_34),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_70),
.A2(n_86),
.B1(n_28),
.B2(n_27),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_34),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_37),
.B(n_32),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_38),
.B(n_22),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_29),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_43),
.A2(n_16),
.B(n_17),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_66),
.C(n_62),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_50),
.A2(n_20),
.B1(n_25),
.B2(n_16),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_61),
.B1(n_40),
.B2(n_45),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_22),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_57),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g94 ( 
.A1(n_44),
.A2(n_29),
.B(n_28),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_42),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_63),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_97),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_101),
.B(n_103),
.Y(n_163)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_104),
.A2(n_122),
.B1(n_123),
.B2(n_131),
.Y(n_159)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_106),
.B(n_115),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_27),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_121),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_84),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_109),
.Y(n_157)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_110),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_111),
.A2(n_124),
.B1(n_125),
.B2(n_129),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_70),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_112),
.Y(n_146)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_114),
.Y(n_141)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_119),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_50),
.B1(n_45),
.B2(n_40),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_48),
.B1(n_54),
.B2(n_49),
.Y(n_136)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_120),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_67),
.B(n_41),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_42),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_42),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_65),
.B1(n_20),
.B2(n_55),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_61),
.C(n_18),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_51),
.B(n_77),
.Y(n_154)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_130),
.A2(n_85),
.B1(n_76),
.B2(n_80),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_62),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_47),
.B1(n_48),
.B2(n_54),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g183 ( 
.A1(n_135),
.A2(n_136),
.B1(n_143),
.B2(n_88),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_99),
.A2(n_128),
.B1(n_107),
.B2(n_126),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_137),
.A2(n_140),
.B1(n_142),
.B2(n_156),
.Y(n_176)
);

OAI32xp33_ASAP7_75t_L g139 ( 
.A1(n_99),
.A2(n_46),
.A3(n_79),
.B1(n_39),
.B2(n_83),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_80),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_103),
.A2(n_49),
.B1(n_47),
.B2(n_59),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_104),
.A2(n_68),
.B1(n_53),
.B2(n_83),
.Y(n_142)
);

NAND2x1p5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_117),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_64),
.B1(n_59),
.B2(n_81),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_147),
.A2(n_149),
.B1(n_165),
.B2(n_58),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_68),
.B1(n_46),
.B2(n_35),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_151),
.B(n_18),
.Y(n_193)
);

NOR3xp33_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_8),
.C(n_2),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_102),
.C(n_130),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_116),
.A2(n_65),
.B(n_77),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_155),
.A2(n_113),
.B(n_129),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_110),
.A2(n_88),
.B1(n_20),
.B2(n_58),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_166),
.A2(n_200),
.B1(n_145),
.B2(n_161),
.Y(n_216)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_192),
.C(n_155),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_114),
.Y(n_169)
);

INVxp33_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_163),
.B(n_98),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_171),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_105),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_172),
.A2(n_175),
.B(n_189),
.Y(n_202)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_173),
.Y(n_226)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_174),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_96),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_19),
.B(n_31),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_178),
.A2(n_194),
.B(n_198),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_125),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_181),
.Y(n_207)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_120),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_141),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_184),
.Y(n_214)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_183),
.Y(n_235)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_137),
.A2(n_100),
.B1(n_111),
.B2(n_124),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_185),
.A2(n_201),
.B1(n_4),
.B2(n_5),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_80),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_186),
.B(n_144),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_141),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_196),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_27),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_190),
.Y(n_220)
);

A2O1A1O1Ixp25_ASAP7_75t_L g189 ( 
.A1(n_164),
.A2(n_143),
.B(n_151),
.C(n_159),
.D(n_160),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_31),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_31),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_195),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_143),
.B(n_116),
.C(n_55),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_165),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_160),
.A2(n_18),
.B(n_17),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_17),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_132),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_0),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_0),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_164),
.A2(n_0),
.B(n_1),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_198),
.A2(n_148),
.B(n_158),
.Y(n_222)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_133),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_148),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_142),
.A2(n_8),
.B1(n_2),
.B2(n_3),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_197),
.A2(n_140),
.B1(n_139),
.B2(n_154),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_204),
.A2(n_208),
.B1(n_209),
.B2(n_216),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_166),
.A2(n_135),
.B1(n_144),
.B2(n_136),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_172),
.B1(n_176),
.B2(n_191),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_211),
.C(n_215),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_149),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_212),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_141),
.C(n_158),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_194),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_182),
.A2(n_161),
.B1(n_145),
.B2(n_150),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_223),
.A2(n_224),
.B1(n_232),
.B2(n_9),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_176),
.A2(n_147),
.B1(n_145),
.B2(n_133),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_189),
.A2(n_161),
.B(n_2),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_233),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_186),
.B(n_3),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_234),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_190),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_171),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_179),
.B(n_4),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_236),
.A2(n_167),
.B1(n_173),
.B2(n_188),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_237),
.A2(n_240),
.B1(n_243),
.B2(n_245),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_235),
.A2(n_195),
.B1(n_168),
.B2(n_183),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_219),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_241),
.B(n_259),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_235),
.A2(n_183),
.B1(n_187),
.B2(n_185),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_244),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_183),
.B1(n_175),
.B2(n_196),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_193),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_246),
.B(n_250),
.Y(n_292)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_247),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_212),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_199),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_202),
.B(n_178),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_254),
.C(n_257),
.Y(n_278)
);

INVx3_ASAP7_75t_SL g252 ( 
.A(n_224),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_221),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_202),
.B(n_180),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_206),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_261),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_174),
.C(n_184),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_214),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_210),
.B(n_201),
.C(n_9),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_263),
.C(n_230),
.Y(n_284)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_6),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_262),
.B(n_232),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_6),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_265),
.A2(n_236),
.B1(n_229),
.B2(n_234),
.Y(n_269)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_227),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_269),
.A2(n_260),
.B1(n_247),
.B2(n_267),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_270),
.B(n_251),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_258),
.A2(n_225),
.B1(n_205),
.B2(n_207),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_271),
.A2(n_290),
.B(n_13),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_272),
.B(n_273),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_264),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_239),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_275),
.A2(n_287),
.B1(n_11),
.B2(n_12),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_240),
.A2(n_209),
.B1(n_245),
.B2(n_243),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_276),
.A2(n_281),
.B1(n_289),
.B2(n_293),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_255),
.A2(n_207),
.B1(n_217),
.B2(n_205),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_277),
.A2(n_279),
.B1(n_249),
.B2(n_257),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_258),
.A2(n_218),
.B1(n_204),
.B2(n_226),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_252),
.A2(n_208),
.B1(n_214),
.B2(n_219),
.Y(n_281)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_237),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_283),
.B(n_284),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_238),
.B(n_211),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_248),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_242),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_253),
.A2(n_228),
.B1(n_227),
.B2(n_231),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_253),
.A2(n_222),
.B(n_228),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_249),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_242),
.Y(n_295)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_295),
.Y(n_330)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_296),
.Y(n_318)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_312),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_238),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_298),
.B(n_302),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_299),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_304),
.C(n_305),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_254),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_303),
.B(n_313),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_270),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_269),
.A2(n_267),
.B1(n_266),
.B2(n_263),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_306),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_9),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_293),
.C(n_280),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_279),
.A2(n_271),
.B1(n_282),
.B2(n_290),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_311),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_289),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_276),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_274),
.A2(n_14),
.B1(n_11),
.B2(n_13),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_314),
.B(n_316),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_286),
.B(n_280),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_281),
.B(n_14),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_319),
.A2(n_300),
.B1(n_314),
.B2(n_291),
.Y(n_341)
);

INVx13_ASAP7_75t_L g321 ( 
.A(n_294),
.Y(n_321)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_321),
.Y(n_335)
);

FAx1_ASAP7_75t_SL g322 ( 
.A(n_295),
.B(n_284),
.CI(n_292),
.CON(n_322),
.SN(n_322)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_322),
.B(n_328),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_294),
.B(n_274),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_326),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_307),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_298),
.B(n_286),
.C(n_291),
.Y(n_328)
);

INVx13_ASAP7_75t_L g333 ( 
.A(n_296),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_333),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_334),
.B(n_336),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_332),
.B(n_303),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_320),
.Y(n_337)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_337),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_325),
.A2(n_300),
.B1(n_316),
.B2(n_313),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_338),
.B(n_324),
.Y(n_350)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_318),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_340),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_305),
.C(n_301),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_341),
.A2(n_329),
.B1(n_330),
.B2(n_326),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_328),
.B(n_302),
.C(n_310),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_346),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_317),
.B(n_309),
.C(n_304),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_323),
.A2(n_308),
.B1(n_315),
.B2(n_330),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_347),
.A2(n_319),
.B1(n_329),
.B2(n_327),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_336),
.B(n_317),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_348),
.B(n_342),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_350),
.B(n_356),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_352),
.A2(n_343),
.B1(n_344),
.B2(n_341),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_335),
.B(n_318),
.Y(n_355)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_355),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_345),
.B(n_324),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_347),
.B(n_322),
.Y(n_357)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_357),
.Y(n_363)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_358),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_360),
.B(n_361),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_322),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_362),
.B(n_365),
.Y(n_372)
);

MAJx2_ASAP7_75t_L g365 ( 
.A(n_353),
.B(n_346),
.C(n_340),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_326),
.C(n_334),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_SL g370 ( 
.A(n_366),
.B(n_358),
.Y(n_370)
);

AO21x1_ASAP7_75t_L g368 ( 
.A1(n_363),
.A2(n_344),
.B(n_351),
.Y(n_368)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_368),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_364),
.A2(n_353),
.B(n_354),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_369),
.A2(n_370),
.B(n_373),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_331),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_371),
.A2(n_367),
.B(n_366),
.Y(n_374)
);

A2O1A1O1Ixp25_ASAP7_75t_L g379 ( 
.A1(n_374),
.A2(n_365),
.B(n_333),
.C(n_360),
.D(n_352),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_372),
.B(n_362),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_376),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_379),
.B(n_377),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_380),
.B(n_378),
.C(n_375),
.Y(n_381)
);

MAJx2_ASAP7_75t_L g382 ( 
.A(n_381),
.B(n_333),
.C(n_321),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_382),
.B(n_331),
.Y(n_383)
);


endmodule