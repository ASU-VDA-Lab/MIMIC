module fake_netlist_6_328_n_1671 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1671);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1671;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_34),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_54),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_61),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_86),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_55),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_133),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_76),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_119),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_57),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_87),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_66),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_98),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_142),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_75),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_93),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_9),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_53),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_91),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_43),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_19),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_58),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_35),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_33),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_43),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_73),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_5),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_104),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_11),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_42),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_83),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_28),
.Y(n_189)
);

BUFx8_ASAP7_75t_SL g190 ( 
.A(n_30),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_41),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_44),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_136),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_7),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_85),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_143),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_112),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_11),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_90),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_59),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_81),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_101),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_41),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_71),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_130),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_15),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_147),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_70),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_25),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_31),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_118),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_128),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_134),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_109),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_97),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_114),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_107),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_117),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_25),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_47),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_69),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_126),
.Y(n_224)
);

BUFx2_ASAP7_75t_SL g225 ( 
.A(n_64),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_31),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_49),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_45),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_82),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_56),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_37),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_39),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_148),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_51),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_48),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_3),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_29),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_12),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_127),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_35),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_121),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_52),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_77),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_49),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_47),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_122),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_7),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_28),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_78),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_50),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_60),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_40),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_33),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_125),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_74),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_6),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_2),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_13),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_45),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_15),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_103),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_129),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_12),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_151),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_140),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_84),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_1),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_5),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_149),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_80),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_16),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_32),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_88),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_13),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_124),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_137),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_6),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_110),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_18),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_37),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_116),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_131),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_32),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_40),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_10),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_92),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_63),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_19),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_68),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_48),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_34),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_106),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_18),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_44),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_14),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_23),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_22),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_4),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_96),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_16),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_67),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_38),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_190),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_272),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_174),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_272),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_160),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_154),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_239),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_156),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_180),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_272),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_180),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_272),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_155),
.B(n_0),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_291),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_243),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_158),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_200),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_201),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_272),
.Y(n_321)
);

INVxp33_ASAP7_75t_SL g322 ( 
.A(n_174),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_159),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_161),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_184),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_187),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_187),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_199),
.B(n_0),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_199),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_184),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_162),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_189),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_208),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_164),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_207),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_208),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_165),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_246),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_200),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_170),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_280),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_280),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_189),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_232),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_166),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_168),
.B(n_1),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_167),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_232),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_173),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_256),
.B(n_2),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_256),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_169),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_273),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_258),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_171),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_291),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_172),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_176),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_258),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_188),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_267),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_267),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_200),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_178),
.Y(n_364)
);

NOR2xp67_ASAP7_75t_L g365 ( 
.A(n_211),
.B(n_3),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_193),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_179),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_271),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_271),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_197),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_198),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_284),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_155),
.B(n_4),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_304),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_311),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_308),
.B(n_168),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_330),
.B(n_253),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_304),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_310),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_306),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_318),
.B(n_183),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_323),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_324),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_306),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_331),
.B(n_183),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_312),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_316),
.B(n_185),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_312),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_334),
.Y(n_389)
);

BUFx8_ASAP7_75t_L g390 ( 
.A(n_325),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_313),
.B(n_216),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_337),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_325),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_319),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_316),
.B(n_181),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_340),
.Y(n_396)
);

OAI21x1_ASAP7_75t_L g397 ( 
.A1(n_319),
.A2(n_281),
.B(n_265),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_321),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_321),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_345),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_314),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_309),
.B(n_253),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_347),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_R g404 ( 
.A(n_358),
.B(n_203),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_319),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_343),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_322),
.B(n_153),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_363),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_352),
.B(n_265),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_363),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_343),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_355),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_344),
.Y(n_413)
);

BUFx8_ASAP7_75t_L g414 ( 
.A(n_350),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_344),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_357),
.B(n_281),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_R g417 ( 
.A(n_366),
.B(n_204),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_309),
.B(n_284),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_360),
.B(n_206),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_309),
.B(n_317),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_307),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_348),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_348),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_339),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_351),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_351),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_354),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_339),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_339),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_354),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_359),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_370),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_371),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_363),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_320),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_359),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_363),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_317),
.B(n_296),
.Y(n_438)
);

OA21x2_ASAP7_75t_L g439 ( 
.A1(n_346),
.A2(n_163),
.B(n_157),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_303),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_317),
.B(n_296),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_335),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_421),
.B(n_338),
.Y(n_443)
);

INVx5_ASAP7_75t_L g444 ( 
.A(n_437),
.Y(n_444)
);

AND2x6_ASAP7_75t_L g445 ( 
.A(n_418),
.B(n_157),
.Y(n_445)
);

AND2x6_ASAP7_75t_L g446 ( 
.A(n_418),
.B(n_163),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_437),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_437),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g449 ( 
.A1(n_439),
.A2(n_373),
.B1(n_315),
.B2(n_346),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_401),
.B(n_349),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_376),
.B(n_364),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_420),
.B(n_367),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_381),
.B(n_305),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_406),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_393),
.B(n_356),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_437),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_442),
.Y(n_457)
);

BUFx10_ASAP7_75t_L g458 ( 
.A(n_440),
.Y(n_458)
);

OAI22xp33_ASAP7_75t_L g459 ( 
.A1(n_391),
.A2(n_350),
.B1(n_305),
.B2(n_226),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_420),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_406),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_393),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_411),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_411),
.Y(n_465)
);

AO22x2_ASAP7_75t_L g466 ( 
.A1(n_387),
.A2(n_297),
.B1(n_298),
.B2(n_195),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_402),
.B(n_361),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_L g468 ( 
.A(n_385),
.B(n_200),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_396),
.A2(n_353),
.B1(n_365),
.B2(n_254),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_437),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_394),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_394),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_439),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_408),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_413),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_413),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_420),
.B(n_200),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_377),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_375),
.B(n_209),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_402),
.B(n_361),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_415),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_379),
.B(n_214),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_382),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_377),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_415),
.Y(n_485)
);

BUFx4f_ASAP7_75t_L g486 ( 
.A(n_439),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_422),
.Y(n_487)
);

OAI22xp33_ASAP7_75t_L g488 ( 
.A1(n_409),
.A2(n_191),
.B1(n_212),
.B2(n_238),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_439),
.A2(n_328),
.B1(n_365),
.B2(n_332),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_383),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_420),
.B(n_218),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_389),
.Y(n_492)
);

INVx5_ASAP7_75t_L g493 ( 
.A(n_394),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_392),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_394),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_422),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_410),
.Y(n_497)
);

NAND2xp33_ASAP7_75t_SL g498 ( 
.A(n_404),
.B(n_228),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_438),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_394),
.Y(n_500)
);

INVx5_ASAP7_75t_L g501 ( 
.A(n_394),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_416),
.B(n_220),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_438),
.A2(n_328),
.B1(n_332),
.B2(n_247),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_410),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_419),
.B(n_223),
.Y(n_505)
);

BUFx4f_ASAP7_75t_L g506 ( 
.A(n_441),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_423),
.Y(n_507)
);

OR2x6_ASAP7_75t_L g508 ( 
.A(n_395),
.B(n_225),
.Y(n_508)
);

OAI22xp33_ASAP7_75t_L g509 ( 
.A1(n_400),
.A2(n_283),
.B1(n_302),
.B2(n_300),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_390),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_403),
.B(n_362),
.Y(n_511)
);

NAND2x1_ASAP7_75t_L g512 ( 
.A(n_374),
.B(n_175),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_424),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_414),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_390),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_434),
.Y(n_516)
);

INVx5_ASAP7_75t_L g517 ( 
.A(n_424),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_412),
.B(n_362),
.Y(n_518)
);

AND2x2_ASAP7_75t_SL g519 ( 
.A(n_441),
.B(n_175),
.Y(n_519)
);

NAND2xp33_ASAP7_75t_L g520 ( 
.A(n_432),
.B(n_224),
.Y(n_520)
);

OR2x6_ASAP7_75t_L g521 ( 
.A(n_390),
.B(n_225),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_433),
.B(n_368),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_390),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_374),
.B(n_230),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_424),
.Y(n_525)
);

NAND2xp33_ASAP7_75t_L g526 ( 
.A(n_417),
.B(n_234),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_414),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_378),
.B(n_241),
.Y(n_528)
);

BUFx8_ASAP7_75t_SL g529 ( 
.A(n_407),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_414),
.A2(n_242),
.B1(n_250),
.B2(n_299),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_414),
.B(n_177),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_378),
.B(n_262),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_380),
.B(n_266),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_423),
.A2(n_261),
.B1(n_182),
.B2(n_195),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_435),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_380),
.B(n_368),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_425),
.B(n_269),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_384),
.B(n_270),
.Y(n_538)
);

INVx5_ASAP7_75t_L g539 ( 
.A(n_424),
.Y(n_539)
);

OAI22xp33_ASAP7_75t_L g540 ( 
.A1(n_425),
.A2(n_222),
.B1(n_295),
.B2(n_294),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_384),
.B(n_369),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_424),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_386),
.B(n_369),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_407),
.B(n_372),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_424),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_386),
.B(n_372),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g547 ( 
.A(n_426),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_426),
.B(n_326),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_434),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_428),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_388),
.B(n_275),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_427),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_388),
.B(n_278),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_427),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_430),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_428),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_428),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_398),
.B(n_186),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_430),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_431),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_431),
.B(n_177),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_436),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_398),
.B(n_192),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_436),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_399),
.B(n_282),
.Y(n_565)
);

BUFx10_ASAP7_75t_L g566 ( 
.A(n_399),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_428),
.B(n_289),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_405),
.B(n_194),
.Y(n_568)
);

INVx5_ASAP7_75t_L g569 ( 
.A(n_428),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_428),
.B(n_182),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_405),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_397),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_429),
.B(n_196),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_405),
.B(n_429),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_429),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_397),
.B(n_205),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_401),
.B(n_221),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_391),
.B(n_227),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_391),
.B(n_231),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_401),
.B(n_235),
.Y(n_580)
);

INVxp67_ASAP7_75t_SL g581 ( 
.A(n_401),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_437),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_401),
.B(n_196),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_437),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_554),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_453),
.B(n_236),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_506),
.B(n_202),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_489),
.B(n_202),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_460),
.Y(n_589)
);

O2A1O1Ixp5_ASAP7_75t_L g590 ( 
.A1(n_486),
.A2(n_215),
.B(n_301),
.C(n_292),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_499),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_544),
.B(n_237),
.Y(n_592)
);

A2O1A1Ixp33_ASAP7_75t_L g593 ( 
.A1(n_453),
.A2(n_449),
.B(n_486),
.C(n_534),
.Y(n_593)
);

O2A1O1Ixp33_ASAP7_75t_L g594 ( 
.A1(n_478),
.A2(n_215),
.B(n_301),
.C(n_292),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_485),
.B(n_210),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_485),
.B(n_213),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_547),
.B(n_213),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_506),
.B(n_217),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_519),
.B(n_217),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_547),
.B(n_219),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_516),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_548),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_454),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_511),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_549),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_581),
.B(n_219),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_581),
.B(n_229),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_467),
.B(n_233),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_519),
.B(n_233),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_461),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_575),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_474),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_451),
.B(n_240),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_451),
.B(n_249),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_447),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_484),
.B(n_449),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_473),
.B(n_249),
.Y(n_617)
);

INVxp67_ASAP7_75t_SL g618 ( 
.A(n_448),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_559),
.B(n_251),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_473),
.B(n_511),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_464),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_518),
.B(n_255),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_567),
.A2(n_286),
.B(n_287),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_465),
.Y(n_624)
);

AND2x2_ASAP7_75t_SL g625 ( 
.A(n_534),
.B(n_261),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_518),
.B(n_264),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_522),
.B(n_452),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_475),
.B(n_264),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_522),
.B(n_276),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_564),
.B(n_276),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_476),
.B(n_286),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_481),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_487),
.B(n_287),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_467),
.B(n_480),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_497),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_496),
.B(n_507),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_552),
.B(n_555),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_560),
.B(n_277),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_508),
.A2(n_279),
.B1(n_245),
.B2(n_248),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_562),
.B(n_285),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_463),
.Y(n_641)
);

INVx8_ASAP7_75t_L g642 ( 
.A(n_521),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_480),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_455),
.B(n_342),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_504),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_535),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_450),
.B(n_342),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_570),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_571),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_571),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_505),
.B(n_274),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_491),
.B(n_288),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_566),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_448),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_448),
.Y(n_655)
);

AND2x6_ASAP7_75t_SL g656 ( 
.A(n_508),
.B(n_521),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_466),
.Y(n_657)
);

OR2x6_ASAP7_75t_L g658 ( 
.A(n_521),
.B(n_510),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_566),
.Y(n_659)
);

NAND3xp33_ASAP7_75t_L g660 ( 
.A(n_450),
.B(n_268),
.C(n_252),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_577),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_531),
.B(n_336),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_512),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_508),
.A2(n_290),
.B1(n_257),
.B2(n_259),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_502),
.B(n_244),
.Y(n_665)
);

NAND3xp33_ASAP7_75t_L g666 ( 
.A(n_577),
.B(n_580),
.C(n_503),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_483),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_576),
.B(n_260),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_576),
.B(n_293),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_568),
.B(n_263),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_568),
.B(n_341),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_524),
.B(n_336),
.Y(n_672)
);

A2O1A1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_536),
.A2(n_333),
.B(n_329),
.C(n_327),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_466),
.Y(n_674)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_578),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_459),
.A2(n_333),
.B1(n_329),
.B2(n_327),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_528),
.B(n_62),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_459),
.B(n_462),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_532),
.B(n_65),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_579),
.B(n_533),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_538),
.B(n_8),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_470),
.B(n_150),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_445),
.A2(n_145),
.B1(n_139),
.B2(n_135),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_466),
.A2(n_8),
.B1(n_10),
.B2(n_14),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_551),
.B(n_132),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_477),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_447),
.Y(n_687)
);

NOR2xp67_ASAP7_75t_L g688 ( 
.A(n_490),
.B(n_123),
.Y(n_688)
);

OR2x6_ASAP7_75t_L g689 ( 
.A(n_515),
.B(n_17),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_503),
.B(n_17),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_553),
.B(n_120),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_477),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_472),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_456),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_583),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_469),
.A2(n_113),
.B1(n_108),
.B2(n_102),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_536),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_445),
.B(n_100),
.Y(n_698)
);

AND2x4_ASAP7_75t_SL g699 ( 
.A(n_458),
.B(n_457),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_445),
.B(n_99),
.Y(n_700)
);

NAND2xp33_ASAP7_75t_L g701 ( 
.A(n_445),
.B(n_95),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_445),
.B(n_446),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_582),
.B(n_94),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_482),
.B(n_540),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_540),
.B(n_20),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_446),
.B(n_89),
.Y(n_706)
);

INVx4_ASAP7_75t_L g707 ( 
.A(n_472),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_456),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_446),
.B(n_79),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_541),
.Y(n_710)
);

NOR3xp33_ASAP7_75t_L g711 ( 
.A(n_488),
.B(n_20),
.C(n_21),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_584),
.B(n_72),
.Y(n_712)
);

NOR2xp67_ASAP7_75t_L g713 ( 
.A(n_492),
.B(n_21),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_561),
.B(n_22),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_541),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_471),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_498),
.B(n_23),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_446),
.B(n_24),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_446),
.B(n_24),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_558),
.B(n_563),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_509),
.B(n_26),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_558),
.B(n_46),
.Y(n_722)
);

OAI22xp5_ASAP7_75t_L g723 ( 
.A1(n_530),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_537),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_509),
.B(n_27),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_556),
.B(n_30),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_471),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_563),
.B(n_46),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_572),
.B(n_36),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_500),
.B(n_545),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_500),
.B(n_513),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_513),
.B(n_36),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_545),
.B(n_38),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_543),
.Y(n_734)
);

BUFx12f_ASAP7_75t_L g735 ( 
.A(n_458),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_557),
.B(n_39),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_557),
.B(n_42),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_472),
.B(n_525),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_546),
.B(n_472),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_546),
.B(n_542),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_488),
.A2(n_561),
.B1(n_468),
.B2(n_573),
.Y(n_741)
);

AO22x1_ASAP7_75t_L g742 ( 
.A1(n_514),
.A2(n_527),
.B1(n_523),
.B2(n_494),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_520),
.A2(n_526),
.B1(n_565),
.B2(n_479),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_666),
.A2(n_574),
.B(n_525),
.C(n_542),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_589),
.Y(n_745)
);

BUFx12f_ASAP7_75t_L g746 ( 
.A(n_667),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_695),
.B(n_574),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_720),
.B(n_525),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_610),
.Y(n_749)
);

OAI21xp5_ASAP7_75t_L g750 ( 
.A1(n_593),
.A2(n_550),
.B(n_444),
.Y(n_750)
);

CKINVDCx8_ASAP7_75t_R g751 ( 
.A(n_656),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_589),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_731),
.A2(n_550),
.B(n_525),
.Y(n_753)
);

HB1xp67_ASAP7_75t_L g754 ( 
.A(n_641),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_621),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_593),
.B(n_542),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_604),
.B(n_443),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_661),
.B(n_529),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_627),
.B(n_495),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_616),
.A2(n_444),
.B(n_493),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_589),
.Y(n_761)
);

NOR3xp33_ASAP7_75t_L g762 ( 
.A(n_613),
.B(n_495),
.C(n_444),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_627),
.B(n_495),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_588),
.A2(n_495),
.B(n_493),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_589),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_624),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_634),
.Y(n_767)
);

BUFx12f_ASAP7_75t_L g768 ( 
.A(n_735),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_586),
.B(n_613),
.Y(n_769)
);

CKINVDCx10_ASAP7_75t_R g770 ( 
.A(n_689),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_632),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_697),
.B(n_444),
.Y(n_772)
);

NAND2xp33_ASAP7_75t_L g773 ( 
.A(n_722),
.B(n_493),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_710),
.B(n_501),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_641),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_617),
.A2(n_738),
.B(n_707),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_704),
.B(n_501),
.Y(n_777)
);

AND2x6_ASAP7_75t_L g778 ( 
.A(n_690),
.B(n_501),
.Y(n_778)
);

NOR3xp33_ASAP7_75t_L g779 ( 
.A(n_586),
.B(n_517),
.C(n_539),
.Y(n_779)
);

NAND3xp33_ASAP7_75t_L g780 ( 
.A(n_704),
.B(n_517),
.C(n_539),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_646),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_636),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_637),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_591),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_715),
.B(n_517),
.Y(n_785)
);

NOR2xp67_ASAP7_75t_SL g786 ( 
.A(n_721),
.B(n_569),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_612),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_647),
.B(n_569),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_620),
.A2(n_590),
.B(n_609),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_592),
.B(n_614),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_699),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_693),
.A2(n_707),
.B(n_650),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_649),
.A2(n_730),
.B(n_702),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_635),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_734),
.B(n_680),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_625),
.A2(n_684),
.B1(n_657),
.B2(n_674),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_645),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_615),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_675),
.B(n_680),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_668),
.A2(n_669),
.B1(n_620),
.B2(n_743),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_599),
.A2(n_625),
.B1(n_728),
.B2(n_668),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_653),
.B(n_659),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_730),
.A2(n_618),
.B(n_701),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_671),
.B(n_606),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_SL g805 ( 
.A(n_705),
.B(n_725),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_599),
.A2(n_678),
.B(n_729),
.Y(n_806)
);

O2A1O1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_622),
.A2(n_629),
.B(n_626),
.C(n_721),
.Y(n_807)
);

INVx4_ASAP7_75t_L g808 ( 
.A(n_634),
.Y(n_808)
);

AO21x2_ASAP7_75t_L g809 ( 
.A1(n_669),
.A2(n_587),
.B(n_598),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_699),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_686),
.A2(n_692),
.B(n_587),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_665),
.B(n_651),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_615),
.Y(n_813)
);

AOI33xp33_ASAP7_75t_L g814 ( 
.A1(n_676),
.A2(n_684),
.A3(n_644),
.B1(n_602),
.B2(n_664),
.B3(n_639),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_630),
.B(n_643),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_670),
.B(n_672),
.Y(n_816)
);

NOR2xp67_ASAP7_75t_L g817 ( 
.A(n_660),
.B(n_724),
.Y(n_817)
);

NAND2x1_ASAP7_75t_L g818 ( 
.A(n_687),
.B(n_694),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_607),
.B(n_595),
.Y(n_819)
);

O2A1O1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_622),
.A2(n_629),
.B(n_626),
.C(n_678),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_608),
.B(n_585),
.Y(n_821)
);

O2A1O1Ixp5_ASAP7_75t_L g822 ( 
.A1(n_598),
.A2(n_652),
.B(n_596),
.C(n_597),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_677),
.A2(n_685),
.B(n_679),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_691),
.A2(n_716),
.B(n_727),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_708),
.A2(n_663),
.B(n_655),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_601),
.Y(n_826)
);

O2A1O1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_729),
.A2(n_674),
.B(n_657),
.C(n_705),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_608),
.B(n_662),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_600),
.B(n_681),
.Y(n_829)
);

CKINVDCx16_ASAP7_75t_R g830 ( 
.A(n_658),
.Y(n_830)
);

O2A1O1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_732),
.A2(n_733),
.B(n_726),
.C(n_725),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_605),
.Y(n_832)
);

O2A1O1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_732),
.A2(n_733),
.B(n_726),
.C(n_673),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_654),
.A2(n_706),
.B(n_698),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_741),
.A2(n_594),
.B(n_623),
.C(n_638),
.Y(n_835)
);

O2A1O1Ixp5_ASAP7_75t_L g836 ( 
.A1(n_736),
.A2(n_737),
.B(n_628),
.C(n_631),
.Y(n_836)
);

AND2x6_ASAP7_75t_L g837 ( 
.A(n_714),
.B(n_683),
.Y(n_837)
);

O2A1O1Ixp5_ASAP7_75t_SL g838 ( 
.A1(n_723),
.A2(n_682),
.B(n_703),
.C(n_712),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_700),
.A2(n_709),
.B(n_611),
.Y(n_839)
);

NOR3xp33_ASAP7_75t_L g840 ( 
.A(n_742),
.B(n_711),
.C(n_717),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_633),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_741),
.B(n_619),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_640),
.B(n_713),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_688),
.B(n_658),
.Y(n_844)
);

NOR2xp67_ASAP7_75t_L g845 ( 
.A(n_718),
.B(n_719),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_673),
.A2(n_682),
.B(n_712),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_703),
.A2(n_696),
.B(n_714),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_676),
.B(n_642),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_642),
.B(n_658),
.Y(n_849)
);

NOR3xp33_ASAP7_75t_L g850 ( 
.A(n_689),
.B(n_613),
.C(n_586),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_689),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_641),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_720),
.B(n_627),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_603),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_739),
.A2(n_506),
.B(n_740),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_593),
.A2(n_666),
.B1(n_720),
.B2(n_489),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_603),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_704),
.A2(n_720),
.B1(n_666),
.B2(n_627),
.Y(n_858)
);

AOI21x1_ASAP7_75t_L g859 ( 
.A1(n_738),
.A2(n_617),
.B(n_730),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_SL g860 ( 
.A1(n_725),
.A2(n_320),
.B1(n_335),
.B2(n_307),
.Y(n_860)
);

AOI21xp33_ASAP7_75t_L g861 ( 
.A1(n_720),
.A2(n_666),
.B(n_704),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_739),
.A2(n_506),
.B(n_740),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_695),
.B(n_593),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_603),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_739),
.A2(n_506),
.B(n_740),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_739),
.A2(n_506),
.B(n_740),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_739),
.A2(n_506),
.B(n_740),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_589),
.Y(n_868)
);

NOR2x1p5_ASAP7_75t_SL g869 ( 
.A(n_648),
.B(n_572),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_739),
.A2(n_506),
.B(n_740),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_604),
.B(n_661),
.Y(n_871)
);

O2A1O1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_593),
.A2(n_720),
.B(n_614),
.C(n_599),
.Y(n_872)
);

NAND2xp33_ASAP7_75t_L g873 ( 
.A(n_593),
.B(n_720),
.Y(n_873)
);

AND2x6_ASAP7_75t_L g874 ( 
.A(n_690),
.B(n_702),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_739),
.A2(n_506),
.B(n_740),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_720),
.B(n_627),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_604),
.B(n_661),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_604),
.B(n_661),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_593),
.A2(n_720),
.B(n_614),
.C(n_599),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_739),
.A2(n_506),
.B(n_740),
.Y(n_880)
);

A2O1A1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_666),
.A2(n_720),
.B(n_613),
.C(n_586),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_720),
.B(n_627),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_739),
.A2(n_506),
.B(n_740),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_739),
.A2(n_506),
.B(n_740),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_666),
.A2(n_720),
.B(n_613),
.C(n_586),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_604),
.B(n_453),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_603),
.Y(n_887)
);

NAND2x1p5_ASAP7_75t_L g888 ( 
.A(n_589),
.B(n_460),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_589),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_720),
.B(n_627),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_666),
.A2(n_720),
.B1(n_704),
.B2(n_599),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_720),
.B(n_627),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_739),
.A2(n_506),
.B(n_740),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_589),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_666),
.A2(n_720),
.B(n_613),
.C(n_586),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_603),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_593),
.A2(n_666),
.B1(n_720),
.B2(n_489),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_720),
.B(n_627),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_739),
.A2(n_506),
.B(n_740),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_666),
.A2(n_720),
.B(n_613),
.C(n_586),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_739),
.A2(n_506),
.B(n_740),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_593),
.A2(n_666),
.B1(n_720),
.B2(n_489),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_720),
.B(n_627),
.Y(n_903)
);

CKINVDCx6p67_ASAP7_75t_R g904 ( 
.A(n_735),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_603),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_739),
.A2(n_506),
.B(n_740),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_603),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_661),
.B(n_720),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_720),
.B(n_627),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_604),
.B(n_661),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_604),
.B(n_661),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_589),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_739),
.A2(n_506),
.B(n_740),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_589),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_739),
.A2(n_506),
.B(n_740),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_603),
.Y(n_916)
);

OAI21x1_ASAP7_75t_L g917 ( 
.A1(n_834),
.A2(n_839),
.B(n_750),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_853),
.B(n_876),
.Y(n_918)
);

BUFx2_ASAP7_75t_L g919 ( 
.A(n_775),
.Y(n_919)
);

OAI21x1_ASAP7_75t_L g920 ( 
.A1(n_750),
.A2(n_756),
.B(n_824),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_882),
.B(n_890),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_798),
.Y(n_922)
);

OAI21x1_ASAP7_75t_L g923 ( 
.A1(n_793),
.A2(n_753),
.B(n_859),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_769),
.B(n_805),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_754),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_855),
.A2(n_865),
.B(n_862),
.Y(n_926)
);

A2O1A1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_892),
.A2(n_898),
.B(n_903),
.C(n_909),
.Y(n_927)
);

INVx3_ASAP7_75t_SL g928 ( 
.A(n_791),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_861),
.A2(n_805),
.B1(n_837),
.B2(n_858),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_866),
.A2(n_870),
.B(n_867),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_795),
.B(n_812),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_799),
.B(n_782),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_761),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_881),
.A2(n_895),
.B(n_885),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_891),
.B(n_900),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_746),
.Y(n_936)
);

OAI21x1_ASAP7_75t_L g937 ( 
.A1(n_875),
.A2(n_883),
.B(n_880),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_886),
.B(n_871),
.Y(n_938)
);

OAI21x1_ASAP7_75t_SL g939 ( 
.A1(n_806),
.A2(n_847),
.B(n_827),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_877),
.B(n_878),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_813),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_783),
.B(n_816),
.Y(n_942)
);

OAI21x1_ASAP7_75t_L g943 ( 
.A1(n_884),
.A2(n_899),
.B(n_893),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_861),
.B(n_800),
.Y(n_944)
);

AOI211x1_ASAP7_75t_L g945 ( 
.A1(n_806),
.A2(n_908),
.B(n_796),
.C(n_863),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_804),
.B(n_829),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_872),
.A2(n_879),
.B(n_902),
.C(n_856),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_804),
.B(n_819),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_747),
.B(n_910),
.Y(n_949)
);

OAI21xp33_ASAP7_75t_SL g950 ( 
.A1(n_863),
.A2(n_801),
.B(n_814),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_856),
.A2(n_897),
.B(n_902),
.C(n_873),
.Y(n_951)
);

AOI21xp33_ASAP7_75t_L g952 ( 
.A1(n_807),
.A2(n_790),
.B(n_831),
.Y(n_952)
);

AND2x6_ASAP7_75t_SL g953 ( 
.A(n_758),
.B(n_757),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_901),
.A2(n_915),
.B(n_906),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_SL g955 ( 
.A(n_810),
.B(n_768),
.Y(n_955)
);

NOR3xp33_ASAP7_75t_L g956 ( 
.A(n_860),
.B(n_850),
.C(n_848),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_852),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_747),
.B(n_911),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_841),
.B(n_843),
.Y(n_959)
);

AOI21x1_ASAP7_75t_L g960 ( 
.A1(n_845),
.A2(n_777),
.B(n_913),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_748),
.A2(n_823),
.B(n_803),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_897),
.B(n_820),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_759),
.B(n_763),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_749),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_766),
.Y(n_965)
);

AO21x1_ASAP7_75t_L g966 ( 
.A1(n_842),
.A2(n_833),
.B(n_789),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_776),
.A2(n_788),
.B(n_792),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_828),
.B(n_808),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_815),
.B(n_821),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_771),
.B(n_854),
.Y(n_970)
);

OA21x2_ASAP7_75t_L g971 ( 
.A1(n_789),
.A2(n_760),
.B(n_846),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_857),
.B(n_864),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_837),
.A2(n_840),
.B1(n_817),
.B2(n_874),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_761),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_811),
.A2(n_764),
.B(n_760),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_846),
.A2(n_836),
.B(n_838),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_835),
.A2(n_796),
.B(n_822),
.C(n_905),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_744),
.A2(n_780),
.B(n_825),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_818),
.A2(n_888),
.B(n_774),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_887),
.B(n_896),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_755),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_904),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_781),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_907),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_761),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_916),
.B(n_784),
.Y(n_986)
);

NOR2xp67_ASAP7_75t_L g987 ( 
.A(n_802),
.B(n_844),
.Y(n_987)
);

AO21x1_ASAP7_75t_L g988 ( 
.A1(n_762),
.A2(n_773),
.B(n_779),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_809),
.A2(n_772),
.B(n_785),
.Y(n_989)
);

AOI21x1_ASAP7_75t_L g990 ( 
.A1(n_786),
.A2(n_826),
.B(n_832),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_745),
.A2(n_889),
.B(n_752),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_752),
.A2(n_889),
.B(n_912),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_837),
.B(n_778),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_808),
.B(n_767),
.Y(n_994)
);

AO21x1_ASAP7_75t_L g995 ( 
.A1(n_844),
.A2(n_837),
.B(n_797),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_787),
.A2(n_794),
.B(n_765),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_778),
.A2(n_874),
.B(n_849),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_765),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_767),
.B(n_851),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_765),
.A2(n_914),
.B(n_894),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_868),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_868),
.A2(n_914),
.B(n_894),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_778),
.B(n_874),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_868),
.Y(n_1004)
);

NAND2x1p5_ASAP7_75t_L g1005 ( 
.A(n_894),
.B(n_914),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_778),
.B(n_874),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_767),
.B(n_869),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_830),
.B(n_751),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_770),
.B(n_853),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_855),
.A2(n_486),
.B(n_913),
.Y(n_1010)
);

O2A1O1Ixp5_ASAP7_75t_L g1011 ( 
.A1(n_769),
.A2(n_720),
.B(n_885),
.C(n_881),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_881),
.A2(n_895),
.B(n_885),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_834),
.A2(n_839),
.B(n_750),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_881),
.A2(n_885),
.B(n_900),
.C(n_895),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_855),
.A2(n_486),
.B(n_913),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_853),
.B(n_876),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_834),
.A2(n_839),
.B(n_750),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_775),
.Y(n_1018)
);

OAI21x1_ASAP7_75t_L g1019 ( 
.A1(n_824),
.A2(n_793),
.B(n_839),
.Y(n_1019)
);

OA21x2_ASAP7_75t_L g1020 ( 
.A1(n_789),
.A2(n_760),
.B(n_806),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_886),
.B(n_604),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_853),
.B(n_876),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_798),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_886),
.B(n_604),
.Y(n_1024)
);

AOI21xp33_ASAP7_75t_L g1025 ( 
.A1(n_769),
.A2(n_613),
.B(n_586),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_881),
.A2(n_895),
.B(n_885),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_834),
.A2(n_839),
.B(n_750),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_834),
.A2(n_839),
.B(n_750),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_798),
.Y(n_1029)
);

AO31x2_ASAP7_75t_L g1030 ( 
.A1(n_856),
.A2(n_902),
.A3(n_897),
.B(n_881),
.Y(n_1030)
);

AOI21xp33_ASAP7_75t_L g1031 ( 
.A1(n_769),
.A2(n_613),
.B(n_586),
.Y(n_1031)
);

AOI22xp33_ASAP7_75t_SL g1032 ( 
.A1(n_805),
.A2(n_769),
.B1(n_613),
.B2(n_586),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_761),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_855),
.A2(n_486),
.B(n_913),
.Y(n_1034)
);

OAI21x1_ASAP7_75t_L g1035 ( 
.A1(n_834),
.A2(n_839),
.B(n_750),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_761),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_853),
.B(n_876),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_855),
.A2(n_486),
.B(n_913),
.Y(n_1038)
);

AOI21x1_ASAP7_75t_L g1039 ( 
.A1(n_845),
.A2(n_777),
.B(n_855),
.Y(n_1039)
);

AOI21xp33_ASAP7_75t_L g1040 ( 
.A1(n_769),
.A2(n_613),
.B(n_586),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_834),
.A2(n_839),
.B(n_750),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_881),
.A2(n_895),
.B(n_885),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_834),
.A2(n_839),
.B(n_750),
.Y(n_1043)
);

CKINVDCx6p67_ASAP7_75t_R g1044 ( 
.A(n_746),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_SL g1045 ( 
.A1(n_806),
.A2(n_847),
.B(n_827),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_SL g1046 ( 
.A1(n_872),
.A2(n_702),
.B(n_593),
.Y(n_1046)
);

INVxp67_ASAP7_75t_L g1047 ( 
.A(n_754),
.Y(n_1047)
);

O2A1O1Ixp5_ASAP7_75t_L g1048 ( 
.A1(n_769),
.A2(n_720),
.B(n_885),
.C(n_881),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_834),
.A2(n_839),
.B(n_750),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_775),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_834),
.A2(n_839),
.B(n_750),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_775),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_828),
.B(n_808),
.Y(n_1053)
);

CKINVDCx11_ASAP7_75t_R g1054 ( 
.A(n_768),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_881),
.A2(n_895),
.B(n_885),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_855),
.A2(n_486),
.B(n_913),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_933),
.Y(n_1057)
);

CKINVDCx8_ASAP7_75t_R g1058 ( 
.A(n_953),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_1050),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_940),
.B(n_969),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_924),
.B(n_1025),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_933),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_965),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_931),
.B(n_948),
.Y(n_1064)
);

OR2x6_ASAP7_75t_L g1065 ( 
.A(n_994),
.B(n_968),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_SL g1066 ( 
.A(n_982),
.B(n_1044),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_933),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_1032),
.A2(n_1022),
.B1(n_1037),
.B2(n_918),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_961),
.A2(n_930),
.B(n_926),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_954),
.A2(n_1012),
.B(n_934),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_942),
.B(n_949),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_919),
.Y(n_1072)
);

INVx5_ASAP7_75t_L g1073 ( 
.A(n_933),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_921),
.B(n_1016),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1026),
.A2(n_1042),
.B(n_1055),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_1018),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_1054),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_1031),
.A2(n_1040),
.B(n_927),
.C(n_946),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_929),
.B(n_924),
.Y(n_1079)
);

AND2x2_ASAP7_75t_SL g1080 ( 
.A(n_929),
.B(n_956),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_1052),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_938),
.B(n_1021),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_967),
.A2(n_1014),
.B(n_1038),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_958),
.B(n_932),
.Y(n_1084)
);

BUFx12f_ASAP7_75t_L g1085 ( 
.A(n_1054),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_970),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_972),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_980),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_982),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1010),
.A2(n_1056),
.B(n_1034),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_935),
.A2(n_944),
.B1(n_962),
.B2(n_952),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_927),
.B(n_973),
.Y(n_1092)
);

OR2x6_ASAP7_75t_L g1093 ( 
.A(n_994),
.B(n_968),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_1024),
.B(n_959),
.Y(n_1094)
);

INVx1_ASAP7_75t_SL g1095 ( 
.A(n_925),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_945),
.B(n_986),
.Y(n_1096)
);

BUFx2_ASAP7_75t_SL g1097 ( 
.A(n_987),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_986),
.B(n_963),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_1047),
.B(n_1009),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_983),
.Y(n_1100)
);

INVx5_ASAP7_75t_L g1101 ( 
.A(n_974),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_936),
.Y(n_1102)
);

BUFx12f_ASAP7_75t_L g1103 ( 
.A(n_936),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_968),
.B(n_1053),
.Y(n_1104)
);

CKINVDCx6p67_ASAP7_75t_R g1105 ( 
.A(n_928),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_974),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_1053),
.B(n_999),
.Y(n_1107)
);

AO21x1_ASAP7_75t_L g1108 ( 
.A1(n_935),
.A2(n_944),
.B(n_962),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_1011),
.A2(n_1048),
.B(n_950),
.C(n_977),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_964),
.B(n_984),
.Y(n_1110)
);

NOR3xp33_ASAP7_75t_L g1111 ( 
.A(n_951),
.B(n_947),
.C(n_1008),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_947),
.A2(n_951),
.B1(n_993),
.B2(n_981),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_957),
.B(n_941),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_941),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_928),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_939),
.A2(n_1045),
.B1(n_966),
.B2(n_995),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1008),
.B(n_985),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_955),
.A2(n_997),
.B1(n_1006),
.B2(n_1003),
.Y(n_1118)
);

BUFx2_ASAP7_75t_L g1119 ( 
.A(n_974),
.Y(n_1119)
);

NAND2x1p5_ASAP7_75t_L g1120 ( 
.A(n_1033),
.B(n_998),
.Y(n_1120)
);

NAND2x1p5_ASAP7_75t_L g1121 ( 
.A(n_1033),
.B(n_998),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_976),
.A2(n_920),
.B(n_978),
.C(n_917),
.Y(n_1122)
);

CKINVDCx6p67_ASAP7_75t_R g1123 ( 
.A(n_1033),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_922),
.B(n_1029),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_1023),
.B(n_1046),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1030),
.B(n_1023),
.Y(n_1126)
);

INVx1_ASAP7_75t_SL g1127 ( 
.A(n_1001),
.Y(n_1127)
);

OR2x6_ASAP7_75t_L g1128 ( 
.A(n_1005),
.B(n_1000),
.Y(n_1128)
);

INVx8_ASAP7_75t_L g1129 ( 
.A(n_1001),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1030),
.B(n_1004),
.Y(n_1130)
);

INVx6_ASAP7_75t_L g1131 ( 
.A(n_1005),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_1004),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_1036),
.B(n_1007),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_971),
.A2(n_1020),
.B1(n_976),
.B2(n_920),
.Y(n_1134)
);

OR2x6_ASAP7_75t_L g1135 ( 
.A(n_1002),
.B(n_996),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1030),
.B(n_971),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1020),
.B(n_960),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1039),
.B(n_988),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_991),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_979),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_979),
.Y(n_1141)
);

CKINVDCx6p67_ASAP7_75t_R g1142 ( 
.A(n_992),
.Y(n_1142)
);

INVx1_ASAP7_75t_SL g1143 ( 
.A(n_989),
.Y(n_1143)
);

BUFx8_ASAP7_75t_L g1144 ( 
.A(n_990),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_937),
.B(n_943),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_923),
.A2(n_937),
.B(n_943),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1015),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_975),
.B(n_917),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1013),
.A2(n_1017),
.B1(n_1049),
.B2(n_1027),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1013),
.B(n_1017),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_1027),
.Y(n_1151)
);

O2A1O1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1028),
.A2(n_1035),
.B(n_1041),
.C(n_1043),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_1028),
.B(n_1035),
.Y(n_1153)
);

INVx3_ASAP7_75t_SL g1154 ( 
.A(n_1041),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1043),
.A2(n_1049),
.B1(n_1051),
.B2(n_1019),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_919),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1032),
.A2(n_769),
.B1(n_805),
.B2(n_1025),
.Y(n_1157)
);

NOR2x1_ASAP7_75t_SL g1158 ( 
.A(n_993),
.B(n_809),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_933),
.Y(n_1159)
);

OAI21xp33_ASAP7_75t_L g1160 ( 
.A1(n_1025),
.A2(n_613),
.B(n_586),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_919),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_965),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_931),
.B(n_853),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_919),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_931),
.B(n_853),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_919),
.Y(n_1166)
);

INVx4_ASAP7_75t_L g1167 ( 
.A(n_933),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_968),
.B(n_1053),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_931),
.B(n_853),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_931),
.B(n_853),
.Y(n_1170)
);

OAI22x1_ASAP7_75t_L g1171 ( 
.A1(n_924),
.A2(n_858),
.B1(n_725),
.B2(n_705),
.Y(n_1171)
);

INVx5_ASAP7_75t_L g1172 ( 
.A(n_933),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_965),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1032),
.A2(n_853),
.B1(n_882),
.B2(n_876),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_919),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1032),
.B(n_769),
.Y(n_1176)
);

OR2x6_ASAP7_75t_L g1177 ( 
.A(n_994),
.B(n_642),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_931),
.B(n_853),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_931),
.B(n_853),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_1050),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_965),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_965),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1089),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1074),
.B(n_1064),
.Y(n_1184)
);

BUFx2_ASAP7_75t_SL g1185 ( 
.A(n_1115),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1111),
.B(n_1080),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_1135),
.Y(n_1187)
);

OAI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1163),
.A2(n_1178),
.B1(n_1165),
.B2(n_1179),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1161),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1063),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1071),
.B(n_1169),
.Y(n_1191)
);

OR2x6_ASAP7_75t_L g1192 ( 
.A(n_1075),
.B(n_1092),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1160),
.A2(n_1080),
.B1(n_1111),
.B2(n_1171),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_1100),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1073),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_1135),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_SL g1197 ( 
.A1(n_1061),
.A2(n_1094),
.B1(n_1115),
.B2(n_1097),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1170),
.B(n_1084),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1162),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_1161),
.Y(n_1200)
);

OR2x6_ASAP7_75t_L g1201 ( 
.A(n_1075),
.B(n_1092),
.Y(n_1201)
);

BUFx2_ASAP7_75t_R g1202 ( 
.A(n_1077),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1089),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1085),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1061),
.B(n_1060),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1146),
.A2(n_1090),
.B(n_1083),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1135),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_1166),
.Y(n_1208)
);

OAI21xp33_ASAP7_75t_L g1209 ( 
.A1(n_1157),
.A2(n_1094),
.B(n_1176),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1090),
.A2(n_1083),
.B(n_1069),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1166),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1173),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1181),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1182),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1069),
.A2(n_1152),
.B(n_1141),
.Y(n_1215)
);

OAI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1058),
.A2(n_1098),
.B1(n_1174),
.B2(n_1068),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1130),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1065),
.B(n_1093),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1157),
.B(n_1079),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1175),
.Y(n_1220)
);

NAND2x1p5_ASAP7_75t_L g1221 ( 
.A(n_1151),
.B(n_1125),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1175),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1117),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1095),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1114),
.Y(n_1225)
);

INVx3_ASAP7_75t_L g1226 ( 
.A(n_1065),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1110),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1086),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1065),
.Y(n_1229)
);

BUFx12f_ASAP7_75t_L g1230 ( 
.A(n_1103),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1082),
.B(n_1087),
.Y(n_1231)
);

AOI22x1_ASAP7_75t_L g1232 ( 
.A1(n_1070),
.A2(n_1147),
.B1(n_1139),
.B2(n_1143),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1091),
.A2(n_1088),
.B1(n_1099),
.B2(n_1096),
.Y(n_1233)
);

INVx1_ASAP7_75t_SL g1234 ( 
.A(n_1076),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1124),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1152),
.A2(n_1141),
.B(n_1155),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1091),
.A2(n_1108),
.B1(n_1125),
.B2(n_1112),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1118),
.A2(n_1156),
.B1(n_1164),
.B2(n_1116),
.Y(n_1238)
);

CKINVDCx20_ASAP7_75t_R g1239 ( 
.A(n_1105),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1155),
.A2(n_1153),
.B(n_1149),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1113),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1126),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_SL g1243 ( 
.A1(n_1066),
.A2(n_1070),
.B1(n_1072),
.B2(n_1107),
.Y(n_1243)
);

INVxp67_ASAP7_75t_SL g1244 ( 
.A(n_1072),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1133),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1107),
.A2(n_1081),
.B1(n_1104),
.B2(n_1168),
.Y(n_1246)
);

INVx4_ASAP7_75t_L g1247 ( 
.A(n_1073),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1059),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1133),
.B(n_1078),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1093),
.B(n_1168),
.Y(n_1250)
);

AOI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1104),
.A2(n_1093),
.B1(n_1177),
.B2(n_1180),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1102),
.A2(n_1158),
.B1(n_1138),
.B2(n_1144),
.Y(n_1252)
);

INVx2_ASAP7_75t_SL g1253 ( 
.A(n_1129),
.Y(n_1253)
);

CKINVDCx6p67_ASAP7_75t_R g1254 ( 
.A(n_1073),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1123),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1127),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1109),
.B(n_1116),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1177),
.B(n_1057),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1109),
.B(n_1136),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1129),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1177),
.B(n_1067),
.Y(n_1261)
);

INVx3_ASAP7_75t_SL g1262 ( 
.A(n_1129),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1144),
.Y(n_1263)
);

AO21x1_ASAP7_75t_L g1264 ( 
.A1(n_1148),
.A2(n_1137),
.B(n_1150),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1119),
.Y(n_1265)
);

AOI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1145),
.A2(n_1150),
.B(n_1128),
.Y(n_1266)
);

NAND2x1p5_ASAP7_75t_L g1267 ( 
.A(n_1073),
.B(n_1172),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1142),
.A2(n_1154),
.B1(n_1131),
.B2(n_1128),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1154),
.A2(n_1131),
.B1(n_1137),
.B2(n_1132),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1134),
.B(n_1106),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1131),
.Y(n_1271)
);

BUFx12f_ASAP7_75t_L g1272 ( 
.A(n_1062),
.Y(n_1272)
);

AOI21xp33_ASAP7_75t_SL g1273 ( 
.A1(n_1120),
.A2(n_1121),
.B(n_1122),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1132),
.Y(n_1274)
);

AOI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1122),
.A2(n_1140),
.B(n_1120),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1101),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1132),
.A2(n_1167),
.B1(n_1159),
.B2(n_1062),
.Y(n_1277)
);

NAND2x1p5_ASAP7_75t_L g1278 ( 
.A(n_1101),
.B(n_1172),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1101),
.B(n_1172),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_SL g1280 ( 
.A1(n_1167),
.A2(n_805),
.B1(n_769),
.B2(n_613),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1135),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1063),
.Y(n_1282)
);

OAI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1064),
.A2(n_805),
.B1(n_876),
.B2(n_853),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1089),
.Y(n_1284)
);

BUFx2_ASAP7_75t_R g1285 ( 
.A(n_1077),
.Y(n_1285)
);

INVx2_ASAP7_75t_SL g1286 ( 
.A(n_1220),
.Y(n_1286)
);

OR2x6_ASAP7_75t_L g1287 ( 
.A(n_1187),
.B(n_1196),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1220),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1188),
.B(n_1216),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1187),
.B(n_1196),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1206),
.A2(n_1215),
.B(n_1210),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1186),
.A2(n_1193),
.B1(n_1209),
.B2(n_1219),
.Y(n_1292)
);

INVx2_ASAP7_75t_SL g1293 ( 
.A(n_1189),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1266),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1242),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1259),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1259),
.Y(n_1297)
);

INVx1_ASAP7_75t_SL g1298 ( 
.A(n_1200),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1280),
.A2(n_1237),
.B(n_1283),
.Y(n_1299)
);

OA21x2_ASAP7_75t_L g1300 ( 
.A1(n_1236),
.A2(n_1264),
.B(n_1240),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1217),
.B(n_1186),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1270),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1217),
.B(n_1249),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1270),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1275),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1192),
.Y(n_1306)
);

OAI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1233),
.A2(n_1232),
.B(n_1184),
.Y(n_1307)
);

OR2x6_ASAP7_75t_L g1308 ( 
.A(n_1207),
.B(n_1281),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1201),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1201),
.Y(n_1310)
);

AO21x2_ASAP7_75t_L g1311 ( 
.A1(n_1273),
.A2(n_1257),
.B(n_1249),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1205),
.B(n_1191),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1223),
.B(n_1219),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1201),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1221),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1223),
.B(n_1221),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1221),
.B(n_1235),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1245),
.B(n_1198),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1225),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1228),
.B(n_1227),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1208),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1211),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1190),
.Y(n_1323)
);

INVxp67_ASAP7_75t_L g1324 ( 
.A(n_1224),
.Y(n_1324)
);

AO21x2_ASAP7_75t_L g1325 ( 
.A1(n_1199),
.A2(n_1213),
.B(n_1282),
.Y(n_1325)
);

OA21x2_ASAP7_75t_L g1326 ( 
.A1(n_1269),
.A2(n_1214),
.B(n_1212),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1222),
.Y(n_1327)
);

NAND3xp33_ASAP7_75t_L g1328 ( 
.A(n_1197),
.B(n_1238),
.C(n_1243),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1256),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_1226),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1268),
.A2(n_1231),
.B(n_1252),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1241),
.B(n_1226),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1234),
.B(n_1194),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1226),
.B(n_1229),
.Y(n_1334)
);

OR2x6_ASAP7_75t_L g1335 ( 
.A(n_1229),
.B(n_1218),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1218),
.Y(n_1336)
);

INVxp67_ASAP7_75t_L g1337 ( 
.A(n_1248),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1265),
.Y(n_1338)
);

OR2x6_ASAP7_75t_L g1339 ( 
.A(n_1218),
.B(n_1278),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1244),
.Y(n_1340)
);

INVx4_ASAP7_75t_L g1341 ( 
.A(n_1195),
.Y(n_1341)
);

BUFx8_ASAP7_75t_L g1342 ( 
.A(n_1230),
.Y(n_1342)
);

INVx5_ASAP7_75t_L g1343 ( 
.A(n_1195),
.Y(n_1343)
);

OR2x6_ASAP7_75t_L g1344 ( 
.A(n_1267),
.B(n_1278),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1326),
.Y(n_1345)
);

INVxp67_ASAP7_75t_L g1346 ( 
.A(n_1340),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1325),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1312),
.B(n_1183),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1325),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1302),
.B(n_1263),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1323),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1302),
.B(n_1263),
.Y(n_1352)
);

NOR2x1p5_ASAP7_75t_L g1353 ( 
.A(n_1328),
.B(n_1254),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1319),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1326),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1296),
.B(n_1274),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1326),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1310),
.B(n_1258),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1310),
.B(n_1261),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1296),
.B(n_1194),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1314),
.B(n_1261),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1314),
.B(n_1250),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1326),
.Y(n_1363)
);

NOR2x1_ASAP7_75t_L g1364 ( 
.A(n_1307),
.B(n_1328),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1304),
.B(n_1250),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1304),
.B(n_1185),
.Y(n_1366)
);

OAI33xp33_ASAP7_75t_L g1367 ( 
.A1(n_1289),
.A2(n_1183),
.A3(n_1284),
.B1(n_1203),
.B2(n_1255),
.B3(n_1204),
.Y(n_1367)
);

NAND2x1_ASAP7_75t_L g1368 ( 
.A(n_1287),
.B(n_1247),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1306),
.B(n_1251),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1297),
.B(n_1271),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1290),
.B(n_1271),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1295),
.B(n_1277),
.Y(n_1372)
);

OA21x2_ASAP7_75t_L g1373 ( 
.A1(n_1347),
.A2(n_1291),
.B(n_1305),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1358),
.B(n_1309),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1364),
.A2(n_1292),
.B1(n_1299),
.B2(n_1331),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_SL g1376 ( 
.A(n_1364),
.B(n_1307),
.Y(n_1376)
);

OAI21xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1353),
.A2(n_1299),
.B(n_1345),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1360),
.B(n_1321),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1360),
.B(n_1322),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1370),
.B(n_1298),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1358),
.B(n_1359),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_SL g1382 ( 
.A1(n_1353),
.A2(n_1344),
.B(n_1339),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1370),
.B(n_1298),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1358),
.B(n_1303),
.Y(n_1384)
);

NAND4xp25_ASAP7_75t_L g1385 ( 
.A(n_1372),
.B(n_1318),
.C(n_1327),
.D(n_1324),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1359),
.B(n_1303),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1366),
.B(n_1327),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1359),
.B(n_1361),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1366),
.B(n_1288),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1361),
.B(n_1316),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1361),
.B(n_1316),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1362),
.B(n_1313),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1366),
.B(n_1329),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1350),
.B(n_1313),
.Y(n_1394)
);

NOR3xp33_ASAP7_75t_L g1395 ( 
.A(n_1367),
.B(n_1331),
.C(n_1318),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1351),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1348),
.A2(n_1246),
.B1(n_1352),
.B2(n_1350),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1362),
.B(n_1301),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1350),
.B(n_1311),
.Y(n_1399)
);

NAND3xp33_ASAP7_75t_L g1400 ( 
.A(n_1345),
.B(n_1337),
.C(n_1338),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1352),
.B(n_1311),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1352),
.B(n_1311),
.Y(n_1402)
);

OA211x2_ASAP7_75t_L g1403 ( 
.A1(n_1368),
.A2(n_1333),
.B(n_1279),
.C(n_1320),
.Y(n_1403)
);

NAND3xp33_ASAP7_75t_L g1404 ( 
.A(n_1355),
.B(n_1340),
.C(n_1320),
.Y(n_1404)
);

OAI221xp5_ASAP7_75t_L g1405 ( 
.A1(n_1369),
.A2(n_1315),
.B1(n_1293),
.B2(n_1204),
.C(n_1334),
.Y(n_1405)
);

NAND2x1p5_ASAP7_75t_L g1406 ( 
.A(n_1368),
.B(n_1294),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_SL g1407 ( 
.A(n_1367),
.B(n_1202),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1365),
.B(n_1311),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1362),
.B(n_1301),
.Y(n_1409)
);

OA211x2_ASAP7_75t_L g1410 ( 
.A1(n_1372),
.A2(n_1342),
.B(n_1343),
.C(n_1344),
.Y(n_1410)
);

NOR3xp33_ASAP7_75t_L g1411 ( 
.A(n_1369),
.B(n_1315),
.C(n_1330),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1354),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1351),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_SL g1414 ( 
.A(n_1371),
.B(n_1285),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1369),
.A2(n_1339),
.B1(n_1203),
.B2(n_1284),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1365),
.B(n_1317),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1371),
.A2(n_1339),
.B1(n_1335),
.B2(n_1344),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1365),
.B(n_1286),
.Y(n_1418)
);

NOR3xp33_ASAP7_75t_L g1419 ( 
.A(n_1356),
.B(n_1330),
.C(n_1341),
.Y(n_1419)
);

OAI221xp5_ASAP7_75t_SL g1420 ( 
.A1(n_1355),
.A2(n_1332),
.B1(n_1335),
.B2(n_1339),
.C(n_1308),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_SL g1421 ( 
.A1(n_1357),
.A2(n_1336),
.B(n_1290),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1399),
.B(n_1346),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1396),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1412),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1401),
.B(n_1346),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1381),
.B(n_1357),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1402),
.B(n_1363),
.Y(n_1427)
);

AND2x2_ASAP7_75t_SL g1428 ( 
.A(n_1411),
.B(n_1363),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1376),
.B(n_1371),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1396),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1373),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1408),
.B(n_1347),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1388),
.B(n_1300),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1400),
.B(n_1349),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1413),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1373),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1412),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1374),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1406),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1389),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1406),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1404),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1406),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1392),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1404),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1400),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1394),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1392),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1380),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1390),
.B(n_1391),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1377),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1384),
.Y(n_1452)
);

INVx1_ASAP7_75t_SL g1453 ( 
.A(n_1393),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1383),
.B(n_1349),
.Y(n_1454)
);

NOR2x1p5_ASAP7_75t_L g1455 ( 
.A(n_1385),
.B(n_1336),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1384),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1375),
.B(n_1371),
.Y(n_1457)
);

OAI221xp5_ASAP7_75t_L g1458 ( 
.A1(n_1451),
.A2(n_1377),
.B1(n_1395),
.B2(n_1420),
.C(n_1421),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1427),
.B(n_1387),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1424),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1424),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1449),
.B(n_1239),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1451),
.B(n_1391),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1437),
.Y(n_1464)
);

INVx1_ASAP7_75t_SL g1465 ( 
.A(n_1453),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1427),
.B(n_1378),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1437),
.Y(n_1467)
);

INVx1_ASAP7_75t_SL g1468 ( 
.A(n_1453),
.Y(n_1468)
);

OAI31xp33_ASAP7_75t_L g1469 ( 
.A1(n_1451),
.A2(n_1405),
.A3(n_1415),
.B(n_1407),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1444),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1423),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1427),
.B(n_1379),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1423),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1430),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1430),
.Y(n_1475)
);

INVxp67_ASAP7_75t_SL g1476 ( 
.A(n_1429),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1444),
.B(n_1386),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1435),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1441),
.B(n_1419),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1444),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1449),
.B(n_1386),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1422),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1435),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1444),
.B(n_1398),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1440),
.B(n_1398),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1448),
.B(n_1409),
.Y(n_1486)
);

NAND2x1p5_ASAP7_75t_L g1487 ( 
.A(n_1441),
.B(n_1300),
.Y(n_1487)
);

INVx1_ASAP7_75t_SL g1488 ( 
.A(n_1440),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1438),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1438),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1438),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1448),
.B(n_1409),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1446),
.B(n_1416),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1448),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1432),
.B(n_1418),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1448),
.Y(n_1496)
);

INVx2_ASAP7_75t_SL g1497 ( 
.A(n_1479),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_SL g1498 ( 
.A(n_1469),
.B(n_1414),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1466),
.B(n_1446),
.Y(n_1499)
);

NAND2x1p5_ASAP7_75t_L g1500 ( 
.A(n_1465),
.B(n_1455),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1460),
.Y(n_1501)
);

NAND2xp33_ASAP7_75t_L g1502 ( 
.A(n_1468),
.B(n_1455),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1463),
.B(n_1476),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1470),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1460),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1463),
.B(n_1450),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1461),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1479),
.B(n_1450),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1479),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1482),
.B(n_1450),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1488),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1493),
.B(n_1429),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1461),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1491),
.B(n_1439),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1467),
.Y(n_1515)
);

INVxp67_ASAP7_75t_L g1516 ( 
.A(n_1462),
.Y(n_1516)
);

AOI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1458),
.A2(n_1457),
.B1(n_1403),
.B2(n_1410),
.Y(n_1517)
);

NAND3xp33_ASAP7_75t_L g1518 ( 
.A(n_1466),
.B(n_1445),
.C(n_1442),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1472),
.B(n_1422),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1472),
.B(n_1425),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_SL g1521 ( 
.A1(n_1485),
.A2(n_1457),
.B(n_1445),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1481),
.B(n_1442),
.Y(n_1522)
);

INVxp67_ASAP7_75t_L g1523 ( 
.A(n_1459),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1470),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1459),
.B(n_1454),
.Y(n_1525)
);

INVx3_ASAP7_75t_SL g1526 ( 
.A(n_1495),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1467),
.Y(n_1527)
);

OAI33xp33_ASAP7_75t_L g1528 ( 
.A1(n_1471),
.A2(n_1434),
.A3(n_1454),
.B1(n_1432),
.B2(n_1425),
.B3(n_1397),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1495),
.B(n_1447),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1480),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1477),
.B(n_1433),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1477),
.B(n_1447),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1484),
.B(n_1452),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_R g1534 ( 
.A(n_1484),
.B(n_1434),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1464),
.Y(n_1535)
);

NOR2x2_ASAP7_75t_L g1536 ( 
.A(n_1480),
.B(n_1439),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1486),
.B(n_1426),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1486),
.B(n_1426),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1492),
.B(n_1433),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1511),
.B(n_1492),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1526),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1501),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1512),
.B(n_1452),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1499),
.B(n_1494),
.Y(n_1544)
);

INVx1_ASAP7_75t_SL g1545 ( 
.A(n_1526),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1505),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1506),
.B(n_1494),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1519),
.B(n_1432),
.Y(n_1548)
);

NAND3xp33_ASAP7_75t_L g1549 ( 
.A(n_1518),
.B(n_1428),
.C(n_1342),
.Y(n_1549)
);

CKINVDCx16_ASAP7_75t_R g1550 ( 
.A(n_1498),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1503),
.Y(n_1551)
);

INVx2_ASAP7_75t_SL g1552 ( 
.A(n_1509),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1516),
.B(n_1452),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1507),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1503),
.B(n_1452),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1523),
.B(n_1456),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1506),
.B(n_1491),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1536),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1517),
.A2(n_1521),
.B1(n_1500),
.B2(n_1497),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1528),
.B(n_1230),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1536),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1508),
.B(n_1471),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1502),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1513),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1514),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1514),
.Y(n_1566)
);

INVxp67_ASAP7_75t_SL g1567 ( 
.A(n_1500),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1509),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1515),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1508),
.B(n_1473),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1527),
.Y(n_1571)
);

NOR2x1_ASAP7_75t_L g1572 ( 
.A(n_1509),
.B(n_1473),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1497),
.B(n_1474),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1510),
.Y(n_1574)
);

INVx2_ASAP7_75t_SL g1575 ( 
.A(n_1510),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1542),
.Y(n_1576)
);

AOI31xp33_ASAP7_75t_L g1577 ( 
.A1(n_1541),
.A2(n_1255),
.A3(n_1522),
.B(n_1342),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1550),
.A2(n_1502),
.B(n_1428),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1542),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1541),
.B(n_1525),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1552),
.Y(n_1581)
);

AOI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1550),
.A2(n_1428),
.B1(n_1525),
.B2(n_1403),
.Y(n_1582)
);

NOR4xp25_ASAP7_75t_SL g1583 ( 
.A(n_1567),
.B(n_1534),
.C(n_1535),
.D(n_1474),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1546),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1559),
.A2(n_1428),
.B1(n_1520),
.B2(n_1537),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1546),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1554),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1563),
.A2(n_1538),
.B1(n_1532),
.B2(n_1529),
.Y(n_1588)
);

O2A1O1Ixp33_ASAP7_75t_SL g1589 ( 
.A1(n_1560),
.A2(n_1239),
.B(n_1342),
.C(n_1475),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1554),
.Y(n_1590)
);

NAND3xp33_ASAP7_75t_L g1591 ( 
.A(n_1549),
.B(n_1524),
.C(n_1504),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1552),
.Y(n_1592)
);

INVxp67_ASAP7_75t_L g1593 ( 
.A(n_1545),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1572),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1540),
.B(n_1533),
.Y(n_1595)
);

OAI31xp33_ASAP7_75t_L g1596 ( 
.A1(n_1549),
.A2(n_1487),
.A3(n_1441),
.B(n_1443),
.Y(n_1596)
);

AOI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1545),
.A2(n_1410),
.B1(n_1417),
.B2(n_1441),
.Y(n_1597)
);

AOI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1551),
.A2(n_1441),
.B1(n_1443),
.B2(n_1439),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1564),
.Y(n_1599)
);

O2A1O1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1558),
.A2(n_1487),
.B(n_1478),
.C(n_1483),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1580),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1593),
.B(n_1574),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1593),
.B(n_1568),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1577),
.B(n_1568),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1576),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1581),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1592),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1589),
.B(n_1575),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1594),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1597),
.B(n_1575),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1588),
.B(n_1562),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1589),
.B(n_1553),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1579),
.B(n_1562),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1584),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1586),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1587),
.B(n_1570),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1595),
.B(n_1555),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1590),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1599),
.Y(n_1619)
);

AOI221xp5_ASAP7_75t_L g1620 ( 
.A1(n_1603),
.A2(n_1585),
.B1(n_1578),
.B2(n_1600),
.C(n_1591),
.Y(n_1620)
);

OAI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1611),
.A2(n_1582),
.B1(n_1578),
.B2(n_1561),
.Y(n_1621)
);

AOI221xp5_ASAP7_75t_L g1622 ( 
.A1(n_1603),
.A2(n_1600),
.B1(n_1596),
.B2(n_1558),
.C(n_1561),
.Y(n_1622)
);

AOI221xp5_ASAP7_75t_L g1623 ( 
.A1(n_1601),
.A2(n_1583),
.B1(n_1571),
.B2(n_1564),
.C(n_1569),
.Y(n_1623)
);

NAND4xp25_ASAP7_75t_L g1624 ( 
.A(n_1604),
.B(n_1572),
.C(n_1598),
.D(n_1573),
.Y(n_1624)
);

OAI211xp5_ASAP7_75t_L g1625 ( 
.A1(n_1604),
.A2(n_1571),
.B(n_1569),
.C(n_1573),
.Y(n_1625)
);

AOI221x1_ASAP7_75t_L g1626 ( 
.A1(n_1602),
.A2(n_1566),
.B1(n_1565),
.B2(n_1570),
.C(n_1556),
.Y(n_1626)
);

OAI21xp33_ASAP7_75t_L g1627 ( 
.A1(n_1610),
.A2(n_1548),
.B(n_1543),
.Y(n_1627)
);

AOI221xp5_ASAP7_75t_L g1628 ( 
.A1(n_1609),
.A2(n_1566),
.B1(n_1565),
.B2(n_1557),
.C(n_1547),
.Y(n_1628)
);

NOR2x1_ASAP7_75t_SL g1629 ( 
.A(n_1607),
.B(n_1544),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1608),
.A2(n_1548),
.B1(n_1557),
.B2(n_1544),
.Y(n_1630)
);

NOR3xp33_ASAP7_75t_L g1631 ( 
.A(n_1621),
.B(n_1606),
.C(n_1608),
.Y(n_1631)
);

NAND3xp33_ASAP7_75t_L g1632 ( 
.A(n_1623),
.B(n_1612),
.C(n_1605),
.Y(n_1632)
);

NOR3xp33_ASAP7_75t_L g1633 ( 
.A(n_1620),
.B(n_1612),
.C(n_1614),
.Y(n_1633)
);

NOR2x1_ASAP7_75t_L g1634 ( 
.A(n_1624),
.B(n_1625),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1627),
.B(n_1617),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1629),
.B(n_1613),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1630),
.B(n_1616),
.Y(n_1637)
);

AOI211xp5_ASAP7_75t_L g1638 ( 
.A1(n_1622),
.A2(n_1619),
.B(n_1618),
.C(n_1615),
.Y(n_1638)
);

XNOR2x1_ASAP7_75t_SL g1639 ( 
.A(n_1626),
.B(n_1547),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1628),
.A2(n_1557),
.B(n_1524),
.Y(n_1640)
);

NOR4xp25_ASAP7_75t_L g1641 ( 
.A(n_1632),
.B(n_1504),
.C(n_1530),
.D(n_1475),
.Y(n_1641)
);

OAI221xp5_ASAP7_75t_L g1642 ( 
.A1(n_1633),
.A2(n_1631),
.B1(n_1634),
.B2(n_1638),
.C(n_1637),
.Y(n_1642)
);

NOR2x1_ASAP7_75t_L g1643 ( 
.A(n_1636),
.B(n_1557),
.Y(n_1643)
);

AOI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1635),
.A2(n_1640),
.B1(n_1639),
.B2(n_1530),
.C(n_1514),
.Y(n_1644)
);

OAI211xp5_ASAP7_75t_SL g1645 ( 
.A1(n_1634),
.A2(n_1382),
.B(n_1478),
.C(n_1483),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1643),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1642),
.B(n_1496),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1644),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1641),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1645),
.Y(n_1650)
);

AOI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1642),
.A2(n_1539),
.B1(n_1531),
.B2(n_1439),
.Y(n_1651)
);

NAND4xp75_ASAP7_75t_L g1652 ( 
.A(n_1648),
.B(n_1539),
.C(n_1531),
.D(n_1253),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1646),
.B(n_1496),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1650),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1649),
.Y(n_1655)
);

OAI211xp5_ASAP7_75t_SL g1656 ( 
.A1(n_1651),
.A2(n_1382),
.B(n_1443),
.C(n_1490),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1654),
.Y(n_1657)
);

NAND3xp33_ASAP7_75t_SL g1658 ( 
.A(n_1655),
.B(n_1647),
.C(n_1267),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1653),
.Y(n_1659)
);

XNOR2x1_ASAP7_75t_L g1660 ( 
.A(n_1657),
.B(n_1652),
.Y(n_1660)
);

XNOR2xp5_ASAP7_75t_L g1661 ( 
.A(n_1660),
.B(n_1659),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1661),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1661),
.Y(n_1663)
);

NAND3x2_ASAP7_75t_L g1664 ( 
.A(n_1663),
.B(n_1658),
.C(n_1656),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1662),
.A2(n_1443),
.B1(n_1262),
.B2(n_1487),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1664),
.A2(n_1260),
.B(n_1489),
.Y(n_1666)
);

INVxp33_ASAP7_75t_L g1667 ( 
.A(n_1665),
.Y(n_1667)
);

OAI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1666),
.A2(n_1260),
.B(n_1443),
.Y(n_1668)
);

AOI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1668),
.A2(n_1667),
.B1(n_1262),
.B2(n_1272),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1669),
.A2(n_1272),
.B1(n_1254),
.B2(n_1436),
.Y(n_1670)
);

AOI211xp5_ASAP7_75t_L g1671 ( 
.A1(n_1670),
.A2(n_1195),
.B(n_1276),
.C(n_1431),
.Y(n_1671)
);


endmodule