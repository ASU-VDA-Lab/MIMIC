module fake_netlist_1_1229_n_1406 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1406);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1406;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_1399;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_641;
wire n_379;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_659;
wire n_386;
wire n_432;
wire n_1329;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1390;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g319 ( .A(n_41), .Y(n_319) );
INVxp67_ASAP7_75t_L g320 ( .A(n_134), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_57), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_130), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_263), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_12), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_185), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_244), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_293), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_9), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_142), .Y(n_329) );
INVxp67_ASAP7_75t_SL g330 ( .A(n_73), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_186), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_265), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_8), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_87), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_203), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_29), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_255), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_128), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_288), .Y(n_339) );
INVxp33_ASAP7_75t_SL g340 ( .A(n_200), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_34), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_164), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_239), .Y(n_343) );
CKINVDCx16_ASAP7_75t_R g344 ( .A(n_180), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_95), .Y(n_345) );
NOR2xp67_ASAP7_75t_L g346 ( .A(n_66), .B(n_90), .Y(n_346) );
CKINVDCx20_ASAP7_75t_R g347 ( .A(n_269), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_162), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_235), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_280), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_20), .Y(n_351) );
INVxp33_ASAP7_75t_L g352 ( .A(n_82), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_123), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_11), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_57), .Y(n_355) );
INVx1_ASAP7_75t_SL g356 ( .A(n_204), .Y(n_356) );
INVxp67_ASAP7_75t_SL g357 ( .A(n_78), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_136), .Y(n_358) );
INVxp33_ASAP7_75t_SL g359 ( .A(n_70), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_284), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_107), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_236), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_241), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_206), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_68), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_116), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_277), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_131), .Y(n_368) );
INVx4_ASAP7_75t_R g369 ( .A(n_222), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_84), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_313), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_223), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_189), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_315), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_301), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_286), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_209), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_184), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_215), .Y(n_379) );
BUFx2_ASAP7_75t_L g380 ( .A(n_192), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_292), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_67), .Y(n_382) );
INVxp67_ASAP7_75t_SL g383 ( .A(n_88), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_167), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_160), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_205), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_213), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_92), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_85), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_195), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_51), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_176), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_226), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_312), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_48), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_67), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_154), .Y(n_397) );
INVxp67_ASAP7_75t_SL g398 ( .A(n_190), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_40), .Y(n_399) );
INVxp67_ASAP7_75t_L g400 ( .A(n_243), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_26), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_31), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_156), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_201), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_141), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_140), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_258), .Y(n_407) );
INVxp33_ASAP7_75t_SL g408 ( .A(n_221), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_246), .Y(n_409) );
CKINVDCx16_ASAP7_75t_R g410 ( .A(n_233), .Y(n_410) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_4), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_147), .B(n_207), .Y(n_412) );
BUFx3_ASAP7_75t_L g413 ( .A(n_6), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_83), .Y(n_414) );
CKINVDCx16_ASAP7_75t_R g415 ( .A(n_31), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_251), .Y(n_416) );
BUFx2_ASAP7_75t_L g417 ( .A(n_303), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_238), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_289), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_191), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_80), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_308), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_187), .Y(n_423) );
CKINVDCx16_ASAP7_75t_R g424 ( .A(n_39), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_299), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_39), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_218), .B(n_318), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_310), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_272), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_115), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_22), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_250), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_120), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_173), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_282), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_106), .Y(n_436) );
INVx1_ASAP7_75t_SL g437 ( .A(n_135), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_12), .Y(n_438) );
CKINVDCx16_ASAP7_75t_R g439 ( .A(n_254), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_297), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_170), .Y(n_441) );
INVxp33_ASAP7_75t_L g442 ( .A(n_232), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_110), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_99), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_76), .Y(n_445) );
CKINVDCx16_ASAP7_75t_R g446 ( .A(n_9), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_79), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_117), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_300), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_317), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g451 ( .A(n_86), .Y(n_451) );
INVxp67_ASAP7_75t_L g452 ( .A(n_211), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_68), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_34), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_72), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_281), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_172), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_225), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_129), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_193), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_267), .Y(n_461) );
INVxp33_ASAP7_75t_SL g462 ( .A(n_276), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_271), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_159), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_304), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_197), .Y(n_466) );
INVxp33_ASAP7_75t_L g467 ( .A(n_126), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_51), .Y(n_468) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_29), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_0), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_91), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_74), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_114), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_234), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_256), .Y(n_475) );
CKINVDCx14_ASAP7_75t_R g476 ( .A(n_101), .Y(n_476) );
INVx1_ASAP7_75t_SL g477 ( .A(n_59), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_270), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_181), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_165), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_119), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_380), .B(n_0), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_344), .Y(n_483) );
BUFx8_ASAP7_75t_L g484 ( .A(n_417), .Y(n_484) );
AND2x4_ASAP7_75t_L g485 ( .A(n_413), .B(n_1), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_410), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_415), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_394), .B(n_1), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_439), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_424), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_389), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_372), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_352), .B(n_2), .Y(n_493) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_374), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_389), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_352), .B(n_2), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_446), .A2(n_454), .B1(n_451), .B2(n_359), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_372), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_451), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_376), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_471), .Y(n_501) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_374), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_442), .B(n_3), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_376), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_402), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_413), .B(n_5), .Y(n_506) );
INVxp67_ASAP7_75t_L g507 ( .A(n_319), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_402), .Y(n_508) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_390), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_421), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_421), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_322), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_323), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_326), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_324), .B(n_6), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_327), .Y(n_516) );
INVxp67_ASAP7_75t_L g517 ( .A(n_333), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_329), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_331), .Y(n_519) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_388), .A2(n_93), .B(n_89), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_492), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_501), .B(n_512), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_492), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_512), .B(n_442), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_494), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_494), .Y(n_526) );
INVx3_ASAP7_75t_L g527 ( .A(n_485), .Y(n_527) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_520), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_498), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_485), .B(n_334), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_498), .Y(n_531) );
CKINVDCx16_ASAP7_75t_R g532 ( .A(n_487), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_494), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_513), .B(n_467), .Y(n_534) );
AND2x4_ASAP7_75t_L g535 ( .A(n_485), .B(n_336), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_507), .B(n_467), .Y(n_536) );
AND2x6_ASAP7_75t_L g537 ( .A(n_506), .B(n_390), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_500), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_494), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_500), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_494), .Y(n_541) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_483), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_504), .Y(n_543) );
INVx4_ASAP7_75t_L g544 ( .A(n_506), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_502), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_506), .B(n_341), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_502), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_504), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_513), .B(n_320), .Y(n_549) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_520), .Y(n_550) );
AND2x4_ASAP7_75t_L g551 ( .A(n_493), .B(n_351), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_493), .B(n_354), .Y(n_552) );
INVx2_ASAP7_75t_SL g553 ( .A(n_496), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_491), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_514), .B(n_400), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_491), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_517), .B(n_325), .Y(n_557) );
INVxp67_ASAP7_75t_L g558 ( .A(n_496), .Y(n_558) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_520), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_514), .B(n_365), .Y(n_560) );
AND2x4_ASAP7_75t_L g561 ( .A(n_516), .B(n_370), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_515), .A2(n_401), .B1(n_414), .B2(n_396), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_516), .B(n_426), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_490), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_495), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_518), .B(n_454), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_515), .A2(n_438), .B1(n_445), .B2(n_431), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_518), .A2(n_453), .B1(n_455), .B2(n_447), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_534), .B(n_519), .Y(n_569) );
NAND3xp33_ASAP7_75t_SL g570 ( .A(n_562), .B(n_382), .C(n_321), .Y(n_570) );
CKINVDCx11_ASAP7_75t_R g571 ( .A(n_564), .Y(n_571) );
INVxp67_ASAP7_75t_L g572 ( .A(n_553), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_554), .Y(n_573) );
BUFx3_ASAP7_75t_L g574 ( .A(n_537), .Y(n_574) );
INVx3_ASAP7_75t_L g575 ( .A(n_544), .Y(n_575) );
BUFx3_ASAP7_75t_L g576 ( .A(n_537), .Y(n_576) );
NAND2xp33_ASAP7_75t_L g577 ( .A(n_537), .B(n_483), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_524), .B(n_503), .Y(n_578) );
CKINVDCx11_ASAP7_75t_R g579 ( .A(n_532), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_554), .Y(n_580) );
INVx5_ASAP7_75t_L g581 ( .A(n_537), .Y(n_581) );
NOR3xp33_ASAP7_75t_SL g582 ( .A(n_532), .B(n_489), .C(n_486), .Y(n_582) );
BUFx2_ASAP7_75t_L g583 ( .A(n_542), .Y(n_583) );
INVx5_ASAP7_75t_L g584 ( .A(n_537), .Y(n_584) );
OR2x6_ASAP7_75t_L g585 ( .A(n_553), .B(n_499), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_558), .B(n_482), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_566), .B(n_522), .Y(n_587) );
NOR2xp67_ASAP7_75t_L g588 ( .A(n_536), .B(n_497), .Y(n_588) );
NAND3xp33_ASAP7_75t_SL g589 ( .A(n_567), .B(n_395), .C(n_391), .Y(n_589) );
AND2x4_ASAP7_75t_L g590 ( .A(n_551), .B(n_488), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_556), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_551), .A2(n_489), .B1(n_486), .B2(n_484), .Y(n_592) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_551), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_556), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_552), .Y(n_595) );
CKINVDCx16_ASAP7_75t_R g596 ( .A(n_552), .Y(n_596) );
INVx2_ASAP7_75t_SL g597 ( .A(n_552), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_560), .B(n_484), .Y(n_598) );
BUFx3_ASAP7_75t_L g599 ( .A(n_537), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_565), .Y(n_600) );
INVx4_ASAP7_75t_L g601 ( .A(n_537), .Y(n_601) );
NOR2x2_ASAP7_75t_L g602 ( .A(n_544), .B(n_484), .Y(n_602) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_528), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_565), .Y(n_604) );
AND2x4_ASAP7_75t_L g605 ( .A(n_561), .B(n_510), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_568), .B(n_477), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_560), .B(n_325), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_521), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_523), .Y(n_609) );
INVxp33_ASAP7_75t_L g610 ( .A(n_549), .Y(n_610) );
INVx2_ASAP7_75t_SL g611 ( .A(n_530), .Y(n_611) );
BUFx4f_ASAP7_75t_L g612 ( .A(n_530), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_523), .Y(n_613) );
BUFx3_ASAP7_75t_L g614 ( .A(n_530), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_529), .Y(n_615) );
NOR3xp33_ASAP7_75t_SL g616 ( .A(n_557), .B(n_345), .C(n_339), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_525), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_529), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_531), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_527), .B(n_332), .Y(n_620) );
AND2x4_ASAP7_75t_L g621 ( .A(n_561), .B(n_347), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_527), .B(n_335), .Y(n_622) );
INVx3_ASAP7_75t_SL g623 ( .A(n_560), .Y(n_623) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_530), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_560), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_535), .B(n_340), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_531), .Y(n_627) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_528), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_538), .Y(n_629) );
INVx3_ASAP7_75t_L g630 ( .A(n_527), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_538), .Y(n_631) );
OR2x6_ASAP7_75t_L g632 ( .A(n_535), .B(n_355), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_535), .B(n_337), .Y(n_633) );
NOR2x1p5_ASAP7_75t_L g634 ( .A(n_561), .B(n_330), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_563), .B(n_339), .Y(n_635) );
INVxp67_ASAP7_75t_L g636 ( .A(n_563), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_563), .B(n_345), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_540), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_563), .B(n_371), .Y(n_639) );
NOR2x2_ASAP7_75t_L g640 ( .A(n_535), .B(n_328), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_540), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_543), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_555), .B(n_371), .Y(n_643) );
INVxp67_ASAP7_75t_SL g644 ( .A(n_543), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_546), .B(n_378), .Y(n_645) );
NAND2x1_ASAP7_75t_L g646 ( .A(n_546), .B(n_369), .Y(n_646) );
INVx2_ASAP7_75t_SL g647 ( .A(n_546), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_548), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_546), .B(n_357), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_548), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_528), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_528), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_528), .A2(n_359), .B1(n_505), .B2(n_495), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_550), .B(n_378), .Y(n_654) );
NAND2x1p5_ASAP7_75t_L g655 ( .A(n_550), .B(n_468), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_550), .Y(n_656) );
INVxp67_ASAP7_75t_SL g657 ( .A(n_550), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_559), .Y(n_658) );
XNOR2xp5_ASAP7_75t_L g659 ( .A(n_525), .B(n_328), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_526), .Y(n_660) );
INVx1_ASAP7_75t_SL g661 ( .A(n_559), .Y(n_661) );
NOR2xp33_ASAP7_75t_SL g662 ( .A(n_601), .B(n_347), .Y(n_662) );
INVx2_ASAP7_75t_SL g663 ( .A(n_596), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_587), .B(n_340), .Y(n_664) );
O2A1O1Ixp33_ASAP7_75t_L g665 ( .A1(n_593), .A2(n_469), .B(n_472), .C(n_470), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_621), .B(n_411), .Y(n_666) );
O2A1O1Ixp33_ASAP7_75t_L g667 ( .A1(n_593), .A2(n_508), .B(n_511), .C(n_505), .Y(n_667) );
OR2x2_ASAP7_75t_L g668 ( .A(n_583), .B(n_621), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_625), .A2(n_384), .B1(n_418), .B2(n_397), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_657), .A2(n_559), .B(n_520), .Y(n_670) );
AO22x1_ASAP7_75t_L g671 ( .A1(n_602), .A2(n_462), .B1(n_408), .B2(n_441), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_636), .A2(n_384), .B1(n_418), .B2(n_397), .Y(n_672) );
A2O1A1Ixp33_ASAP7_75t_L g673 ( .A1(n_573), .A2(n_559), .B(n_346), .C(n_511), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_644), .Y(n_674) );
BUFx2_ASAP7_75t_L g675 ( .A(n_632), .Y(n_675) );
INVx5_ASAP7_75t_L g676 ( .A(n_601), .Y(n_676) );
BUFx3_ASAP7_75t_L g677 ( .A(n_579), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_644), .Y(n_678) );
AND2x4_ASAP7_75t_L g679 ( .A(n_595), .B(n_433), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_598), .B(n_408), .Y(n_680) );
NOR2xp33_ASAP7_75t_SL g681 ( .A(n_574), .B(n_433), .Y(n_681) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_574), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_597), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_630), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_636), .A2(n_481), .B1(n_480), .B2(n_462), .Y(n_685) );
BUFx3_ASAP7_75t_L g686 ( .A(n_579), .Y(n_686) );
INVx3_ASAP7_75t_L g687 ( .A(n_575), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_630), .Y(n_688) );
INVx4_ASAP7_75t_L g689 ( .A(n_623), .Y(n_689) );
INVx4_ASAP7_75t_L g690 ( .A(n_623), .Y(n_690) );
A2O1A1Ixp33_ASAP7_75t_L g691 ( .A1(n_594), .A2(n_559), .B(n_508), .C(n_342), .Y(n_691) );
OR2x2_ASAP7_75t_L g692 ( .A(n_659), .B(n_411), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_575), .Y(n_693) );
A2O1A1Ixp33_ASAP7_75t_L g694 ( .A1(n_580), .A2(n_343), .B(n_348), .C(n_338), .Y(n_694) );
CKINVDCx5p33_ASAP7_75t_R g695 ( .A(n_571), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_591), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_614), .Y(n_697) );
BUFx12f_ASAP7_75t_L g698 ( .A(n_571), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_605), .Y(n_699) );
O2A1O1Ixp5_ASAP7_75t_L g700 ( .A1(n_578), .A2(n_633), .B(n_646), .C(n_622), .Y(n_700) );
AND2x4_ASAP7_75t_SL g701 ( .A(n_632), .B(n_480), .Y(n_701) );
INVx1_ASAP7_75t_SL g702 ( .A(n_581), .Y(n_702) );
BUFx3_ASAP7_75t_L g703 ( .A(n_590), .Y(n_703) );
A2O1A1Ixp33_ASAP7_75t_L g704 ( .A1(n_600), .A2(n_350), .B(n_358), .C(n_349), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_605), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_582), .Y(n_706) );
CKINVDCx5p33_ASAP7_75t_R g707 ( .A(n_582), .Y(n_707) );
NOR2x1_ASAP7_75t_L g708 ( .A(n_570), .B(n_481), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_569), .B(n_420), .Y(n_709) );
AND2x4_ASAP7_75t_L g710 ( .A(n_590), .B(n_383), .Y(n_710) );
AND2x6_ASAP7_75t_L g711 ( .A(n_576), .B(n_360), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_586), .B(n_420), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_572), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_604), .Y(n_714) );
INVx3_ASAP7_75t_L g715 ( .A(n_576), .Y(n_715) );
INVx6_ASAP7_75t_L g716 ( .A(n_634), .Y(n_716) );
BUFx2_ASAP7_75t_L g717 ( .A(n_632), .Y(n_717) );
INVxp67_ASAP7_75t_L g718 ( .A(n_607), .Y(n_718) );
AOI21x1_ASAP7_75t_L g719 ( .A1(n_651), .A2(n_533), .B(n_526), .Y(n_719) );
INVx5_ASAP7_75t_L g720 ( .A(n_581), .Y(n_720) );
AOI22xp33_ASAP7_75t_SL g721 ( .A1(n_624), .A2(n_476), .B1(n_441), .B2(n_457), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_626), .B(n_449), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_608), .Y(n_723) );
NAND2x2_ASAP7_75t_L g724 ( .A(n_602), .B(n_427), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_612), .A2(n_476), .B1(n_449), .B2(n_461), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g726 ( .A1(n_657), .A2(n_539), .B(n_533), .Y(n_726) );
BUFx8_ASAP7_75t_SL g727 ( .A(n_585), .Y(n_727) );
BUFx2_ASAP7_75t_SL g728 ( .A(n_581), .Y(n_728) );
NAND2x1_ASAP7_75t_SL g729 ( .A(n_592), .B(n_361), .Y(n_729) );
O2A1O1Ixp33_ASAP7_75t_L g730 ( .A1(n_570), .A2(n_452), .B(n_362), .C(n_364), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_613), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_572), .Y(n_732) );
NOR2xp67_ASAP7_75t_L g733 ( .A(n_584), .B(n_94), .Y(n_733) );
INVx4_ASAP7_75t_L g734 ( .A(n_584), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_626), .B(n_461), .Y(n_735) );
CKINVDCx5p33_ASAP7_75t_R g736 ( .A(n_616), .Y(n_736) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_612), .Y(n_737) );
AOI21xp5_ASAP7_75t_L g738 ( .A1(n_654), .A2(n_541), .B(n_539), .Y(n_738) );
AO21x2_ASAP7_75t_L g739 ( .A1(n_652), .A2(n_366), .B(n_363), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_585), .A2(n_398), .B1(n_367), .B2(n_373), .Y(n_740) );
NAND2x1p5_ASAP7_75t_L g741 ( .A(n_584), .B(n_399), .Y(n_741) );
BUFx12f_ASAP7_75t_L g742 ( .A(n_585), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_619), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_638), .Y(n_744) );
BUFx6f_ASAP7_75t_L g745 ( .A(n_599), .Y(n_745) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_611), .Y(n_746) );
BUFx8_ASAP7_75t_L g747 ( .A(n_649), .Y(n_747) );
INVx3_ASAP7_75t_L g748 ( .A(n_599), .Y(n_748) );
AND2x4_ASAP7_75t_L g749 ( .A(n_647), .B(n_588), .Y(n_749) );
OAI21xp5_ASAP7_75t_L g750 ( .A1(n_656), .A2(n_547), .B(n_545), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g751 ( .A(n_616), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_610), .B(n_464), .Y(n_752) );
O2A1O1Ixp33_ASAP7_75t_L g753 ( .A1(n_589), .A2(n_368), .B(n_377), .C(n_375), .Y(n_753) );
NAND2xp33_ASAP7_75t_L g754 ( .A(n_655), .B(n_464), .Y(n_754) );
INVx1_ASAP7_75t_SL g755 ( .A(n_640), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_641), .Y(n_756) );
NOR3xp33_ASAP7_75t_L g757 ( .A(n_589), .B(n_474), .C(n_465), .Y(n_757) );
INVx1_ASAP7_75t_SL g758 ( .A(n_640), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_610), .A2(n_399), .B1(n_509), .B2(n_502), .Y(n_759) );
INVx3_ASAP7_75t_L g760 ( .A(n_648), .Y(n_760) );
AND2x4_ASAP7_75t_L g761 ( .A(n_633), .B(n_379), .Y(n_761) );
BUFx3_ASAP7_75t_L g762 ( .A(n_650), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_606), .B(n_465), .Y(n_763) );
O2A1O1Ixp5_ASAP7_75t_L g764 ( .A1(n_620), .A2(n_388), .B(n_385), .C(n_386), .Y(n_764) );
AOI21xp5_ASAP7_75t_L g765 ( .A1(n_658), .A2(n_387), .B(n_381), .Y(n_765) );
CKINVDCx10_ASAP7_75t_R g766 ( .A(n_577), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_643), .B(n_474), .Y(n_767) );
INVx2_ASAP7_75t_SL g768 ( .A(n_635), .Y(n_768) );
OAI22xp33_ASAP7_75t_L g769 ( .A1(n_637), .A2(n_475), .B1(n_399), .B2(n_393), .Y(n_769) );
INVx3_ASAP7_75t_L g770 ( .A(n_609), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_639), .B(n_475), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_615), .Y(n_772) );
BUFx12f_ASAP7_75t_L g773 ( .A(n_655), .Y(n_773) );
INVx3_ASAP7_75t_L g774 ( .A(n_618), .Y(n_774) );
NAND2xp5_ASAP7_75t_SL g775 ( .A(n_645), .B(n_353), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_627), .Y(n_776) );
INVx3_ASAP7_75t_L g777 ( .A(n_629), .Y(n_777) );
BUFx2_ASAP7_75t_L g778 ( .A(n_631), .Y(n_778) );
AND3x1_ASAP7_75t_SL g779 ( .A(n_642), .B(n_403), .C(n_392), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_653), .A2(n_399), .B1(n_509), .B2(n_502), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_617), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_653), .A2(n_509), .B1(n_404), .B2(n_406), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_620), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_617), .Y(n_784) );
INVxp67_ASAP7_75t_SL g785 ( .A(n_603), .Y(n_785) );
A2O1A1Ixp33_ASAP7_75t_L g786 ( .A1(n_661), .A2(n_405), .B(n_409), .C(n_407), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_603), .A2(n_416), .B1(n_422), .B2(n_419), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_603), .B(n_356), .Y(n_788) );
INVx4_ASAP7_75t_L g789 ( .A(n_628), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_660), .Y(n_790) );
OAI21xp5_ASAP7_75t_L g791 ( .A1(n_660), .A2(n_425), .B(n_423), .Y(n_791) );
A2O1A1Ixp33_ASAP7_75t_SL g792 ( .A1(n_628), .A2(n_412), .B(n_429), .C(n_428), .Y(n_792) );
BUFx6f_ASAP7_75t_L g793 ( .A(n_628), .Y(n_793) );
INVx4_ASAP7_75t_L g794 ( .A(n_628), .Y(n_794) );
BUFx12f_ASAP7_75t_L g795 ( .A(n_579), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_598), .B(n_437), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_585), .A2(n_509), .B1(n_432), .B2(n_434), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_625), .A2(n_435), .B1(n_436), .B2(n_430), .Y(n_798) );
INVx3_ASAP7_75t_L g799 ( .A(n_575), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_593), .Y(n_800) );
NAND3xp33_ASAP7_75t_L g801 ( .A(n_757), .B(n_509), .C(n_443), .Y(n_801) );
OA21x2_ASAP7_75t_L g802 ( .A1(n_673), .A2(n_479), .B(n_444), .Y(n_802) );
AO21x2_ASAP7_75t_L g803 ( .A1(n_691), .A2(n_448), .B(n_440), .Y(n_803) );
OAI21x1_ASAP7_75t_L g804 ( .A1(n_719), .A2(n_456), .B(n_450), .Y(n_804) );
INVx2_ASAP7_75t_L g805 ( .A(n_781), .Y(n_805) );
NAND2xp5_ASAP7_75t_SL g806 ( .A(n_662), .B(n_458), .Y(n_806) );
OAI21x1_ASAP7_75t_L g807 ( .A1(n_738), .A2(n_460), .B(n_459), .Y(n_807) );
BUFx2_ASAP7_75t_L g808 ( .A(n_773), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_713), .Y(n_809) );
INVxp67_ASAP7_75t_L g810 ( .A(n_662), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_732), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_701), .B(n_7), .Y(n_812) );
OAI21x1_ASAP7_75t_SL g813 ( .A1(n_791), .A2(n_466), .B(n_463), .Y(n_813) );
INVx1_ASAP7_75t_SL g814 ( .A(n_675), .Y(n_814) );
INVx2_ASAP7_75t_L g815 ( .A(n_790), .Y(n_815) );
AOI21xp33_ASAP7_75t_SL g816 ( .A1(n_695), .A2(n_7), .B(n_8), .Y(n_816) );
INVxp67_ASAP7_75t_SL g817 ( .A(n_681), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_778), .Y(n_818) );
AO31x2_ASAP7_75t_L g819 ( .A1(n_786), .A2(n_473), .A3(n_13), .B(n_10), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_718), .B(n_10), .Y(n_820) );
OA21x2_ASAP7_75t_L g821 ( .A1(n_750), .A2(n_478), .B(n_97), .Y(n_821) );
AO21x2_ASAP7_75t_L g822 ( .A1(n_739), .A2(n_98), .B(n_96), .Y(n_822) );
OAI21x1_ASAP7_75t_L g823 ( .A1(n_726), .A2(n_102), .B(n_100), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_800), .Y(n_824) );
BUFx3_ASAP7_75t_L g825 ( .A(n_689), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_674), .A2(n_14), .B1(n_11), .B2(n_13), .Y(n_826) );
OAI21xp5_ASAP7_75t_L g827 ( .A1(n_765), .A2(n_104), .B(n_103), .Y(n_827) );
OR2x2_ASAP7_75t_L g828 ( .A(n_692), .B(n_14), .Y(n_828) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_678), .Y(n_829) );
INVx1_ASAP7_75t_SL g830 ( .A(n_717), .Y(n_830) );
NAND2x1p5_ASAP7_75t_L g831 ( .A(n_689), .B(n_15), .Y(n_831) );
OAI21x1_ASAP7_75t_L g832 ( .A1(n_785), .A2(n_108), .B(n_105), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_770), .Y(n_833) );
BUFx3_ASAP7_75t_L g834 ( .A(n_690), .Y(n_834) );
O2A1O1Ixp33_ASAP7_75t_L g835 ( .A1(n_694), .A2(n_15), .B(n_16), .C(n_17), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_795), .Y(n_836) );
AO21x2_ASAP7_75t_L g837 ( .A1(n_739), .A2(n_111), .B(n_109), .Y(n_837) );
INVx2_ASAP7_75t_L g838 ( .A(n_770), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_742), .A2(n_776), .B1(n_772), .B2(n_768), .Y(n_839) );
BUFx2_ASAP7_75t_L g840 ( .A(n_747), .Y(n_840) );
OAI22xp33_ASAP7_75t_L g841 ( .A1(n_681), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_841) );
AO31x2_ASAP7_75t_L g842 ( .A1(n_704), .A2(n_18), .A3(n_19), .B(n_20), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_699), .Y(n_843) );
NOR2xp67_ASAP7_75t_L g844 ( .A(n_698), .B(n_19), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_774), .Y(n_845) );
OAI21x1_ASAP7_75t_L g846 ( .A1(n_700), .A2(n_113), .B(n_112), .Y(n_846) );
OAI21x1_ASAP7_75t_L g847 ( .A1(n_733), .A2(n_121), .B(n_118), .Y(n_847) );
OAI21x1_ASAP7_75t_L g848 ( .A1(n_733), .A2(n_124), .B(n_122), .Y(n_848) );
BUFx10_ASAP7_75t_L g849 ( .A(n_679), .Y(n_849) );
INVx2_ASAP7_75t_SL g850 ( .A(n_677), .Y(n_850) );
CKINVDCx16_ASAP7_75t_R g851 ( .A(n_686), .Y(n_851) );
AND2x4_ASAP7_75t_L g852 ( .A(n_749), .B(n_21), .Y(n_852) );
INVx3_ASAP7_75t_L g853 ( .A(n_690), .Y(n_853) );
INVx2_ASAP7_75t_SL g854 ( .A(n_747), .Y(n_854) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_664), .B(n_680), .Y(n_855) );
AOI21x1_ASAP7_75t_L g856 ( .A1(n_791), .A2(n_127), .B(n_125), .Y(n_856) );
CKINVDCx16_ASAP7_75t_R g857 ( .A(n_669), .Y(n_857) );
NAND2xp33_ASAP7_75t_SL g858 ( .A(n_793), .B(n_21), .Y(n_858) );
OAI21x1_ASAP7_75t_L g859 ( .A1(n_741), .A2(n_133), .B(n_132), .Y(n_859) );
INVx2_ASAP7_75t_L g860 ( .A(n_774), .Y(n_860) );
OR2x6_ASAP7_75t_L g861 ( .A(n_679), .B(n_22), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_705), .Y(n_862) );
AO21x2_ASAP7_75t_L g863 ( .A1(n_792), .A2(n_138), .B(n_137), .Y(n_863) );
OAI21xp5_ASAP7_75t_L g864 ( .A1(n_783), .A2(n_143), .B(n_139), .Y(n_864) );
INVx2_ASAP7_75t_SL g865 ( .A(n_716), .Y(n_865) );
BUFx5_ASAP7_75t_L g866 ( .A(n_711), .Y(n_866) );
OAI22xp33_ASAP7_75t_SL g867 ( .A1(n_669), .A2(n_23), .B1(n_24), .B2(n_25), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_683), .Y(n_868) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_685), .A2(n_23), .B1(n_24), .B2(n_26), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_740), .B(n_27), .Y(n_870) );
BUFx12f_ASAP7_75t_L g871 ( .A(n_663), .Y(n_871) );
OAI21x1_ASAP7_75t_L g872 ( .A1(n_777), .A2(n_145), .B(n_144), .Y(n_872) );
AO21x2_ASAP7_75t_L g873 ( .A1(n_787), .A2(n_148), .B(n_146), .Y(n_873) );
OAI21x1_ASAP7_75t_L g874 ( .A1(n_777), .A2(n_150), .B(n_149), .Y(n_874) );
AO21x2_ASAP7_75t_L g875 ( .A1(n_787), .A2(n_152), .B(n_151), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_703), .Y(n_876) );
INVx2_ASAP7_75t_L g877 ( .A(n_784), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_740), .B(n_763), .Y(n_878) );
OA21x2_ASAP7_75t_L g879 ( .A1(n_764), .A2(n_155), .B(n_153), .Y(n_879) );
OAI21xp5_ASAP7_75t_L g880 ( .A1(n_696), .A2(n_714), .B(n_723), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_762), .Y(n_881) );
OA21x2_ASAP7_75t_L g882 ( .A1(n_759), .A2(n_158), .B(n_157), .Y(n_882) );
AOI21xp33_ASAP7_75t_L g883 ( .A1(n_752), .A2(n_27), .B(n_28), .Y(n_883) );
OAI21x1_ASAP7_75t_L g884 ( .A1(n_780), .A2(n_163), .B(n_161), .Y(n_884) );
OR2x6_ASAP7_75t_L g885 ( .A(n_671), .B(n_28), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_731), .Y(n_886) );
AOI21xp33_ASAP7_75t_L g887 ( .A1(n_796), .A2(n_30), .B(n_32), .Y(n_887) );
OAI21x1_ASAP7_75t_L g888 ( .A1(n_760), .A2(n_168), .B(n_166), .Y(n_888) );
NOR2xp33_ASAP7_75t_L g889 ( .A(n_668), .B(n_30), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_743), .Y(n_890) );
NOR2x1_ASAP7_75t_L g891 ( .A(n_706), .B(n_32), .Y(n_891) );
OAI21x1_ASAP7_75t_L g892 ( .A1(n_760), .A2(n_171), .B(n_169), .Y(n_892) );
AND2x4_ASAP7_75t_L g893 ( .A(n_749), .B(n_33), .Y(n_893) );
O2A1O1Ixp5_ASAP7_75t_L g894 ( .A1(n_788), .A2(n_199), .B(n_314), .C(n_311), .Y(n_894) );
CKINVDCx20_ASAP7_75t_R g895 ( .A(n_727), .Y(n_895) );
INVx3_ASAP7_75t_L g896 ( .A(n_676), .Y(n_896) );
XNOR2xp5_ASAP7_75t_L g897 ( .A(n_685), .B(n_33), .Y(n_897) );
INVx1_ASAP7_75t_SL g898 ( .A(n_716), .Y(n_898) );
CKINVDCx20_ASAP7_75t_R g899 ( .A(n_779), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_709), .B(n_35), .Y(n_900) );
OA21x2_ASAP7_75t_L g901 ( .A1(n_797), .A2(n_198), .B(n_309), .Y(n_901) );
OAI21x1_ASAP7_75t_L g902 ( .A1(n_744), .A2(n_196), .B(n_307), .Y(n_902) );
OAI21x1_ASAP7_75t_L g903 ( .A1(n_756), .A2(n_194), .B(n_306), .Y(n_903) );
NAND2xp5_ASAP7_75t_SL g904 ( .A(n_789), .B(n_174), .Y(n_904) );
BUFx4f_ASAP7_75t_L g905 ( .A(n_711), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_761), .A2(n_35), .B1(n_36), .B2(n_37), .Y(n_906) );
OAI21x1_ASAP7_75t_L g907 ( .A1(n_667), .A2(n_202), .B(n_305), .Y(n_907) );
HB1xp67_ASAP7_75t_L g908 ( .A(n_676), .Y(n_908) );
BUFx12f_ASAP7_75t_L g909 ( .A(n_707), .Y(n_909) );
BUFx2_ASAP7_75t_L g910 ( .A(n_711), .Y(n_910) );
BUFx2_ASAP7_75t_L g911 ( .A(n_711), .Y(n_911) );
OAI21x1_ASAP7_75t_L g912 ( .A1(n_688), .A2(n_188), .B(n_302), .Y(n_912) );
INVx3_ASAP7_75t_L g913 ( .A(n_676), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_746), .Y(n_914) );
OAI21x1_ASAP7_75t_L g915 ( .A1(n_684), .A2(n_183), .B(n_298), .Y(n_915) );
OAI21x1_ASAP7_75t_L g916 ( .A1(n_782), .A2(n_182), .B(n_296), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_708), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_917) );
INVx1_ASAP7_75t_SL g918 ( .A(n_666), .Y(n_918) );
A2O1A1Ixp33_ASAP7_75t_L g919 ( .A1(n_730), .A2(n_38), .B(n_40), .C(n_41), .Y(n_919) );
OAI21x1_ASAP7_75t_L g920 ( .A1(n_687), .A2(n_212), .B(n_295), .Y(n_920) );
BUFx12f_ASAP7_75t_L g921 ( .A(n_736), .Y(n_921) );
OAI21xp5_ASAP7_75t_L g922 ( .A1(n_722), .A2(n_210), .B(n_294), .Y(n_922) );
NOR2x1_ASAP7_75t_R g923 ( .A(n_751), .B(n_42), .Y(n_923) );
CKINVDCx5p33_ASAP7_75t_R g924 ( .A(n_766), .Y(n_924) );
AO21x2_ASAP7_75t_L g925 ( .A1(n_754), .A2(n_208), .B(n_291), .Y(n_925) );
OR2x6_ASAP7_75t_L g926 ( .A(n_737), .B(n_42), .Y(n_926) );
OAI21x1_ASAP7_75t_L g927 ( .A1(n_687), .A2(n_179), .B(n_290), .Y(n_927) );
OAI21x1_ASAP7_75t_L g928 ( .A1(n_715), .A2(n_178), .B(n_287), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_712), .B(n_43), .Y(n_929) );
BUFx4f_ASAP7_75t_L g930 ( .A(n_710), .Y(n_930) );
OAI21x1_ASAP7_75t_L g931 ( .A1(n_799), .A2(n_177), .B(n_285), .Y(n_931) );
AND2x2_ASAP7_75t_L g932 ( .A(n_755), .B(n_43), .Y(n_932) );
AO21x2_ASAP7_75t_L g933 ( .A1(n_798), .A2(n_214), .B(n_283), .Y(n_933) );
AO21x2_ASAP7_75t_L g934 ( .A1(n_769), .A2(n_175), .B(n_279), .Y(n_934) );
HB1xp67_ASAP7_75t_L g935 ( .A(n_682), .Y(n_935) );
AND2x2_ASAP7_75t_L g936 ( .A(n_755), .B(n_44), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_710), .B(n_44), .Y(n_937) );
OAI21xp5_ASAP7_75t_L g938 ( .A1(n_735), .A2(n_247), .B(n_278), .Y(n_938) );
OAI21xp5_ASAP7_75t_L g939 ( .A1(n_771), .A2(n_245), .B(n_275), .Y(n_939) );
OAI21xp5_ASAP7_75t_L g940 ( .A1(n_693), .A2(n_242), .B(n_274), .Y(n_940) );
OAI21x1_ASAP7_75t_L g941 ( .A1(n_799), .A2(n_316), .B(n_273), .Y(n_941) );
AND2x2_ASAP7_75t_L g942 ( .A(n_758), .B(n_45), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_758), .B(n_721), .Y(n_943) );
OAI21x1_ASAP7_75t_L g944 ( .A1(n_715), .A2(n_268), .B(n_266), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_665), .B(n_45), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_725), .B(n_46), .Y(n_946) );
BUFx3_ASAP7_75t_L g947 ( .A(n_720), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_697), .Y(n_948) );
OAI21xp5_ASAP7_75t_L g949 ( .A1(n_767), .A2(n_264), .B(n_262), .Y(n_949) );
OAI21x1_ASAP7_75t_L g950 ( .A1(n_748), .A2(n_261), .B(n_260), .Y(n_950) );
OAI222xp33_ASAP7_75t_L g951 ( .A1(n_766), .A2(n_46), .B1(n_47), .B2(n_48), .C1(n_49), .C2(n_50), .Y(n_951) );
AND2x2_ASAP7_75t_L g952 ( .A(n_775), .B(n_47), .Y(n_952) );
OAI21x1_ASAP7_75t_L g953 ( .A1(n_748), .A2(n_259), .B(n_257), .Y(n_953) );
INVx2_ASAP7_75t_SL g954 ( .A(n_724), .Y(n_954) );
OAI21x1_ASAP7_75t_L g955 ( .A1(n_729), .A2(n_253), .B(n_252), .Y(n_955) );
INVxp67_ASAP7_75t_L g956 ( .A(n_808), .Y(n_956) );
O2A1O1Ixp33_ASAP7_75t_L g957 ( .A1(n_878), .A2(n_702), .B(n_728), .C(n_52), .Y(n_957) );
NOR2x1_ASAP7_75t_SL g958 ( .A(n_926), .B(n_720), .Y(n_958) );
OAI21x1_ASAP7_75t_L g959 ( .A1(n_846), .A2(n_794), .B(n_789), .Y(n_959) );
OAI211xp5_ASAP7_75t_SL g960 ( .A1(n_839), .A2(n_702), .B(n_50), .C(n_52), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_855), .B(n_745), .Y(n_961) );
AOI222xp33_ASAP7_75t_L g962 ( .A1(n_897), .A2(n_734), .B1(n_745), .B2(n_682), .C1(n_794), .C2(n_56), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_861), .A2(n_734), .B1(n_53), .B2(n_54), .Y(n_963) );
HB1xp67_ASAP7_75t_L g964 ( .A(n_861), .Y(n_964) );
BUFx6f_ASAP7_75t_L g965 ( .A(n_947), .Y(n_965) );
INVx2_ASAP7_75t_L g966 ( .A(n_877), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_824), .Y(n_967) );
BUFx8_ASAP7_75t_L g968 ( .A(n_840), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_809), .Y(n_969) );
A2O1A1Ixp33_ASAP7_75t_L g970 ( .A1(n_855), .A2(n_49), .B(n_53), .C(n_54), .Y(n_970) );
BUFx4f_ASAP7_75t_SL g971 ( .A(n_836), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_918), .B(n_55), .Y(n_972) );
OAI221xp5_ASAP7_75t_L g973 ( .A1(n_839), .A2(n_55), .B1(n_56), .B2(n_58), .C(n_59), .Y(n_973) );
AOI221xp5_ASAP7_75t_L g974 ( .A1(n_889), .A2(n_58), .B1(n_60), .B2(n_61), .C(n_62), .Y(n_974) );
AOI21xp5_ASAP7_75t_L g975 ( .A1(n_821), .A2(n_249), .B(n_248), .Y(n_975) );
INVx3_ASAP7_75t_L g976 ( .A(n_947), .Y(n_976) );
INVx2_ASAP7_75t_L g977 ( .A(n_877), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_811), .Y(n_978) );
NAND3xp33_ASAP7_75t_L g979 ( .A(n_919), .B(n_60), .C(n_61), .Y(n_979) );
AO21x2_ASAP7_75t_L g980 ( .A1(n_813), .A2(n_240), .B(n_237), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_861), .A2(n_62), .B1(n_63), .B2(n_64), .Y(n_981) );
OAI22xp5_ASAP7_75t_L g982 ( .A1(n_905), .A2(n_63), .B1(n_64), .B2(n_65), .Y(n_982) );
BUFx4f_ASAP7_75t_SL g983 ( .A(n_836), .Y(n_983) );
OAI221xp5_ASAP7_75t_SL g984 ( .A1(n_828), .A2(n_65), .B1(n_66), .B2(n_69), .C(n_70), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_899), .A2(n_69), .B1(n_71), .B2(n_72), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_818), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_930), .B(n_71), .Y(n_987) );
INVx2_ASAP7_75t_SL g988 ( .A(n_825), .Y(n_988) );
OAI211xp5_ASAP7_75t_L g989 ( .A1(n_816), .A2(n_73), .B(n_74), .C(n_75), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_843), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_899), .A2(n_893), .B1(n_852), .B2(n_946), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_852), .A2(n_75), .B1(n_76), .B2(n_77), .Y(n_992) );
BUFx3_ASAP7_75t_L g993 ( .A(n_871), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_862), .Y(n_994) );
OR2x6_ASAP7_75t_L g995 ( .A(n_926), .B(n_77), .Y(n_995) );
NOR2x1_ASAP7_75t_L g996 ( .A(n_895), .B(n_78), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_930), .B(n_79), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_852), .A2(n_80), .B1(n_81), .B2(n_82), .Y(n_998) );
AO31x2_ASAP7_75t_L g999 ( .A1(n_919), .A2(n_81), .A3(n_83), .B(n_84), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_893), .A2(n_85), .B1(n_86), .B2(n_87), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_893), .A2(n_216), .B1(n_217), .B2(n_219), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_885), .A2(n_220), .B1(n_224), .B2(n_227), .Y(n_1002) );
AOI211xp5_ASAP7_75t_L g1003 ( .A1(n_951), .A2(n_228), .B(n_229), .C(n_230), .Y(n_1003) );
AOI221xp5_ASAP7_75t_L g1004 ( .A1(n_889), .A2(n_231), .B1(n_869), .B2(n_820), .C(n_945), .Y(n_1004) );
OR2x6_ASAP7_75t_L g1005 ( .A(n_926), .B(n_854), .Y(n_1005) );
AOI21xp33_ASAP7_75t_L g1006 ( .A1(n_810), .A2(n_929), .B(n_900), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_885), .A2(n_943), .B1(n_820), .B2(n_870), .Y(n_1007) );
AO221x2_ASAP7_75t_L g1008 ( .A1(n_951), .A2(n_841), .B1(n_826), .B2(n_949), .C(n_938), .Y(n_1008) );
OAI22xp5_ASAP7_75t_L g1009 ( .A1(n_905), .A2(n_817), .B1(n_810), .B2(n_806), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_885), .A2(n_806), .B1(n_954), .B2(n_952), .Y(n_1010) );
BUFx12f_ASAP7_75t_L g1011 ( .A(n_924), .Y(n_1011) );
AOI222xp33_ASAP7_75t_L g1012 ( .A1(n_923), .A2(n_812), .B1(n_844), .B2(n_924), .C1(n_849), .C2(n_909), .Y(n_1012) );
OAI22xp5_ASAP7_75t_L g1013 ( .A1(n_817), .A2(n_910), .B1(n_911), .B2(n_829), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_886), .Y(n_1014) );
AO221x2_ASAP7_75t_L g1015 ( .A1(n_841), .A2(n_922), .B1(n_939), .B2(n_864), .C(n_940), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_914), .B(n_868), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_937), .B(n_825), .Y(n_1017) );
OA21x2_ASAP7_75t_L g1018 ( .A1(n_807), .A2(n_848), .B(n_847), .Y(n_1018) );
NAND3xp33_ASAP7_75t_L g1019 ( .A(n_917), .B(n_883), .C(n_835), .Y(n_1019) );
OAI22xp33_ASAP7_75t_L g1020 ( .A1(n_831), .A2(n_834), .B1(n_851), .B2(n_895), .Y(n_1020) );
OAI221xp5_ASAP7_75t_L g1021 ( .A1(n_917), .A2(n_887), .B1(n_830), .B2(n_814), .C(n_906), .Y(n_1021) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_906), .A2(n_831), .B1(n_845), .B2(n_833), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_932), .A2(n_942), .B1(n_936), .B2(n_871), .Y(n_1023) );
AOI221xp5_ASAP7_75t_L g1024 ( .A1(n_867), .A2(n_835), .B1(n_876), .B2(n_850), .C(n_881), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_921), .A2(n_801), .B1(n_909), .B2(n_890), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_921), .A2(n_845), .B1(n_860), .B2(n_838), .Y(n_1026) );
INVx2_ASAP7_75t_L g1027 ( .A(n_805), .Y(n_1027) );
AO21x2_ASAP7_75t_L g1028 ( .A1(n_863), .A2(n_804), .B(n_822), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_833), .A2(n_860), .B1(n_838), .B2(n_891), .Y(n_1029) );
AOI222xp33_ASAP7_75t_L g1030 ( .A1(n_948), .A2(n_898), .B1(n_858), .B2(n_865), .C1(n_880), .C2(n_853), .Y(n_1030) );
BUFx2_ASAP7_75t_L g1031 ( .A(n_908), .Y(n_1031) );
A2O1A1Ixp33_ASAP7_75t_L g1032 ( .A1(n_907), .A2(n_916), .B(n_858), .C(n_884), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_853), .A2(n_866), .B1(n_908), .B2(n_803), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_842), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_805), .B(n_815), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g1036 ( .A(n_815), .B(n_803), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_935), .B(n_913), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_935), .B(n_913), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_842), .B(n_819), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_842), .Y(n_1040) );
OAI21xp5_ASAP7_75t_L g1041 ( .A1(n_907), .A2(n_916), .B(n_802), .Y(n_1041) );
AO21x2_ASAP7_75t_L g1042 ( .A1(n_863), .A2(n_822), .B(n_837), .Y(n_1042) );
INVx4_ASAP7_75t_L g1043 ( .A(n_896), .Y(n_1043) );
AND2x4_ASAP7_75t_L g1044 ( .A(n_896), .B(n_904), .Y(n_1044) );
INVx3_ASAP7_75t_L g1045 ( .A(n_866), .Y(n_1045) );
AND2x4_ASAP7_75t_L g1046 ( .A(n_904), .B(n_955), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_866), .A2(n_802), .B1(n_901), .B2(n_934), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_866), .A2(n_802), .B1(n_901), .B2(n_934), .Y(n_1048) );
A2O1A1Ixp33_ASAP7_75t_L g1049 ( .A1(n_884), .A2(n_894), .B(n_955), .C(n_827), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_866), .A2(n_901), .B1(n_933), .B2(n_882), .Y(n_1050) );
BUFx6f_ASAP7_75t_L g1051 ( .A(n_859), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_842), .Y(n_1052) );
INVx2_ASAP7_75t_L g1053 ( .A(n_819), .Y(n_1053) );
AOI22xp33_ASAP7_75t_SL g1054 ( .A1(n_866), .A2(n_882), .B1(n_875), .B2(n_873), .Y(n_1054) );
NAND2xp5_ASAP7_75t_SL g1055 ( .A(n_928), .B(n_856), .Y(n_1055) );
BUFx12f_ASAP7_75t_L g1056 ( .A(n_819), .Y(n_1056) );
AO21x2_ASAP7_75t_L g1057 ( .A1(n_823), .A2(n_925), .B(n_902), .Y(n_1057) );
OAI22xp5_ASAP7_75t_L g1058 ( .A1(n_879), .A2(n_872), .B1(n_874), .B2(n_953), .Y(n_1058) );
AOI22xp5_ASAP7_75t_L g1059 ( .A1(n_912), .A2(n_944), .B1(n_950), .B2(n_920), .Y(n_1059) );
AOI221xp5_ASAP7_75t_L g1060 ( .A1(n_832), .A2(n_927), .B1(n_931), .B2(n_941), .C(n_888), .Y(n_1060) );
A2O1A1Ixp33_ASAP7_75t_L g1061 ( .A1(n_892), .A2(n_855), .B(n_753), .C(n_730), .Y(n_1061) );
AOI221xp5_ASAP7_75t_L g1062 ( .A1(n_915), .A2(n_855), .B1(n_665), .B2(n_878), .C(n_610), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_903), .B(n_855), .Y(n_1063) );
OAI22xp5_ASAP7_75t_L g1064 ( .A1(n_878), .A2(n_669), .B1(n_685), .B2(n_621), .Y(n_1064) );
OAI211xp5_ASAP7_75t_L g1065 ( .A1(n_816), .A2(n_592), .B(n_669), .C(n_579), .Y(n_1065) );
OAI21xp33_ASAP7_75t_L g1066 ( .A1(n_878), .A2(n_662), .B(n_855), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_861), .A2(n_742), .B1(n_855), .B2(n_727), .Y(n_1067) );
BUFx12f_ASAP7_75t_L g1068 ( .A(n_840), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_861), .A2(n_742), .B1(n_855), .B2(n_727), .Y(n_1069) );
OAI22xp33_ASAP7_75t_L g1070 ( .A1(n_857), .A2(n_669), .B1(n_662), .B2(n_681), .Y(n_1070) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_855), .B(n_878), .Y(n_1071) );
CKINVDCx5p33_ASAP7_75t_R g1072 ( .A(n_836), .Y(n_1072) );
BUFx6f_ASAP7_75t_L g1073 ( .A(n_947), .Y(n_1073) );
OAI221xp5_ASAP7_75t_L g1074 ( .A1(n_855), .A2(n_878), .B1(n_839), .B2(n_592), .C(n_740), .Y(n_1074) );
AOI21xp33_ASAP7_75t_L g1075 ( .A1(n_878), .A2(n_855), .B(n_763), .Y(n_1075) );
AOI22xp33_ASAP7_75t_SL g1076 ( .A1(n_857), .A2(n_662), .B1(n_701), .B2(n_672), .Y(n_1076) );
OR2x6_ASAP7_75t_L g1077 ( .A(n_808), .B(n_926), .Y(n_1077) );
OA21x2_ASAP7_75t_L g1078 ( .A1(n_846), .A2(n_670), .B(n_807), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_861), .A2(n_742), .B1(n_855), .B2(n_727), .Y(n_1079) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_855), .B(n_878), .Y(n_1080) );
AOI222xp33_ASAP7_75t_L g1081 ( .A1(n_897), .A2(n_755), .B1(n_758), .B2(n_742), .C1(n_855), .C2(n_701), .Y(n_1081) );
BUFx2_ASAP7_75t_L g1082 ( .A(n_808), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_824), .Y(n_1083) );
OAI22xp5_ASAP7_75t_L g1084 ( .A1(n_878), .A2(n_669), .B1(n_685), .B2(n_621), .Y(n_1084) );
AND2x4_ASAP7_75t_L g1085 ( .A(n_825), .B(n_834), .Y(n_1085) );
INVx3_ASAP7_75t_L g1086 ( .A(n_947), .Y(n_1086) );
INVxp67_ASAP7_75t_L g1087 ( .A(n_808), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1016), .Y(n_1088) );
AND2x2_ASAP7_75t_SL g1089 ( .A(n_1050), .B(n_964), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_1008), .A2(n_1075), .B1(n_1074), .B2(n_995), .Y(n_1090) );
AND2x4_ASAP7_75t_L g1091 ( .A(n_966), .B(n_977), .Y(n_1091) );
INVx2_ASAP7_75t_L g1092 ( .A(n_1035), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1027), .B(n_1039), .Y(n_1093) );
AND2x4_ASAP7_75t_L g1094 ( .A(n_958), .B(n_1043), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1014), .B(n_967), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1034), .Y(n_1096) );
INVx2_ASAP7_75t_L g1097 ( .A(n_1078), .Y(n_1097) );
BUFx2_ASAP7_75t_L g1098 ( .A(n_995), .Y(n_1098) );
INVx4_ASAP7_75t_R g1099 ( .A(n_993), .Y(n_1099) );
AOI22xp5_ASAP7_75t_L g1100 ( .A1(n_1064), .A2(n_1084), .B1(n_1076), .B2(n_1070), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1040), .Y(n_1101) );
INVx4_ASAP7_75t_SL g1102 ( .A(n_995), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1052), .Y(n_1103) );
INVx3_ASAP7_75t_L g1104 ( .A(n_1043), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1083), .B(n_969), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1053), .Y(n_1106) );
HB1xp67_ASAP7_75t_L g1107 ( .A(n_1082), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_986), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1036), .Y(n_1109) );
HB1xp67_ASAP7_75t_L g1110 ( .A(n_1031), .Y(n_1110) );
AND2x4_ASAP7_75t_L g1111 ( .A(n_1044), .B(n_1045), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_978), .B(n_990), .Y(n_1112) );
INVx2_ASAP7_75t_L g1113 ( .A(n_959), .Y(n_1113) );
AND2x4_ASAP7_75t_L g1114 ( .A(n_1044), .B(n_1045), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1115 ( .A(n_1071), .B(n_1080), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_994), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_991), .B(n_1007), .Y(n_1117) );
NAND2x1_ASAP7_75t_L g1118 ( .A(n_1046), .B(n_1018), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_999), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_999), .Y(n_1120) );
INVx2_ASAP7_75t_SL g1121 ( .A(n_1085), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_999), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1056), .Y(n_1123) );
NOR2x1_ASAP7_75t_L g1124 ( .A(n_1020), .B(n_1077), .Y(n_1124) );
INVxp67_ASAP7_75t_SL g1125 ( .A(n_961), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_976), .B(n_1086), .Y(n_1126) );
HB1xp67_ASAP7_75t_L g1127 ( .A(n_1085), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_976), .B(n_1086), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_965), .B(n_1073), .Y(n_1129) );
INVx2_ASAP7_75t_L g1130 ( .A(n_1018), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_965), .B(n_1073), .Y(n_1131) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1063), .Y(n_1132) );
CKINVDCx20_ASAP7_75t_R g1133 ( .A(n_971), .Y(n_1133) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_1008), .A2(n_962), .B1(n_1066), .B2(n_1005), .Y(n_1134) );
INVx3_ASAP7_75t_L g1135 ( .A(n_988), .Y(n_1135) );
HB1xp67_ASAP7_75t_L g1136 ( .A(n_1077), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1003), .B(n_1005), .Y(n_1137) );
HB1xp67_ASAP7_75t_L g1138 ( .A(n_1077), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g1139 ( .A1(n_1066), .A2(n_1005), .B1(n_1081), .B2(n_1062), .Y(n_1139) );
AND2x4_ASAP7_75t_L g1140 ( .A(n_1037), .B(n_1038), .Y(n_1140) );
HB1xp67_ASAP7_75t_L g1141 ( .A(n_956), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1003), .B(n_992), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_998), .B(n_1000), .Y(n_1143) );
HB1xp67_ASAP7_75t_L g1144 ( .A(n_1087), .Y(n_1144) );
CKINVDCx16_ASAP7_75t_R g1145 ( .A(n_1068), .Y(n_1145) );
BUFx3_ASAP7_75t_L g1146 ( .A(n_968), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_1010), .B(n_1079), .Y(n_1147) );
OR2x2_ASAP7_75t_L g1148 ( .A(n_1017), .B(n_1013), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1024), .B(n_981), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1006), .B(n_970), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1022), .Y(n_1151) );
INVxp67_ASAP7_75t_L g1152 ( .A(n_968), .Y(n_1152) );
INVx8_ASAP7_75t_L g1153 ( .A(n_987), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_997), .B(n_1030), .Y(n_1154) );
INVx5_ASAP7_75t_L g1155 ( .A(n_1051), .Y(n_1155) );
NOR2xp33_ASAP7_75t_L g1156 ( .A(n_1065), .B(n_1069), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1061), .B(n_1023), .Y(n_1157) );
NOR2xp33_ASAP7_75t_L g1158 ( .A(n_1067), .B(n_972), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1026), .B(n_963), .Y(n_1159) );
BUFx2_ASAP7_75t_L g1160 ( .A(n_1046), .Y(n_1160) );
INVx2_ASAP7_75t_SL g1161 ( .A(n_983), .Y(n_1161) );
BUFx3_ASAP7_75t_L g1162 ( .A(n_1072), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_974), .B(n_979), .Y(n_1163) );
NOR2xp33_ASAP7_75t_L g1164 ( .A(n_1021), .B(n_996), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_973), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_982), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_989), .Y(n_1167) );
NAND2x1p5_ASAP7_75t_L g1168 ( .A(n_1051), .B(n_1059), .Y(n_1168) );
AND2x4_ASAP7_75t_L g1169 ( .A(n_1033), .B(n_980), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1029), .B(n_1012), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1171 ( .A(n_1004), .B(n_1025), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_979), .B(n_985), .Y(n_1172) );
HB1xp67_ASAP7_75t_L g1173 ( .A(n_1009), .Y(n_1173) );
INVx1_ASAP7_75t_L g1174 ( .A(n_960), .Y(n_1174) );
INVx2_ASAP7_75t_L g1175 ( .A(n_1057), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1047), .B(n_1048), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1041), .B(n_1019), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1019), .B(n_1002), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1001), .B(n_1015), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1015), .B(n_1042), .Y(n_1180) );
CKINVDCx5p33_ASAP7_75t_R g1181 ( .A(n_1011), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1059), .Y(n_1182) );
INVx2_ASAP7_75t_L g1183 ( .A(n_1057), .Y(n_1183) );
INVx2_ASAP7_75t_L g1184 ( .A(n_1028), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1054), .B(n_1028), .Y(n_1185) );
BUFx6f_ASAP7_75t_L g1186 ( .A(n_1055), .Y(n_1186) );
HB1xp67_ASAP7_75t_L g1187 ( .A(n_984), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1032), .B(n_957), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1058), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1049), .B(n_975), .Y(n_1190) );
BUFx3_ASAP7_75t_L g1191 ( .A(n_1094), .Y(n_1191) );
OAI22xp5_ASAP7_75t_L g1192 ( .A1(n_1090), .A2(n_1060), .B1(n_1098), .B2(n_1134), .Y(n_1192) );
AOI22xp5_ASAP7_75t_L g1193 ( .A1(n_1149), .A2(n_1164), .B1(n_1154), .B2(n_1156), .Y(n_1193) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1095), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1105), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_1088), .B(n_1112), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1117), .B(n_1112), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1108), .Y(n_1198) );
NOR2xp33_ASAP7_75t_R g1199 ( .A(n_1133), .B(n_1145), .Y(n_1199) );
NOR2xp33_ASAP7_75t_L g1200 ( .A(n_1115), .B(n_1187), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1116), .Y(n_1201) );
AOI33xp33_ASAP7_75t_L g1202 ( .A1(n_1139), .A2(n_1116), .A3(n_1157), .B1(n_1149), .B2(n_1154), .B3(n_1137), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1140), .B(n_1110), .Y(n_1203) );
NOR3xp33_ASAP7_75t_L g1204 ( .A(n_1158), .B(n_1147), .C(n_1170), .Y(n_1204) );
OAI21xp5_ASAP7_75t_L g1205 ( .A1(n_1171), .A2(n_1167), .B(n_1174), .Y(n_1205) );
INVxp67_ASAP7_75t_SL g1206 ( .A(n_1092), .Y(n_1206) );
INVx1_ASAP7_75t_SL g1207 ( .A(n_1133), .Y(n_1207) );
INVx4_ASAP7_75t_L g1208 ( .A(n_1102), .Y(n_1208) );
NAND2xp5_ASAP7_75t_L g1209 ( .A(n_1140), .B(n_1098), .Y(n_1209) );
AOI322xp5_ASAP7_75t_L g1210 ( .A1(n_1124), .A2(n_1137), .A3(n_1100), .B1(n_1152), .B2(n_1146), .C1(n_1142), .C2(n_1161), .Y(n_1210) );
OR2x2_ASAP7_75t_L g1211 ( .A(n_1107), .B(n_1127), .Y(n_1211) );
INVx4_ASAP7_75t_L g1212 ( .A(n_1102), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1121), .B(n_1102), .Y(n_1213) );
AOI22xp33_ASAP7_75t_L g1214 ( .A1(n_1142), .A2(n_1166), .B1(n_1163), .B2(n_1143), .Y(n_1214) );
OAI21xp33_ASAP7_75t_L g1215 ( .A1(n_1150), .A2(n_1180), .B(n_1179), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1096), .Y(n_1216) );
NOR2xp33_ASAP7_75t_L g1217 ( .A(n_1159), .B(n_1141), .Y(n_1217) );
INVxp67_ASAP7_75t_SL g1218 ( .A(n_1092), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1096), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1101), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1101), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1144), .B(n_1159), .Y(n_1222) );
NAND2xp5_ASAP7_75t_SL g1223 ( .A(n_1104), .B(n_1094), .Y(n_1223) );
AO21x2_ASAP7_75t_L g1224 ( .A1(n_1184), .A2(n_1183), .B(n_1175), .Y(n_1224) );
OR2x2_ASAP7_75t_L g1225 ( .A(n_1093), .B(n_1125), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1177), .B(n_1180), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1103), .B(n_1176), .Y(n_1227) );
INVx2_ASAP7_75t_L g1228 ( .A(n_1097), .Y(n_1228) );
BUFx3_ASAP7_75t_L g1229 ( .A(n_1094), .Y(n_1229) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1130), .Y(n_1230) );
OAI221xp5_ASAP7_75t_L g1231 ( .A1(n_1165), .A2(n_1150), .B1(n_1138), .B2(n_1136), .C(n_1163), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1135), .B(n_1131), .Y(n_1232) );
AOI22xp33_ASAP7_75t_L g1233 ( .A1(n_1143), .A2(n_1172), .B1(n_1179), .B2(n_1178), .Y(n_1233) );
OR2x2_ASAP7_75t_L g1234 ( .A(n_1148), .B(n_1153), .Y(n_1234) );
INVx2_ASAP7_75t_SL g1235 ( .A(n_1104), .Y(n_1235) );
OAI22xp5_ASAP7_75t_L g1236 ( .A1(n_1153), .A2(n_1148), .B1(n_1104), .B2(n_1172), .Y(n_1236) );
HB1xp67_ASAP7_75t_L g1237 ( .A(n_1109), .Y(n_1237) );
NOR2xp33_ASAP7_75t_R g1238 ( .A(n_1146), .B(n_1153), .Y(n_1238) );
OAI21xp5_ASAP7_75t_L g1239 ( .A1(n_1188), .A2(n_1132), .B(n_1151), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1091), .Y(n_1240) );
AND2x2_ASAP7_75t_L g1241 ( .A(n_1176), .B(n_1091), .Y(n_1241) );
OR2x2_ASAP7_75t_L g1242 ( .A(n_1129), .B(n_1131), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1119), .B(n_1122), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_1151), .A2(n_1188), .B1(n_1173), .B2(n_1089), .Y(n_1244) );
OAI31xp33_ASAP7_75t_SL g1245 ( .A1(n_1126), .A2(n_1128), .A3(n_1123), .B(n_1111), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1119), .B(n_1122), .Y(n_1246) );
NOR2xp33_ASAP7_75t_L g1247 ( .A(n_1162), .B(n_1089), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1126), .B(n_1128), .Y(n_1248) );
OR2x6_ASAP7_75t_L g1249 ( .A(n_1160), .B(n_1111), .Y(n_1249) );
BUFx6f_ASAP7_75t_L g1250 ( .A(n_1155), .Y(n_1250) );
INVx5_ASAP7_75t_L g1251 ( .A(n_1250), .Y(n_1251) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1216), .Y(n_1252) );
INVx2_ASAP7_75t_SL g1253 ( .A(n_1191), .Y(n_1253) );
HB1xp67_ASAP7_75t_L g1254 ( .A(n_1237), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1226), .B(n_1120), .Y(n_1255) );
INVx2_ASAP7_75t_L g1256 ( .A(n_1230), .Y(n_1256) );
NOR2xp33_ASAP7_75t_L g1257 ( .A(n_1207), .B(n_1181), .Y(n_1257) );
NAND4xp25_ASAP7_75t_L g1258 ( .A(n_1204), .B(n_1185), .C(n_1169), .D(n_1182), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1219), .Y(n_1259) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1220), .Y(n_1260) );
HB1xp67_ASAP7_75t_L g1261 ( .A(n_1237), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1227), .B(n_1106), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1241), .B(n_1106), .Y(n_1263) );
AND2x4_ASAP7_75t_L g1264 ( .A(n_1208), .B(n_1155), .Y(n_1264) );
INVxp67_ASAP7_75t_SL g1265 ( .A(n_1206), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1233), .B(n_1132), .Y(n_1266) );
AND2x4_ASAP7_75t_L g1267 ( .A(n_1208), .B(n_1155), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1197), .B(n_1189), .Y(n_1268) );
BUFx3_ASAP7_75t_L g1269 ( .A(n_1191), .Y(n_1269) );
NAND2xp5_ASAP7_75t_L g1270 ( .A(n_1233), .B(n_1169), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1214), .B(n_1169), .Y(n_1271) );
NAND2x1p5_ASAP7_75t_L g1272 ( .A(n_1212), .B(n_1155), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_1214), .B(n_1190), .Y(n_1273) );
OR2x2_ASAP7_75t_L g1274 ( .A(n_1222), .B(n_1118), .Y(n_1274) );
NAND5xp2_ASAP7_75t_L g1275 ( .A(n_1210), .B(n_1099), .C(n_1190), .D(n_1168), .E(n_1181), .Y(n_1275) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1221), .Y(n_1276) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1243), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1246), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1239), .B(n_1114), .Y(n_1279) );
AND2x4_ASAP7_75t_L g1280 ( .A(n_1212), .B(n_1114), .Y(n_1280) );
AND2x4_ASAP7_75t_SL g1281 ( .A(n_1212), .B(n_1114), .Y(n_1281) );
INVxp67_ASAP7_75t_L g1282 ( .A(n_1218), .Y(n_1282) );
NOR2x1p5_ASAP7_75t_L g1283 ( .A(n_1229), .B(n_1113), .Y(n_1283) );
INVx4_ASAP7_75t_L g1284 ( .A(n_1229), .Y(n_1284) );
NOR3xp33_ASAP7_75t_SL g1285 ( .A(n_1192), .B(n_1168), .C(n_1186), .Y(n_1285) );
BUFx2_ASAP7_75t_L g1286 ( .A(n_1249), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1248), .B(n_1186), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1201), .B(n_1215), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1194), .B(n_1195), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1217), .B(n_1228), .Y(n_1290) );
INVx2_ASAP7_75t_SL g1291 ( .A(n_1223), .Y(n_1291) );
HB1xp67_ASAP7_75t_SL g1292 ( .A(n_1284), .Y(n_1292) );
NAND2xp33_ASAP7_75t_SL g1293 ( .A(n_1284), .B(n_1238), .Y(n_1293) );
INVxp33_ASAP7_75t_L g1294 ( .A(n_1257), .Y(n_1294) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1252), .Y(n_1295) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1252), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_1268), .B(n_1217), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1259), .Y(n_1298) );
OR2x2_ASAP7_75t_L g1299 ( .A(n_1290), .B(n_1225), .Y(n_1299) );
NOR2x1p5_ASAP7_75t_L g1300 ( .A(n_1284), .B(n_1258), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1255), .B(n_1203), .Y(n_1301) );
INVx2_ASAP7_75t_L g1302 ( .A(n_1256), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1303 ( .A(n_1268), .B(n_1193), .Y(n_1303) );
NOR2xp67_ASAP7_75t_L g1304 ( .A(n_1284), .B(n_1235), .Y(n_1304) );
OR2x2_ASAP7_75t_L g1305 ( .A(n_1290), .B(n_1209), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1263), .B(n_1240), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1259), .Y(n_1307) );
OR2x2_ASAP7_75t_L g1308 ( .A(n_1277), .B(n_1196), .Y(n_1308) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1260), .Y(n_1309) );
NAND2x1p5_ASAP7_75t_L g1310 ( .A(n_1283), .B(n_1223), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1277), .B(n_1224), .Y(n_1311) );
OR2x2_ASAP7_75t_L g1312 ( .A(n_1278), .B(n_1242), .Y(n_1312) );
NOR2x1_ASAP7_75t_L g1313 ( .A(n_1283), .B(n_1211), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1287), .B(n_1249), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1315 ( .A(n_1289), .B(n_1202), .Y(n_1315) );
NAND2xp33_ASAP7_75t_SL g1316 ( .A(n_1285), .B(n_1238), .Y(n_1316) );
INVx1_ASAP7_75t_SL g1317 ( .A(n_1269), .Y(n_1317) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1276), .Y(n_1318) );
OR2x2_ASAP7_75t_L g1319 ( .A(n_1299), .B(n_1282), .Y(n_1319) );
OAI21xp5_ASAP7_75t_L g1320 ( .A1(n_1313), .A2(n_1258), .B(n_1200), .Y(n_1320) );
INVxp67_ASAP7_75t_L g1321 ( .A(n_1292), .Y(n_1321) );
NAND2xp5_ASAP7_75t_L g1322 ( .A(n_1315), .B(n_1273), .Y(n_1322) );
NOR2xp33_ASAP7_75t_L g1323 ( .A(n_1294), .B(n_1247), .Y(n_1323) );
OAI21xp5_ASAP7_75t_L g1324 ( .A1(n_1313), .A2(n_1205), .B(n_1265), .Y(n_1324) );
INVx2_ASAP7_75t_L g1325 ( .A(n_1302), .Y(n_1325) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1295), .Y(n_1326) );
AOI22xp5_ASAP7_75t_L g1327 ( .A1(n_1293), .A2(n_1247), .B1(n_1236), .B2(n_1231), .Y(n_1327) );
AOI22xp5_ASAP7_75t_L g1328 ( .A1(n_1300), .A2(n_1273), .B1(n_1244), .B2(n_1266), .Y(n_1328) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1295), .Y(n_1329) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1296), .Y(n_1330) );
AOI22xp5_ASAP7_75t_L g1331 ( .A1(n_1300), .A2(n_1244), .B1(n_1266), .B2(n_1279), .Y(n_1331) );
NAND2xp5_ASAP7_75t_L g1332 ( .A(n_1303), .B(n_1262), .Y(n_1332) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1296), .Y(n_1333) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1298), .Y(n_1334) );
INVx2_ASAP7_75t_L g1335 ( .A(n_1302), .Y(n_1335) );
OAI22xp5_ASAP7_75t_L g1336 ( .A1(n_1304), .A2(n_1234), .B1(n_1253), .B2(n_1286), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1337 ( .A(n_1297), .B(n_1262), .Y(n_1337) );
NAND3xp33_ASAP7_75t_L g1338 ( .A(n_1316), .B(n_1261), .C(n_1254), .Y(n_1338) );
AOI222xp33_ASAP7_75t_L g1339 ( .A1(n_1304), .A2(n_1271), .B1(n_1198), .B2(n_1270), .C1(n_1288), .C2(n_1279), .Y(n_1339) );
O2A1O1Ixp33_ASAP7_75t_L g1340 ( .A1(n_1308), .A2(n_1275), .B(n_1235), .C(n_1288), .Y(n_1340) );
OR2x2_ASAP7_75t_L g1341 ( .A(n_1305), .B(n_1274), .Y(n_1341) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1307), .Y(n_1342) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1309), .Y(n_1343) );
XOR2xp5_ASAP7_75t_L g1344 ( .A(n_1328), .B(n_1308), .Y(n_1344) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1326), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1339), .B(n_1301), .Y(n_1346) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1329), .Y(n_1347) );
NOR2xp33_ASAP7_75t_SL g1348 ( .A(n_1321), .B(n_1317), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_1322), .B(n_1311), .Y(n_1349) );
INVxp33_ASAP7_75t_L g1350 ( .A(n_1323), .Y(n_1350) );
INVx2_ASAP7_75t_L g1351 ( .A(n_1325), .Y(n_1351) );
INVx2_ASAP7_75t_L g1352 ( .A(n_1335), .Y(n_1352) );
OAI21xp5_ASAP7_75t_L g1353 ( .A1(n_1320), .A2(n_1310), .B(n_1253), .Y(n_1353) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1330), .Y(n_1354) );
XOR2x2_ASAP7_75t_L g1355 ( .A(n_1320), .B(n_1199), .Y(n_1355) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1333), .Y(n_1356) );
NOR2x1p5_ASAP7_75t_L g1357 ( .A(n_1338), .B(n_1269), .Y(n_1357) );
INVx2_ASAP7_75t_L g1358 ( .A(n_1334), .Y(n_1358) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1343), .Y(n_1359) );
OR2x2_ASAP7_75t_L g1360 ( .A(n_1319), .B(n_1312), .Y(n_1360) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1342), .Y(n_1361) );
NOR2xp67_ASAP7_75t_SL g1362 ( .A(n_1324), .B(n_1251), .Y(n_1362) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1345), .Y(n_1363) );
OAI222xp33_ASAP7_75t_L g1364 ( .A1(n_1362), .A2(n_1331), .B1(n_1327), .B2(n_1340), .C1(n_1336), .C2(n_1341), .Y(n_1364) );
INVx3_ASAP7_75t_L g1365 ( .A(n_1355), .Y(n_1365) );
NOR2xp33_ASAP7_75t_L g1366 ( .A(n_1350), .B(n_1332), .Y(n_1366) );
CKINVDCx5p33_ASAP7_75t_R g1367 ( .A(n_1355), .Y(n_1367) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1345), .Y(n_1368) );
NOR2x1_ASAP7_75t_L g1369 ( .A(n_1357), .B(n_1275), .Y(n_1369) );
AOI22xp5_ASAP7_75t_L g1370 ( .A1(n_1346), .A2(n_1314), .B1(n_1270), .B2(n_1337), .Y(n_1370) );
AOI21xp33_ASAP7_75t_SL g1371 ( .A1(n_1353), .A2(n_1245), .B(n_1310), .Y(n_1371) );
AOI22xp5_ASAP7_75t_L g1372 ( .A1(n_1346), .A2(n_1314), .B1(n_1271), .B2(n_1306), .Y(n_1372) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1347), .Y(n_1373) );
AOI21xp5_ASAP7_75t_L g1374 ( .A1(n_1348), .A2(n_1310), .B(n_1281), .Y(n_1374) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1347), .Y(n_1375) );
XNOR2xp5_ASAP7_75t_L g1376 ( .A(n_1367), .B(n_1344), .Y(n_1376) );
OAI211xp5_ASAP7_75t_SL g1377 ( .A1(n_1365), .A2(n_1360), .B(n_1349), .C(n_1361), .Y(n_1377) );
OAI21xp5_ASAP7_75t_L g1378 ( .A1(n_1364), .A2(n_1362), .B(n_1344), .Y(n_1378) );
XNOR2x1_ASAP7_75t_L g1379 ( .A(n_1365), .B(n_1360), .Y(n_1379) );
AOI221xp5_ASAP7_75t_L g1380 ( .A1(n_1371), .A2(n_1361), .B1(n_1359), .B2(n_1354), .C(n_1356), .Y(n_1380) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1363), .Y(n_1381) );
INVx1_ASAP7_75t_SL g1382 ( .A(n_1374), .Y(n_1382) );
OAI22xp33_ASAP7_75t_L g1383 ( .A1(n_1369), .A2(n_1312), .B1(n_1291), .B2(n_1251), .Y(n_1383) );
AND2x4_ASAP7_75t_L g1384 ( .A(n_1382), .B(n_1366), .Y(n_1384) );
OR2x2_ASAP7_75t_L g1385 ( .A(n_1379), .B(n_1368), .Y(n_1385) );
OR2x2_ASAP7_75t_L g1386 ( .A(n_1381), .B(n_1373), .Y(n_1386) );
NOR3xp33_ASAP7_75t_L g1387 ( .A(n_1378), .B(n_1370), .C(n_1375), .Y(n_1387) );
CKINVDCx5p33_ASAP7_75t_R g1388 ( .A(n_1376), .Y(n_1388) );
NOR2xp33_ASAP7_75t_L g1389 ( .A(n_1377), .B(n_1372), .Y(n_1389) );
NAND2xp5_ASAP7_75t_L g1390 ( .A(n_1380), .B(n_1358), .Y(n_1390) );
NOR2xp67_ASAP7_75t_L g1391 ( .A(n_1384), .B(n_1383), .Y(n_1391) );
OAI22xp33_ASAP7_75t_L g1392 ( .A1(n_1385), .A2(n_1251), .B1(n_1272), .B2(n_1358), .Y(n_1392) );
INVx2_ASAP7_75t_L g1393 ( .A(n_1386), .Y(n_1393) );
OR2x2_ASAP7_75t_L g1394 ( .A(n_1390), .B(n_1352), .Y(n_1394) );
XNOR2xp5_ASAP7_75t_L g1395 ( .A(n_1388), .B(n_1232), .Y(n_1395) );
INVx2_ASAP7_75t_L g1396 ( .A(n_1393), .Y(n_1396) );
OA21x2_ASAP7_75t_L g1397 ( .A1(n_1391), .A2(n_1387), .B(n_1389), .Y(n_1397) );
INVx2_ASAP7_75t_L g1398 ( .A(n_1394), .Y(n_1398) );
OAI22xp5_ASAP7_75t_SL g1399 ( .A1(n_1397), .A2(n_1395), .B1(n_1392), .B2(n_1251), .Y(n_1399) );
AND3x4_ASAP7_75t_L g1400 ( .A(n_1396), .B(n_1280), .C(n_1267), .Y(n_1400) );
INVx2_ASAP7_75t_L g1401 ( .A(n_1398), .Y(n_1401) );
NOR2xp33_ASAP7_75t_L g1402 ( .A(n_1397), .B(n_1351), .Y(n_1402) );
OAI22x1_ASAP7_75t_L g1403 ( .A1(n_1401), .A2(n_1402), .B1(n_1400), .B2(n_1399), .Y(n_1403) );
AOI22xp5_ASAP7_75t_L g1404 ( .A1(n_1403), .A2(n_1213), .B1(n_1281), .B2(n_1264), .Y(n_1404) );
XNOR2xp5_ASAP7_75t_L g1405 ( .A(n_1404), .B(n_1272), .Y(n_1405) );
AOI21xp5_ASAP7_75t_L g1406 ( .A1(n_1405), .A2(n_1318), .B(n_1309), .Y(n_1406) );
endmodule