module fake_jpeg_26986_n_246 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_246);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_246;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_3),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_34),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_24),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_43),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_36),
.B1(n_41),
.B2(n_39),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_46),
.A2(n_48),
.B1(n_58),
.B2(n_59),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_27),
.B1(n_33),
.B2(n_23),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_64),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_27),
.B1(n_33),
.B2(n_23),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_61),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_62),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_21),
.B1(n_18),
.B2(n_29),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_57),
.B1(n_32),
.B2(n_31),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_21),
.B1(n_18),
.B2(n_29),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_32),
.B1(n_31),
.B2(n_25),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_32),
.B1(n_31),
.B2(n_25),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_43),
.Y(n_77)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_26),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_70),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_50),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_71),
.A2(n_19),
.B1(n_3),
.B2(n_4),
.Y(n_103)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_87),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_79),
.Y(n_93)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_43),
.B1(n_25),
.B2(n_26),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_78),
.A2(n_49),
.B1(n_52),
.B2(n_50),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_16),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_15),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_54),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_22),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_78),
.B(n_84),
.Y(n_104)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_67),
.Y(n_90)
);

INVx5_ASAP7_75t_SL g111 ( 
.A(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_56),
.B(n_1),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_91),
.B(n_1),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_66),
.B1(n_65),
.B2(n_53),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_101),
.B1(n_107),
.B2(n_78),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_66),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_99),
.Y(n_120)
);

AOI32xp33_ASAP7_75t_L g98 ( 
.A1(n_69),
.A2(n_56),
.A3(n_59),
.B1(n_19),
.B2(n_22),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_98),
.A2(n_74),
.B(n_70),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_51),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_102),
.B(n_4),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_78),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_52),
.B1(n_51),
.B2(n_5),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_86),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_73),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_110),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_2),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_113),
.B(n_116),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_89),
.B(n_88),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_2),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_118),
.A2(n_119),
.B1(n_111),
.B2(n_86),
.Y(n_158)
);

AO32x1_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_77),
.A3(n_78),
.B1(n_76),
.B2(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_127),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_76),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_122),
.B(n_126),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_125),
.B(n_133),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_124),
.B(n_102),
.Y(n_141)
);

HAxp5_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_90),
.CON(n_125),
.SN(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_72),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_92),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_131),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_136),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_135),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_112),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_140),
.A2(n_98),
.B(n_93),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_144),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_108),
.C(n_116),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_148),
.C(n_156),
.Y(n_172)
);

INVx5_ASAP7_75t_SL g144 ( 
.A(n_132),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_108),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_157),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_126),
.C(n_133),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_114),
.C(n_106),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_150),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_152),
.A2(n_155),
.B(n_140),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_132),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_153),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_93),
.C(n_114),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_111),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_159),
.Y(n_167)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_136),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_111),
.B1(n_113),
.B2(n_96),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_162),
.A2(n_138),
.B1(n_121),
.B2(n_127),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_142),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_164),
.Y(n_185)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_175),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_168),
.A2(n_177),
.B(n_74),
.Y(n_199)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_155),
.A2(n_130),
.B(n_123),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_168),
.B(n_149),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_129),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_178),
.Y(n_188)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_176),
.A2(n_143),
.B1(n_147),
.B2(n_156),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_123),
.B(n_130),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_140),
.C(n_125),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_181),
.Y(n_193)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_144),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_182),
.B(n_183),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_118),
.C(n_96),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_181),
.A2(n_163),
.B1(n_151),
.B2(n_160),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_184),
.A2(n_189),
.B1(n_190),
.B2(n_198),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_177),
.Y(n_202)
);

NAND2xp33_ASAP7_75t_SL g189 ( 
.A(n_173),
.B(n_152),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_165),
.A2(n_163),
.B1(n_151),
.B2(n_180),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_179),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_194),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_157),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_197),
.Y(n_211)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_167),
.Y(n_201)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_202),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_172),
.C(n_183),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_204),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_172),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_166),
.C(n_170),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_206),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_178),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_SL g207 ( 
.A1(n_199),
.A2(n_170),
.B(n_174),
.C(n_9),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_192),
.B(n_200),
.Y(n_215)
);

BUFx24_ASAP7_75t_SL g209 ( 
.A(n_185),
.Y(n_209)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_192),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_196),
.C(n_190),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_SL g229 ( 
.A1(n_215),
.A2(n_13),
.B(n_217),
.C(n_219),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_207),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_211),
.A2(n_196),
.B1(n_193),
.B2(n_184),
.Y(n_219)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_208),
.A2(n_193),
.B1(n_194),
.B2(n_198),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_222),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_211),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_212),
.C(n_207),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_228),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_222),
.Y(n_232)
);

OAI211xp5_ASAP7_75t_SL g226 ( 
.A1(n_215),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_220),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_10),
.C(n_13),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_229),
.A2(n_221),
.B(n_218),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_230),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_233),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_232),
.B(n_235),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_214),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_234),
.C(n_229),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_218),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_238),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_240),
.A2(n_227),
.B(n_214),
.Y(n_241)
);

BUFx24_ASAP7_75t_SL g244 ( 
.A(n_241),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_237),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_244),
.B(n_243),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_242),
.Y(n_246)
);


endmodule