module fake_netlist_6_1477_n_937 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_937);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_937;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_341;
wire n_362;
wire n_828;
wire n_462;
wire n_607;
wire n_726;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_761;
wire n_428;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_758;
wire n_720;
wire n_525;
wire n_842;
wire n_611;
wire n_491;
wire n_878;
wire n_772;
wire n_656;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_926;
wire n_927;
wire n_839;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_527;
wire n_608;
wire n_261;
wire n_474;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_322;
wire n_707;
wire n_409;
wire n_345;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_404;
wire n_271;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_515;
wire n_434;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_678;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

BUFx2_ASAP7_75t_SL g242 ( 
.A(n_76),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_30),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_196),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_89),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_20),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_74),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_49),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_53),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_52),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_130),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_60),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_159),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_64),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_98),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_13),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_99),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_37),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_213),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_220),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_90),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_181),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_203),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_18),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_170),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_23),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_48),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_28),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_142),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_63),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_125),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_149),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_145),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_4),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_169),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_17),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_68),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_78),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_55),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_5),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_12),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_119),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_36),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_120),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_22),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_154),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_157),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_132),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_228),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_215),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_92),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_66),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_184),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_238),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_208),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_22),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_134),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_50),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_72),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_87),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_231),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_118),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_112),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_172),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_75),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_8),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_201),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_21),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_91),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_47),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_35),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_6),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_24),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_185),
.Y(n_314)
);

BUFx5_ASAP7_75t_L g315 ( 
.A(n_122),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_35),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_237),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_150),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_200),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_34),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_147),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_62),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_121),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_240),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_226),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_174),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_79),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_69),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_160),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_8),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_186),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_211),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_103),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_155),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_239),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_144),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_123),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_81),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_198),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_233),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_146),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_117),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_163),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_56),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_189),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_54),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_227),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_236),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_13),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_32),
.Y(n_350)
);

BUFx2_ASAP7_75t_R g351 ( 
.A(n_175),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_95),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_105),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_58),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_104),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_113),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_214),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_235),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_210),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_100),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_12),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_164),
.Y(n_362)
);

BUFx10_ASAP7_75t_L g363 ( 
.A(n_41),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_93),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_131),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_138),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_219),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_177),
.Y(n_368)
);

BUFx10_ASAP7_75t_L g369 ( 
.A(n_140),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_0),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_110),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_212),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_101),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_199),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_32),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_234),
.Y(n_376)
);

BUFx10_ASAP7_75t_L g377 ( 
.A(n_161),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_88),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_179),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_25),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_82),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_209),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_26),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_83),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_225),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_29),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_39),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_124),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_57),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_16),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_86),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_67),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_71),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_141),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_136),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_139),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_94),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_106),
.Y(n_398)
);

AND2x6_ASAP7_75t_L g399 ( 
.A(n_265),
.B(n_42),
.Y(n_399)
);

INVx5_ASAP7_75t_L g400 ( 
.A(n_244),
.Y(n_400)
);

AND2x6_ASAP7_75t_L g401 ( 
.A(n_265),
.B(n_43),
.Y(n_401)
);

BUFx8_ASAP7_75t_L g402 ( 
.A(n_383),
.Y(n_402)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_244),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_244),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_261),
.B(n_0),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_243),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_282),
.B(n_1),
.Y(n_407)
);

INVx5_ASAP7_75t_L g408 ( 
.A(n_244),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_374),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_376),
.B(n_1),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_261),
.B(n_2),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_376),
.B(n_2),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_3),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_382),
.B(n_3),
.Y(n_414)
);

INVx5_ASAP7_75t_L g415 ( 
.A(n_374),
.Y(n_415)
);

AND2x6_ASAP7_75t_L g416 ( 
.A(n_374),
.B(n_44),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_352),
.B(n_4),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_264),
.B(n_5),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_319),
.B(n_321),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_259),
.B(n_7),
.Y(n_420)
);

INVx5_ASAP7_75t_L g421 ( 
.A(n_374),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_349),
.Y(n_422)
);

BUFx8_ASAP7_75t_L g423 ( 
.A(n_246),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_318),
.B(n_7),
.Y(n_424)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_245),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_315),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_269),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_326),
.B(n_9),
.Y(n_428)
);

INVx5_ASAP7_75t_L g429 ( 
.A(n_363),
.Y(n_429)
);

INVx6_ASAP7_75t_L g430 ( 
.A(n_363),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_292),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_309),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_369),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_309),
.B(n_10),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_369),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_256),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_317),
.B(n_10),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_317),
.B(n_11),
.Y(n_438)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_248),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_315),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_315),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_315),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_280),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_398),
.B(n_14),
.Y(n_444)
);

AND2x6_ASAP7_75t_L g445 ( 
.A(n_241),
.B(n_45),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_266),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_268),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_377),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_315),
.B(n_14),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_315),
.B(n_15),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_280),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_274),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_247),
.B(n_16),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_306),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_375),
.Y(n_455)
);

BUFx12f_ASAP7_75t_L g456 ( 
.A(n_296),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_250),
.B(n_252),
.Y(n_457)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_258),
.B(n_17),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_257),
.B(n_18),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_377),
.B(n_19),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_273),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_279),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_276),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_296),
.Y(n_464)
);

INVx5_ASAP7_75t_L g465 ( 
.A(n_242),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_284),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_281),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_316),
.B(n_20),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_286),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_288),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_394),
.B(n_21),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_283),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_285),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_295),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_308),
.B(n_24),
.Y(n_475)
);

BUFx12f_ASAP7_75t_L g476 ( 
.A(n_311),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_297),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_302),
.B(n_25),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_249),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_307),
.B(n_26),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_310),
.B(n_27),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_251),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_322),
.B(n_28),
.Y(n_483)
);

INVx5_ASAP7_75t_L g484 ( 
.A(n_313),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_328),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_253),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_331),
.B(n_29),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_355),
.B(n_356),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_255),
.Y(n_489)
);

OAI22xp33_ASAP7_75t_L g490 ( 
.A1(n_419),
.A2(n_458),
.B1(n_428),
.B2(n_420),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_406),
.B(n_260),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_452),
.B(n_262),
.Y(n_492)
);

OAI22xp33_ASAP7_75t_L g493 ( 
.A1(n_443),
.A2(n_361),
.B1(n_370),
.B2(n_350),
.Y(n_493)
);

OAI22xp33_ASAP7_75t_L g494 ( 
.A1(n_443),
.A2(n_390),
.B1(n_380),
.B2(n_320),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_424),
.A2(n_272),
.B1(n_275),
.B2(n_254),
.Y(n_495)
);

BUFx10_ASAP7_75t_L g496 ( 
.A(n_430),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_463),
.B(n_263),
.Y(n_497)
);

AND2x4_ASAP7_75t_SL g498 ( 
.A(n_425),
.B(n_294),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_SL g499 ( 
.A(n_460),
.B(n_312),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_467),
.B(n_267),
.Y(n_500)
);

OR2x6_ASAP7_75t_L g501 ( 
.A(n_476),
.B(n_357),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_407),
.A2(n_334),
.B1(n_338),
.B2(n_329),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_472),
.B(n_270),
.Y(n_503)
);

INVx8_ASAP7_75t_L g504 ( 
.A(n_429),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_471),
.A2(n_348),
.B1(n_368),
.B2(n_366),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_425),
.B(n_360),
.Y(n_506)
);

AND2x2_ASAP7_75t_SL g507 ( 
.A(n_412),
.B(n_367),
.Y(n_507)
);

OAI22xp33_ASAP7_75t_SL g508 ( 
.A1(n_430),
.A2(n_372),
.B1(n_373),
.B2(n_371),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_439),
.B(n_378),
.Y(n_509)
);

AND2x2_ASAP7_75t_SL g510 ( 
.A(n_414),
.B(n_385),
.Y(n_510)
);

OAI22xp33_ASAP7_75t_L g511 ( 
.A1(n_451),
.A2(n_386),
.B1(n_387),
.B2(n_330),
.Y(n_511)
);

AO22x2_ASAP7_75t_L g512 ( 
.A1(n_410),
.A2(n_413),
.B1(n_437),
.B2(n_444),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_404),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_479),
.B(n_388),
.Y(n_514)
);

AND2x6_ASAP7_75t_L g515 ( 
.A(n_437),
.B(n_392),
.Y(n_515)
);

AO22x2_ASAP7_75t_L g516 ( 
.A1(n_410),
.A2(n_395),
.B1(n_351),
.B2(n_34),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_473),
.B(n_271),
.Y(n_517)
);

OAI22xp33_ASAP7_75t_L g518 ( 
.A1(n_464),
.A2(n_379),
.B1(n_381),
.B2(n_396),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_429),
.B(n_277),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_422),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_429),
.B(n_278),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_404),
.Y(n_522)
);

BUFx6f_ASAP7_75t_SL g523 ( 
.A(n_433),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_409),
.Y(n_524)
);

AO22x2_ASAP7_75t_L g525 ( 
.A1(n_413),
.A2(n_31),
.B1(n_33),
.B2(n_36),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_427),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_409),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_422),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_427),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_475),
.A2(n_341),
.B1(n_397),
.B2(n_393),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_427),
.Y(n_531)
);

OR2x6_ASAP7_75t_L g532 ( 
.A(n_456),
.B(n_33),
.Y(n_532)
);

OR2x6_ASAP7_75t_L g533 ( 
.A(n_435),
.B(n_448),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_431),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_468),
.A2(n_391),
.B1(n_389),
.B2(n_384),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_489),
.B(n_482),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_486),
.B(n_287),
.Y(n_537)
);

AO22x2_ASAP7_75t_L g538 ( 
.A1(n_444),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_486),
.B(n_289),
.Y(n_539)
);

AO22x2_ASAP7_75t_L g540 ( 
.A1(n_459),
.A2(n_38),
.B1(n_40),
.B2(n_365),
.Y(n_540)
);

OAI22xp33_ASAP7_75t_SL g541 ( 
.A1(n_417),
.A2(n_364),
.B1(n_362),
.B2(n_359),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_431),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_465),
.B(n_290),
.Y(n_543)
);

AOI22x1_ASAP7_75t_L g544 ( 
.A1(n_418),
.A2(n_358),
.B1(n_354),
.B2(n_353),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_399),
.B(n_291),
.Y(n_545)
);

OR2x6_ASAP7_75t_L g546 ( 
.A(n_454),
.B(n_455),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_431),
.Y(n_547)
);

OAI22xp33_ASAP7_75t_R g548 ( 
.A1(n_488),
.A2(n_347),
.B1(n_346),
.B2(n_345),
.Y(n_548)
);

AO22x2_ASAP7_75t_L g549 ( 
.A1(n_459),
.A2(n_344),
.B1(n_343),
.B2(n_342),
.Y(n_549)
);

OAI22xp33_ASAP7_75t_SL g550 ( 
.A1(n_405),
.A2(n_340),
.B1(n_339),
.B2(n_337),
.Y(n_550)
);

OAI22xp33_ASAP7_75t_L g551 ( 
.A1(n_478),
.A2(n_336),
.B1(n_335),
.B2(n_333),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_432),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_480),
.A2(n_303),
.B1(n_327),
.B2(n_325),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_484),
.B(n_293),
.Y(n_554)
);

INVxp33_ASAP7_75t_L g555 ( 
.A(n_491),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_526),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_542),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_529),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_490),
.B(n_484),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_531),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_547),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_534),
.Y(n_562)
);

INVxp67_ASAP7_75t_SL g563 ( 
.A(n_520),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_512),
.B(n_426),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_513),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_522),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_522),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_552),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_500),
.B(n_466),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_524),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_527),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_527),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_505),
.B(n_495),
.Y(n_573)
);

XOR2x2_ASAP7_75t_L g574 ( 
.A(n_502),
.B(n_453),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_528),
.Y(n_575)
);

AND2x6_ASAP7_75t_L g576 ( 
.A(n_514),
.B(n_480),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_507),
.B(n_457),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_503),
.B(n_492),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_498),
.Y(n_579)
);

NAND2x1p5_ASAP7_75t_L g580 ( 
.A(n_514),
.B(n_481),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_512),
.B(n_440),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_546),
.B(n_481),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_497),
.B(n_470),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_546),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_535),
.B(n_483),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_517),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_554),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_536),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_519),
.B(n_462),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_510),
.Y(n_590)
);

INVxp33_ASAP7_75t_L g591 ( 
.A(n_516),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_515),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_515),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_543),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_506),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_509),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_544),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_538),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_496),
.B(n_462),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_499),
.B(n_483),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_530),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_550),
.B(n_298),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_537),
.B(n_436),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_553),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_545),
.B(n_441),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_538),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_539),
.Y(n_607)
);

INVx8_ASAP7_75t_L g608 ( 
.A(n_504),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_504),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_501),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_L g611 ( 
.A1(n_551),
.A2(n_401),
.B(n_399),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_525),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_540),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_518),
.B(n_416),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_521),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_508),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_540),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_523),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_533),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_501),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_541),
.B(n_549),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_493),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_532),
.Y(n_623)
);

BUFx5_ASAP7_75t_L g624 ( 
.A(n_592),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_599),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_593),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_L g627 ( 
.A1(n_597),
.A2(n_401),
.B(n_399),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_595),
.B(n_487),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_587),
.B(n_399),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_596),
.B(n_436),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_577),
.B(n_446),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_575),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_555),
.B(n_494),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_563),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_590),
.B(n_511),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g636 ( 
.A1(n_611),
.A2(n_401),
.B(n_445),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_603),
.B(n_532),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_616),
.B(n_401),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_560),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_562),
.Y(n_640)
);

NAND2x1p5_ASAP7_75t_L g641 ( 
.A(n_578),
.B(n_594),
.Y(n_641)
);

INVx3_ASAP7_75t_SL g642 ( 
.A(n_618),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_585),
.B(n_445),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_563),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_569),
.B(n_446),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_589),
.B(n_445),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_583),
.B(n_447),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_566),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_568),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_586),
.B(n_434),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_558),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_600),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_576),
.B(n_432),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_607),
.B(n_447),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_614),
.B(n_449),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_566),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_579),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_580),
.B(n_588),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_565),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_561),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_580),
.B(n_405),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_567),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_564),
.B(n_411),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_564),
.B(n_411),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_582),
.B(n_461),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_581),
.B(n_450),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_582),
.B(n_461),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_L g668 ( 
.A1(n_611),
.A2(n_438),
.B(n_442),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_556),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_584),
.B(n_570),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_557),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_615),
.B(n_609),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_567),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_574),
.B(n_469),
.Y(n_674)
);

OR2x2_ASAP7_75t_SL g675 ( 
.A(n_622),
.B(n_548),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_567),
.Y(n_676)
);

INVxp67_ASAP7_75t_SL g677 ( 
.A(n_605),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_602),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_559),
.B(n_469),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_608),
.Y(n_680)
);

INVxp67_ASAP7_75t_SL g681 ( 
.A(n_571),
.Y(n_681)
);

AND2x2_ASAP7_75t_SL g682 ( 
.A(n_614),
.B(n_548),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_632),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_631),
.B(n_573),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_631),
.B(n_591),
.Y(n_685)
);

AND2x6_ASAP7_75t_L g686 ( 
.A(n_638),
.B(n_598),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_665),
.B(n_572),
.Y(n_687)
);

NAND2x1_ASAP7_75t_L g688 ( 
.A(n_638),
.B(n_606),
.Y(n_688)
);

OR2x6_ASAP7_75t_L g689 ( 
.A(n_680),
.B(n_619),
.Y(n_689)
);

BUFx4f_ASAP7_75t_L g690 ( 
.A(n_642),
.Y(n_690)
);

BUFx5_ASAP7_75t_L g691 ( 
.A(n_626),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_677),
.B(n_612),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_674),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_639),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_626),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_648),
.Y(n_696)
);

AND2x6_ASAP7_75t_L g697 ( 
.A(n_638),
.B(n_613),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_675),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_639),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_650),
.B(n_617),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_640),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_SL g702 ( 
.A(n_642),
.B(n_601),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_625),
.B(n_604),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_640),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_637),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_650),
.B(n_621),
.Y(n_706)
);

OR2x6_ASAP7_75t_L g707 ( 
.A(n_652),
.B(n_608),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_667),
.B(n_610),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_651),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_634),
.B(n_299),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_SL g711 ( 
.A(n_682),
.B(n_620),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_645),
.B(n_623),
.Y(n_712)
);

OR2x6_ASAP7_75t_L g713 ( 
.A(n_652),
.B(n_608),
.Y(n_713)
);

OR2x6_ASAP7_75t_L g714 ( 
.A(n_641),
.B(n_469),
.Y(n_714)
);

OR2x6_ASAP7_75t_L g715 ( 
.A(n_641),
.B(n_474),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_644),
.B(n_300),
.Y(n_716)
);

NOR2xp67_ASAP7_75t_L g717 ( 
.A(n_672),
.B(n_301),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_648),
.Y(n_718)
);

INVx5_ASAP7_75t_L g719 ( 
.A(n_648),
.Y(n_719)
);

OR2x6_ASAP7_75t_SL g720 ( 
.A(n_679),
.B(n_304),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_651),
.Y(n_721)
);

INVx3_ASAP7_75t_SL g722 ( 
.A(n_708),
.Y(n_722)
);

INVxp67_ASAP7_75t_SL g723 ( 
.A(n_696),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_701),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_690),
.Y(n_725)
);

NAND2x1p5_ASAP7_75t_L g726 ( 
.A(n_719),
.B(n_655),
.Y(n_726)
);

BUFx2_ASAP7_75t_L g727 ( 
.A(n_693),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_701),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_693),
.Y(n_729)
);

BUFx4_ASAP7_75t_SL g730 ( 
.A(n_689),
.Y(n_730)
);

HB1xp67_ASAP7_75t_L g731 ( 
.A(n_705),
.Y(n_731)
);

BUFx2_ASAP7_75t_SL g732 ( 
.A(n_719),
.Y(n_732)
);

INVx6_ASAP7_75t_L g733 ( 
.A(n_719),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_684),
.B(n_633),
.Y(n_734)
);

NAND2x1p5_ASAP7_75t_L g735 ( 
.A(n_696),
.B(n_655),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_700),
.B(n_663),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_685),
.B(n_664),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_708),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_688),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_688),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_712),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_698),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_696),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_697),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_704),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_718),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_704),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_718),
.Y(n_748)
);

INVx6_ASAP7_75t_L g749 ( 
.A(n_718),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_698),
.Y(n_750)
);

OR2x6_ASAP7_75t_L g751 ( 
.A(n_714),
.B(n_715),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_694),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_724),
.Y(n_753)
);

HB1xp67_ASAP7_75t_L g754 ( 
.A(n_727),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_728),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_747),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_745),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_SL g758 ( 
.A1(n_734),
.A2(n_682),
.B1(n_706),
.B2(n_711),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_727),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_745),
.Y(n_760)
);

INVx8_ASAP7_75t_L g761 ( 
.A(n_746),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_736),
.A2(n_695),
.B1(n_692),
.B2(n_643),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_742),
.Y(n_763)
);

OAI22xp33_ASAP7_75t_L g764 ( 
.A1(n_741),
.A2(n_702),
.B1(n_678),
.B2(n_703),
.Y(n_764)
);

INVx6_ASAP7_75t_L g765 ( 
.A(n_733),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_SL g766 ( 
.A1(n_741),
.A2(n_635),
.B1(n_402),
.B2(n_636),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_752),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_752),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_737),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_735),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_750),
.B(n_647),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_739),
.A2(n_653),
.B(n_627),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_738),
.A2(n_635),
.B1(n_666),
.B2(n_661),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_738),
.A2(n_666),
.B1(n_661),
.B2(n_658),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_725),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_731),
.A2(n_666),
.B1(n_658),
.B2(n_697),
.Y(n_776)
);

CKINVDCx11_ASAP7_75t_R g777 ( 
.A(n_722),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_753),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_L g779 ( 
.A1(n_764),
.A2(n_751),
.B1(n_769),
.B2(n_722),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_766),
.B(n_758),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_758),
.A2(n_654),
.B1(n_717),
.B2(n_687),
.Y(n_781)
);

NAND3xp33_ASAP7_75t_L g782 ( 
.A(n_766),
.B(n_402),
.C(n_423),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_773),
.A2(n_654),
.B1(n_687),
.B2(n_714),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_774),
.A2(n_751),
.B1(n_729),
.B2(n_715),
.Y(n_784)
);

BUFx2_ASAP7_75t_L g785 ( 
.A(n_754),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_771),
.A2(n_654),
.B1(n_721),
.B2(n_709),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_765),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_768),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_757),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_L g790 ( 
.A1(n_776),
.A2(n_763),
.B1(n_759),
.B2(n_754),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_760),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_777),
.A2(n_660),
.B1(n_630),
.B2(n_683),
.Y(n_792)
);

AOI222xp33_ASAP7_75t_L g793 ( 
.A1(n_759),
.A2(n_628),
.B1(n_423),
.B2(n_668),
.C1(n_755),
.C2(n_756),
.Y(n_793)
);

AOI211xp5_ASAP7_75t_SL g794 ( 
.A1(n_762),
.A2(n_716),
.B(n_710),
.C(n_628),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_SL g795 ( 
.A1(n_770),
.A2(n_657),
.B1(n_744),
.B2(n_686),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_765),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_767),
.Y(n_797)
);

BUFx4f_ASAP7_75t_SL g798 ( 
.A(n_765),
.Y(n_798)
);

OAI22xp33_ASAP7_75t_L g799 ( 
.A1(n_772),
.A2(n_720),
.B1(n_713),
.B2(n_707),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_761),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_761),
.Y(n_801)
);

OAI222xp33_ASAP7_75t_L g802 ( 
.A1(n_758),
.A2(n_735),
.B1(n_726),
.B2(n_332),
.C1(n_305),
.C2(n_314),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_775),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_758),
.A2(n_669),
.B1(n_671),
.B2(n_659),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_758),
.A2(n_671),
.B1(n_669),
.B2(n_649),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_780),
.A2(n_793),
.B1(n_782),
.B2(n_779),
.Y(n_806)
);

OAI22xp33_ASAP7_75t_L g807 ( 
.A1(n_794),
.A2(n_713),
.B1(n_707),
.B2(n_726),
.Y(n_807)
);

AOI222xp33_ASAP7_75t_L g808 ( 
.A1(n_802),
.A2(n_670),
.B1(n_681),
.B2(n_323),
.C1(n_324),
.C2(n_629),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_789),
.B(n_743),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_792),
.A2(n_744),
.B1(n_689),
.B2(n_739),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_781),
.A2(n_691),
.B1(n_629),
.B2(n_670),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_789),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_785),
.B(n_699),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_784),
.A2(n_691),
.B1(n_670),
.B2(n_740),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_799),
.A2(n_740),
.B1(n_739),
.B2(n_697),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_785),
.B(n_723),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_791),
.B(n_743),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_783),
.A2(n_740),
.B1(n_646),
.B2(n_656),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_SL g819 ( 
.A1(n_795),
.A2(n_733),
.B1(n_732),
.B2(n_743),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_790),
.A2(n_662),
.B1(n_624),
.B2(n_477),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_788),
.B(n_746),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_791),
.B(n_797),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_804),
.A2(n_662),
.B1(n_624),
.B2(n_477),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_788),
.B(n_746),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_805),
.A2(n_624),
.B1(n_474),
.B2(n_477),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_SL g826 ( 
.A1(n_803),
.A2(n_748),
.B1(n_746),
.B2(n_749),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_786),
.A2(n_749),
.B1(n_748),
.B2(n_676),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_803),
.A2(n_787),
.B1(n_778),
.B2(n_797),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_787),
.B(n_748),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_798),
.A2(n_624),
.B1(n_485),
.B2(n_676),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_796),
.A2(n_624),
.B1(n_676),
.B2(n_673),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_796),
.A2(n_748),
.B1(n_676),
.B2(n_673),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_800),
.A2(n_801),
.B1(n_673),
.B2(n_730),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_801),
.A2(n_673),
.B1(n_421),
.B2(n_415),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_801),
.A2(n_421),
.B1(n_415),
.B2(n_408),
.Y(n_835)
);

NOR3xp33_ASAP7_75t_SL g836 ( 
.A(n_807),
.B(n_801),
.C(n_51),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_806),
.B(n_46),
.Y(n_837)
);

AOI21xp33_ASAP7_75t_SL g838 ( 
.A1(n_808),
.A2(n_59),
.B(n_61),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_822),
.B(n_65),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_812),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_828),
.B(n_70),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_816),
.B(n_73),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_813),
.B(n_77),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_815),
.B(n_833),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_809),
.B(n_80),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_819),
.A2(n_421),
.B1(n_415),
.B2(n_408),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_817),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_817),
.B(n_84),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_829),
.B(n_85),
.Y(n_849)
);

NAND3xp33_ASAP7_75t_L g850 ( 
.A(n_814),
.B(n_810),
.C(n_820),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_821),
.B(n_96),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_824),
.B(n_97),
.Y(n_852)
);

AND2x2_ASAP7_75t_SL g853 ( 
.A(n_831),
.B(n_102),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_826),
.B(n_107),
.Y(n_854)
);

AOI221xp5_ASAP7_75t_L g855 ( 
.A1(n_825),
.A2(n_408),
.B1(n_403),
.B2(n_400),
.C(n_114),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_811),
.A2(n_403),
.B1(n_400),
.B2(n_111),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_831),
.B(n_108),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_823),
.B(n_109),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_832),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_847),
.B(n_818),
.Y(n_860)
);

AOI221xp5_ASAP7_75t_L g861 ( 
.A1(n_838),
.A2(n_827),
.B1(n_830),
.B2(n_834),
.C(n_835),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_840),
.B(n_115),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_840),
.B(n_116),
.Y(n_863)
);

OR2x2_ASAP7_75t_L g864 ( 
.A(n_839),
.B(n_126),
.Y(n_864)
);

AO21x2_ASAP7_75t_L g865 ( 
.A1(n_836),
.A2(n_127),
.B(n_128),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_842),
.B(n_129),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_859),
.Y(n_867)
);

NAND4xp75_ASAP7_75t_L g868 ( 
.A(n_853),
.B(n_133),
.C(n_135),
.D(n_137),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_844),
.B(n_143),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_853),
.B(n_148),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_837),
.A2(n_403),
.B1(n_152),
.B2(n_153),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_845),
.B(n_151),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_857),
.B(n_156),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_844),
.B(n_158),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_848),
.B(n_162),
.Y(n_875)
);

NOR3xp33_ASAP7_75t_L g876 ( 
.A(n_837),
.B(n_165),
.C(n_166),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_867),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_867),
.Y(n_878)
);

NAND4xp75_ASAP7_75t_L g879 ( 
.A(n_869),
.B(n_841),
.C(n_854),
.D(n_843),
.Y(n_879)
);

NAND4xp75_ASAP7_75t_L g880 ( 
.A(n_869),
.B(n_849),
.C(n_855),
.D(n_852),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_874),
.B(n_850),
.Y(n_881)
);

XOR2x2_ASAP7_75t_L g882 ( 
.A(n_868),
.B(n_870),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_863),
.Y(n_883)
);

NAND4xp75_ASAP7_75t_SL g884 ( 
.A(n_870),
.B(n_846),
.C(n_856),
.D(n_851),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_860),
.Y(n_885)
);

OAI22x1_ASAP7_75t_L g886 ( 
.A1(n_874),
.A2(n_858),
.B1(n_856),
.B2(n_167),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_862),
.Y(n_887)
);

OAI22x1_ASAP7_75t_L g888 ( 
.A1(n_873),
.A2(n_168),
.B1(n_171),
.B2(n_173),
.Y(n_888)
);

XNOR2xp5_ASAP7_75t_L g889 ( 
.A(n_882),
.B(n_872),
.Y(n_889)
);

XOR2xp5_ASAP7_75t_L g890 ( 
.A(n_879),
.B(n_872),
.Y(n_890)
);

XOR2x2_ASAP7_75t_L g891 ( 
.A(n_881),
.B(n_876),
.Y(n_891)
);

XNOR2xp5_ASAP7_75t_L g892 ( 
.A(n_886),
.B(n_875),
.Y(n_892)
);

XNOR2xp5_ASAP7_75t_L g893 ( 
.A(n_884),
.B(n_875),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_880),
.A2(n_871),
.B1(n_864),
.B2(n_861),
.Y(n_894)
);

XNOR2xp5_ASAP7_75t_L g895 ( 
.A(n_888),
.B(n_866),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_877),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_885),
.Y(n_897)
);

XNOR2x1_ASAP7_75t_SL g898 ( 
.A(n_887),
.B(n_865),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_883),
.B(n_176),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_885),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_896),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_900),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_896),
.B(n_878),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_897),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_893),
.B(n_178),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_898),
.Y(n_906)
);

XOR2xp5_ASAP7_75t_L g907 ( 
.A(n_889),
.B(n_180),
.Y(n_907)
);

CKINVDCx8_ASAP7_75t_R g908 ( 
.A(n_899),
.Y(n_908)
);

AO22x2_ASAP7_75t_L g909 ( 
.A1(n_894),
.A2(n_182),
.B1(n_183),
.B2(n_187),
.Y(n_909)
);

OA22x2_ASAP7_75t_L g910 ( 
.A1(n_890),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_892),
.B(n_192),
.Y(n_911)
);

XNOR2xp5_ASAP7_75t_L g912 ( 
.A(n_891),
.B(n_193),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_901),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_903),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_902),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_904),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_913),
.Y(n_917)
);

AO22x2_ASAP7_75t_L g918 ( 
.A1(n_915),
.A2(n_906),
.B1(n_907),
.B2(n_911),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_914),
.Y(n_919)
);

NAND4xp75_ASAP7_75t_L g920 ( 
.A(n_916),
.B(n_905),
.C(n_909),
.D(n_910),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_919),
.Y(n_921)
);

AO22x2_ASAP7_75t_SL g922 ( 
.A1(n_920),
.A2(n_914),
.B1(n_912),
.B2(n_908),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_917),
.Y(n_923)
);

NOR2x1_ASAP7_75t_L g924 ( 
.A(n_921),
.B(n_918),
.Y(n_924)
);

NOR2x1_ASAP7_75t_L g925 ( 
.A(n_923),
.B(n_895),
.Y(n_925)
);

NOR4xp25_ASAP7_75t_L g926 ( 
.A(n_922),
.B(n_194),
.C(n_195),
.D(n_197),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_924),
.Y(n_927)
);

AO22x2_ASAP7_75t_L g928 ( 
.A1(n_927),
.A2(n_926),
.B1(n_925),
.B2(n_205),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_928),
.Y(n_929)
);

INVx2_ASAP7_75t_SL g930 ( 
.A(n_929),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_930),
.Y(n_931)
);

AO22x2_ASAP7_75t_L g932 ( 
.A1(n_931),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_932)
);

INVxp67_ASAP7_75t_SL g933 ( 
.A(n_932),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_SL g934 ( 
.A1(n_933),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_934),
.Y(n_935)
);

AOI221xp5_ASAP7_75t_L g936 ( 
.A1(n_935),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.C(n_224),
.Y(n_936)
);

AOI211xp5_ASAP7_75t_L g937 ( 
.A1(n_936),
.A2(n_229),
.B(n_230),
.C(n_232),
.Y(n_937)
);


endmodule