module fake_jpeg_29974_n_519 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_519);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_519;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_55),
.Y(n_137)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_8),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_59),
.B(n_66),
.Y(n_123)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_62),
.Y(n_147)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_63),
.Y(n_153)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_65),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_8),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_69),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_35),
.B(n_8),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_72),
.B(n_73),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_18),
.B(n_52),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_21),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_74),
.Y(n_107)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_18),
.B(n_9),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_77),
.B(n_86),
.Y(n_150)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_79),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx5_ASAP7_75t_SL g155 ( 
.A(n_82),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_19),
.B(n_7),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g140 ( 
.A(n_87),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_90),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_92),
.B(n_94),
.Y(n_157)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_7),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_33),
.B(n_10),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_100),
.Y(n_103)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_33),
.B(n_10),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_46),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_40),
.B(n_10),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_52),
.B1(n_40),
.B2(n_43),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_116),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_81),
.A2(n_49),
.B1(n_24),
.B2(n_27),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_54),
.A2(n_43),
.B1(n_22),
.B2(n_23),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_49),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_113),
.B(n_133),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_90),
.A2(n_24),
.B1(n_27),
.B2(n_38),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_118),
.B(n_28),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_55),
.A2(n_23),
.B1(n_22),
.B2(n_24),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_121),
.A2(n_131),
.B1(n_91),
.B2(n_88),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_80),
.A2(n_65),
.B(n_53),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_124),
.A2(n_56),
.B(n_63),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_SL g125 ( 
.A1(n_93),
.A2(n_23),
.B(n_26),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_159),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_L g131 ( 
.A1(n_61),
.A2(n_42),
.B1(n_38),
.B2(n_27),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_74),
.B(n_41),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_64),
.A2(n_24),
.B1(n_27),
.B2(n_38),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_135),
.A2(n_152),
.B1(n_87),
.B2(n_82),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_76),
.A2(n_68),
.B1(n_58),
.B2(n_82),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_62),
.B(n_41),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_123),
.A2(n_45),
.B1(n_30),
.B2(n_34),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_160),
.B(n_169),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_143),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_161),
.B(n_162),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_144),
.B(n_46),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_157),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_163),
.B(n_186),
.Y(n_226)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_164),
.Y(n_220)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_170),
.Y(n_223)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_171),
.Y(n_230)
);

AO22x2_ASAP7_75t_L g172 ( 
.A1(n_125),
.A2(n_83),
.B1(n_69),
.B2(n_70),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_172),
.B(n_190),
.Y(n_225)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_173),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_108),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_174),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_175),
.Y(n_233)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_176),
.Y(n_238)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_177),
.Y(n_232)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_178),
.Y(n_235)
);

OA22x2_ASAP7_75t_L g179 ( 
.A1(n_116),
.A2(n_71),
.B1(n_26),
.B2(n_97),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_179),
.B(n_194),
.Y(n_241)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_181),
.A2(n_208),
.B1(n_135),
.B2(n_139),
.Y(n_214)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_182),
.Y(n_248)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_126),
.Y(n_183)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_183),
.Y(n_258)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_136),
.Y(n_185)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_185),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_150),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_187),
.A2(n_212),
.B1(n_127),
.B2(n_34),
.Y(n_229)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_141),
.Y(n_188)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_189),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_103),
.A2(n_29),
.B(n_28),
.C(n_30),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_140),
.A2(n_29),
.B1(n_28),
.B2(n_30),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_191),
.A2(n_193),
.B(n_107),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_192),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_140),
.A2(n_29),
.B1(n_50),
.B2(n_45),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_131),
.B(n_101),
.Y(n_194)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_108),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_196),
.B(n_197),
.Y(n_251)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_198),
.B(n_201),
.Y(n_252)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_137),
.Y(n_199)
);

INVx11_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_105),
.A2(n_50),
.B1(n_45),
.B2(n_36),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_114),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_202),
.B(n_203),
.Y(n_255)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_117),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_204),
.B(n_207),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_107),
.B(n_75),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_205),
.B(n_206),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_127),
.B(n_50),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_137),
.A2(n_84),
.B1(n_79),
.B2(n_36),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_146),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_210),
.Y(n_218)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_146),
.Y(n_210)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_117),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_211),
.A2(n_171),
.B1(n_178),
.B2(n_175),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_152),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_213),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_214),
.A2(n_221),
.B1(n_228),
.B2(n_242),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_215),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_119),
.B1(n_139),
.B2(n_148),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_216),
.A2(n_239),
.B1(n_247),
.B2(n_249),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_190),
.A2(n_148),
.B1(n_147),
.B2(n_110),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_169),
.A2(n_36),
.B(n_34),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_229),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_166),
.A2(n_147),
.B1(n_138),
.B2(n_110),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_184),
.B(n_166),
.C(n_165),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_179),
.C(n_183),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_166),
.A2(n_129),
.B1(n_149),
.B2(n_153),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_184),
.A2(n_129),
.B1(n_120),
.B2(n_153),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_201),
.A2(n_129),
.B1(n_120),
.B2(n_38),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_172),
.A2(n_42),
.B1(n_128),
.B2(n_158),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_194),
.A2(n_158),
.B1(n_128),
.B2(n_42),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_250),
.A2(n_256),
.B1(n_195),
.B2(n_199),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_194),
.A2(n_172),
.B1(n_160),
.B2(n_179),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_167),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_259),
.B(n_263),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_225),
.B(n_172),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_225),
.B(n_173),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_268),
.Y(n_302)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_220),
.Y(n_265)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_265),
.Y(n_306)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_266),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_257),
.Y(n_267)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_267),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_217),
.B(n_164),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_238),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_269),
.B(n_272),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_218),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_271),
.B(n_275),
.Y(n_322)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_273),
.B(n_257),
.C(n_251),
.Y(n_314)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_274),
.B(n_276),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_218),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_244),
.B(n_217),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_235),
.Y(n_277)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_277),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_217),
.B(n_180),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_278),
.B(n_279),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_244),
.B(n_176),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_226),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_284),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_252),
.A2(n_179),
.B(n_198),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_281),
.A2(n_283),
.B(n_248),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_229),
.A2(n_213),
.B1(n_230),
.B2(n_235),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_282),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_182),
.Y(n_283)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_236),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_226),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_285),
.A2(n_296),
.B(n_299),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_286),
.A2(n_294),
.B1(n_228),
.B2(n_255),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_168),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_287),
.B(n_289),
.Y(n_312)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_220),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_288),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_253),
.B(n_177),
.Y(n_289)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_231),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_258),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_231),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_256),
.A2(n_188),
.B1(n_185),
.B2(n_174),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_255),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_295),
.B(n_297),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_251),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_219),
.B(n_189),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_258),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_298),
.A2(n_245),
.B1(n_240),
.B2(n_224),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_219),
.B(n_207),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_227),
.B(n_210),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_283),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_263),
.A2(n_290),
.B1(n_264),
.B2(n_275),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_301),
.A2(n_303),
.B1(n_304),
.B2(n_307),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_290),
.A2(n_241),
.B1(n_252),
.B2(n_214),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_271),
.A2(n_241),
.B1(n_249),
.B2(n_250),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_273),
.A2(n_241),
.B1(n_247),
.B2(n_242),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_309),
.A2(n_328),
.B1(n_330),
.B2(n_266),
.Y(n_355)
);

A2O1A1Ixp33_ASAP7_75t_SL g311 ( 
.A1(n_261),
.A2(n_230),
.B(n_255),
.C(n_257),
.Y(n_311)
);

OA22x2_ASAP7_75t_L g339 ( 
.A1(n_311),
.A2(n_267),
.B1(n_281),
.B2(n_261),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_259),
.B(n_251),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_313),
.B(n_314),
.C(n_329),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_315),
.Y(n_363)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_280),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_319),
.B(n_297),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_320),
.B(n_279),
.Y(n_356)
);

OAI21xp33_ASAP7_75t_SL g323 ( 
.A1(n_278),
.A2(n_254),
.B(n_233),
.Y(n_323)
);

XOR2x2_ASAP7_75t_SL g366 ( 
.A(n_323),
.B(n_51),
.Y(n_366)
);

OAI32xp33_ASAP7_75t_L g327 ( 
.A1(n_268),
.A2(n_222),
.A3(n_248),
.B1(n_223),
.B2(n_209),
.Y(n_327)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_327),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_286),
.A2(n_222),
.B1(n_223),
.B2(n_234),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_276),
.B(n_26),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_260),
.A2(n_234),
.B1(n_236),
.B2(n_232),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_332),
.B(n_298),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_285),
.A2(n_236),
.B1(n_232),
.B2(n_224),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_333),
.A2(n_335),
.B1(n_337),
.B2(n_338),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_262),
.A2(n_240),
.B1(n_245),
.B2(n_246),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_289),
.B(n_254),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_336),
.B(n_296),
.C(n_269),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_300),
.A2(n_246),
.B1(n_203),
.B2(n_211),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_260),
.A2(n_42),
.B1(n_233),
.B2(n_51),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_SL g379 ( 
.A1(n_339),
.A2(n_348),
.B(n_366),
.Y(n_379)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_317),
.Y(n_340)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_340),
.Y(n_376)
);

OA21x2_ASAP7_75t_L g341 ( 
.A1(n_322),
.A2(n_261),
.B(n_299),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_341),
.B(n_353),
.Y(n_378)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_317),
.Y(n_344)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_344),
.Y(n_394)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_326),
.Y(n_345)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_345),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_301),
.A2(n_294),
.B1(n_283),
.B2(n_270),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_347),
.A2(n_359),
.B1(n_328),
.B2(n_330),
.Y(n_387)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_308),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_349),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_334),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_350),
.B(n_354),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_352),
.B(n_351),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_312),
.B(n_287),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_334),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_355),
.A2(n_360),
.B1(n_372),
.B2(n_338),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_356),
.B(n_12),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_357),
.B(n_371),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_325),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_358),
.B(n_306),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_304),
.A2(n_274),
.B1(n_292),
.B2(n_272),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_309),
.A2(n_293),
.B1(n_291),
.B2(n_284),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_313),
.B(n_277),
.C(n_288),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_361),
.B(n_367),
.C(n_311),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_316),
.A2(n_265),
.B(n_98),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_362),
.Y(n_383)
);

OAI22x1_ASAP7_75t_L g364 ( 
.A1(n_316),
.A2(n_284),
.B1(n_12),
.B2(n_13),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g400 ( 
.A1(n_364),
.A2(n_6),
.B1(n_15),
.B2(n_14),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_303),
.A2(n_44),
.B1(n_51),
.B2(n_11),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_365),
.A2(n_324),
.B1(n_310),
.B2(n_331),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_305),
.B(n_44),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_318),
.Y(n_368)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_368),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_321),
.B(n_44),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_369),
.Y(n_375)
);

BUFx16f_ASAP7_75t_L g370 ( 
.A(n_325),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_335),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_318),
.A2(n_6),
.B(n_15),
.Y(n_371)
);

OAI22xp33_ASAP7_75t_L g372 ( 
.A1(n_302),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_374),
.B(n_391),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_381),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_382),
.B(n_385),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_384),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_355),
.A2(n_307),
.B1(n_336),
.B2(n_320),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_387),
.A2(n_388),
.B1(n_393),
.B2(n_343),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_342),
.A2(n_302),
.B1(n_324),
.B2(n_314),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_345),
.B(n_312),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_389),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_390),
.B(n_398),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_351),
.B(n_329),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_368),
.B(n_337),
.Y(n_392)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_392),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_342),
.A2(n_327),
.B1(n_315),
.B2(n_311),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_341),
.B(n_311),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_395),
.B(n_396),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_341),
.B(n_11),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_397),
.B(n_371),
.Y(n_415)
);

FAx1_ASAP7_75t_SL g398 ( 
.A(n_353),
.B(n_311),
.CI(n_6),
.CON(n_398),
.SN(n_398)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_400),
.B(n_375),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_352),
.B(n_16),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_401),
.B(n_403),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_343),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_402)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_402),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_403),
.B(n_369),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_391),
.C(n_361),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_404),
.B(n_405),
.C(n_421),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_396),
.B(n_363),
.C(n_344),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_406),
.A2(n_411),
.B1(n_382),
.B2(n_392),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_387),
.A2(n_360),
.B1(n_363),
.B2(n_366),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_380),
.A2(n_347),
.B(n_362),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_412),
.B(n_429),
.Y(n_441)
);

CKINVDCx14_ASAP7_75t_R g447 ( 
.A(n_415),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_416),
.B(n_427),
.Y(n_444)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_399),
.Y(n_417)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_417),
.Y(n_432)
);

XNOR2x2_ASAP7_75t_SL g418 ( 
.A(n_378),
.B(n_339),
.Y(n_418)
);

XOR2x2_ASAP7_75t_L g430 ( 
.A(n_418),
.B(n_379),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_388),
.B(n_339),
.C(n_367),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_422),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_386),
.B(n_349),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_423),
.B(n_424),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_399),
.B(n_370),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_394),
.Y(n_425)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_425),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_385),
.B(n_339),
.C(n_359),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_426),
.B(n_383),
.C(n_401),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_381),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_430),
.B(n_436),
.Y(n_462)
);

AOI21xp33_ASAP7_75t_L g433 ( 
.A1(n_408),
.A2(n_378),
.B(n_376),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_433),
.B(n_398),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_417),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_434),
.B(n_443),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_425),
.B(n_394),
.Y(n_435)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_435),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_437),
.B(n_448),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_411),
.A2(n_383),
.B1(n_373),
.B2(n_375),
.Y(n_438)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_438),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_404),
.B(n_373),
.C(n_395),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_442),
.B(n_405),
.C(n_426),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_407),
.B(n_429),
.Y(n_443)
);

NAND2xp33_ASAP7_75t_SL g445 ( 
.A(n_428),
.B(n_364),
.Y(n_445)
);

NOR2xp67_ASAP7_75t_R g460 ( 
.A(n_445),
.B(n_370),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_428),
.A2(n_402),
.B1(n_376),
.B2(n_346),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_446),
.A2(n_450),
.B1(n_413),
.B2(n_409),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_393),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_406),
.A2(n_409),
.B1(n_414),
.B2(n_413),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_464),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_447),
.A2(n_410),
.B1(n_346),
.B2(n_412),
.Y(n_452)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_452),
.Y(n_472)
);

FAx1_ASAP7_75t_SL g454 ( 
.A(n_443),
.B(n_418),
.CI(n_416),
.CON(n_454),
.SN(n_454)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_463),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_455),
.B(n_442),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_431),
.B(n_420),
.C(n_419),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_465),
.C(n_444),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_441),
.A2(n_407),
.B1(n_414),
.B2(n_410),
.Y(n_458)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_458),
.Y(n_476)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_460),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_441),
.A2(n_421),
.B1(n_365),
.B2(n_348),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_438),
.A2(n_358),
.B(n_420),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_464),
.A2(n_448),
.B(n_435),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_431),
.B(n_427),
.C(n_398),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_449),
.B(n_377),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_466),
.B(n_440),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_467),
.A2(n_439),
.B(n_436),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_468),
.A2(n_459),
.B(n_453),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_469),
.B(n_473),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_470),
.B(n_474),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_477),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_458),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_450),
.C(n_437),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_478),
.B(n_479),
.C(n_481),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_456),
.B(n_430),
.C(n_446),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_444),
.C(n_440),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_462),
.B(n_445),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_482),
.B(n_454),
.C(n_358),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_480),
.B(n_460),
.Y(n_483)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_483),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_481),
.B(n_471),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_485),
.B(n_491),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_472),
.B(n_462),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_486),
.B(n_489),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_476),
.A2(n_459),
.B1(n_457),
.B2(n_451),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_487),
.B(n_490),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_470),
.A2(n_457),
.B1(n_432),
.B2(n_463),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_478),
.A2(n_453),
.B1(n_432),
.B2(n_465),
.Y(n_491)
);

NOR2xp67_ASAP7_75t_L g492 ( 
.A(n_468),
.B(n_454),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_492),
.B(n_494),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_494),
.B(n_479),
.C(n_482),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_495),
.B(n_484),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_496),
.A2(n_501),
.B(n_502),
.Y(n_505)
);

XNOR2x1_ASAP7_75t_L g506 ( 
.A(n_498),
.B(n_488),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_493),
.B(n_475),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_493),
.B(n_369),
.C(n_372),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_503),
.A2(n_486),
.B1(n_489),
.B2(n_483),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_506),
.B(n_507),
.C(n_510),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_497),
.A2(n_496),
.B(n_504),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_508),
.B(n_509),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_504),
.A2(n_13),
.B(n_1),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_500),
.A2(n_0),
.B(n_3),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_505),
.B(n_499),
.C(n_4),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_513),
.A2(n_3),
.B(n_4),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_511),
.A2(n_3),
.B(n_4),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_514),
.B(n_515),
.C(n_512),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_516),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_517),
.B(n_3),
.C(n_5),
.Y(n_518)
);

BUFx24_ASAP7_75t_SL g519 ( 
.A(n_518),
.Y(n_519)
);


endmodule