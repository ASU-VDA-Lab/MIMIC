module real_jpeg_30320_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g200 ( 
.A(n_0),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_0),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_0),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_0),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_1),
.A2(n_267),
.B1(n_270),
.B2(n_271),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_1),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_1),
.A2(n_270),
.B1(n_326),
.B2(n_329),
.Y(n_325)
);

OAI22xp33_ASAP7_75t_L g425 ( 
.A1(n_1),
.A2(n_270),
.B1(n_426),
.B2(n_428),
.Y(n_425)
);

OAI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_1),
.A2(n_270),
.B1(n_458),
.B2(n_460),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_2),
.B(n_535),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_2),
.A2(n_532),
.B1(n_539),
.B2(n_542),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_3),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_3),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_3),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_5),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_5),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_5),
.Y(n_207)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_5),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_6),
.A2(n_114),
.B1(n_120),
.B2(n_121),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_6),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_6),
.A2(n_120),
.B1(n_168),
.B2(n_172),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_6),
.A2(n_120),
.B1(n_219),
.B2(n_222),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_6),
.A2(n_120),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_7),
.A2(n_40),
.B1(n_44),
.B2(n_48),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_7),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_7),
.A2(n_48),
.B1(n_103),
.B2(n_107),
.Y(n_102)
);

AO22x1_ASAP7_75t_L g209 ( 
.A1(n_7),
.A2(n_48),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_7),
.B(n_153),
.Y(n_384)
);

NAND2xp33_ASAP7_75t_SL g417 ( 
.A(n_7),
.B(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_7),
.B(n_24),
.Y(n_453)
);

OAI32xp33_ASAP7_75t_L g469 ( 
.A1(n_7),
.A2(n_470),
.A3(n_472),
.B1(n_473),
.B2(n_479),
.Y(n_469)
);

INVxp33_ASAP7_75t_L g535 ( 
.A(n_8),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_9),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_9),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_10),
.Y(n_127)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_10),
.Y(n_133)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_11),
.Y(n_485)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_12),
.Y(n_129)
);

AO22x1_ASAP7_75t_SL g51 ( 
.A1(n_13),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_13),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_13),
.A2(n_56),
.B1(n_122),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_13),
.A2(n_56),
.B1(n_219),
.B2(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_13),
.A2(n_56),
.B1(n_205),
.B2(n_257),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_188),
.B(n_526),
.C(n_536),
.Y(n_14)
);

HB1xp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_16),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_178),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_17),
.B(n_178),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_150),
.C(n_162),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_18),
.A2(n_150),
.B1(n_164),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_18),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_111),
.B1(n_112),
.B2(n_149),
.Y(n_18)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_19),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_76),
.B2(n_110),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_21),
.Y(n_187)
);

NOR2x1_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_49),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_23),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_38),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_24),
.B(n_51),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_24),
.A2(n_49),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_24),
.B(n_325),
.Y(n_367)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g183 ( 
.A1(n_25),
.A2(n_39),
.B(n_62),
.Y(n_183)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AO21x2_ASAP7_75t_L g62 ( 
.A1(n_26),
.A2(n_63),
.B(n_70),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_30),
.B1(n_33),
.B2(n_36),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_27),
.A2(n_93),
.B1(n_97),
.B2(n_100),
.Y(n_92)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_29),
.Y(n_427)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_37),
.Y(n_221)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2x1_ASAP7_75t_L g263 ( 
.A(n_39),
.B(n_62),
.Y(n_263)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AO22x2_ASAP7_75t_L g125 ( 
.A1(n_46),
.A2(n_126),
.B1(n_128),
.B2(n_130),
.Y(n_125)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_47),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_48),
.A2(n_156),
.B(n_158),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_48),
.B(n_159),
.Y(n_158)
);

AOI32xp33_ASAP7_75t_L g412 ( 
.A1(n_48),
.A2(n_413),
.A3(n_415),
.B1(n_416),
.B2(n_417),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_48),
.B(n_474),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_48),
.B(n_501),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_48),
.B(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_50),
.B(n_367),
.Y(n_366)
);

NAND2x1_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_61),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_53),
.Y(n_338)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_61),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_61),
.B(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_64),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_64),
.Y(n_415)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_66),
.Y(n_171)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVxp33_ASAP7_75t_L g416 ( 
.A(n_70),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_76),
.B(n_164),
.C(n_165),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_R g186 ( 
.A(n_76),
.B(n_111),
.C(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_76),
.A2(n_110),
.B1(n_166),
.B2(n_195),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g365 ( 
.A(n_76),
.B(n_366),
.C(n_368),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_76),
.A2(n_110),
.B1(n_366),
.B2(n_378),
.Y(n_377)
);

OA21x2_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_91),
.B(n_102),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_77),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_77),
.B(n_102),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_77),
.B(n_218),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_77),
.B(n_425),
.Y(n_438)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_92),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_78),
.Y(n_501)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_85),
.B2(n_87),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_84),
.Y(n_459)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_84),
.Y(n_462)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_87),
.Y(n_303)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_90),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_91),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_91),
.B(n_226),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_91),
.B(n_102),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_91),
.B(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_106),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_106),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_106),
.Y(n_430)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_109),
.Y(n_422)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_124),
.B(n_134),
.Y(n_112)
);

OAI21x1_ASAP7_75t_SL g180 ( 
.A1(n_113),
.A2(n_151),
.B(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_119),
.Y(n_345)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_124),
.B(n_181),
.Y(n_234)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2x1p5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_125),
.B(n_266),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_127),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_127),
.Y(n_350)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_129),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_134),
.B(n_274),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_135),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_140),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_138),
.A2(n_142),
.B1(n_144),
.B2(n_147),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_139),
.Y(n_269)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_139),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_140),
.B(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_150),
.A2(n_164),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_152),
.B(n_265),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_153),
.B(n_155),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_154),
.B(n_309),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_155),
.B(n_234),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_158),
.Y(n_355)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_163),
.B(n_244),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_175),
.B(n_176),
.Y(n_166)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_167),
.Y(n_238)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_176),
.B(n_324),
.Y(n_382)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NOR2x1_ASAP7_75t_L g262 ( 
.A(n_177),
.B(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_186),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_180),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_180),
.B(n_184),
.C(n_186),
.Y(n_530)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

INVxp67_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2x1_ASAP7_75t_L g315 ( 
.A(n_183),
.B(n_308),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_184),
.B(n_296),
.C(n_308),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_188),
.A2(n_537),
.B(n_541),
.Y(n_536)
);

AO21x2_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_283),
.B(n_522),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_242),
.B1(n_246),
.B2(n_279),
.Y(n_189)
);

INVxp33_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NOR2x1_ASAP7_75t_L g523 ( 
.A(n_191),
.B(n_243),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_191),
.B(n_243),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_196),
.C(n_235),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_192),
.A2(n_235),
.B1(n_236),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_192),
.Y(n_282)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_196),
.B(n_281),
.Y(n_280)
);

OAI21xp33_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_215),
.B(n_232),
.Y(n_196)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_197),
.B(n_233),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_197),
.A2(n_216),
.B1(n_231),
.B2(n_294),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_197),
.B(n_412),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_197),
.A2(n_231),
.B1(n_412),
.B2(n_444),
.Y(n_443)
);

AO21x2_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_201),
.B(n_208),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_198),
.A2(n_255),
.B(n_301),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_200),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_201),
.A2(n_301),
.B(n_304),
.Y(n_300)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_202),
.B(n_256),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_202),
.B(n_209),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_202),
.B(n_457),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx8_ASAP7_75t_L g496 ( 
.A(n_204),
.Y(n_496)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_205),
.Y(n_471)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_207),
.Y(n_259)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_207),
.Y(n_302)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_209),
.B(n_253),
.Y(n_252)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2x1_ASAP7_75t_L g277 ( 
.A(n_215),
.B(n_278),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_231),
.Y(n_215)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_216),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_224),
.B(n_225),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_221),
.Y(n_223)
);

INVx5_ASAP7_75t_L g472 ( 
.A(n_221),
.Y(n_472)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_225),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_225),
.B(n_424),
.Y(n_451)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVxp67_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp33_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

XOR2x2_ASAP7_75t_L g275 ( 
.A(n_237),
.B(n_239),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_240),
.B(n_424),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_241),
.B(n_250),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_241),
.B(n_438),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_SL g246 ( 
.A(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_247),
.B(n_280),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_275),
.C(n_276),
.Y(n_247)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_248),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_260),
.C(n_264),
.Y(n_248)
);

XNOR2x1_ASAP7_75t_L g290 ( 
.A(n_249),
.B(n_291),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_251),
.B(n_319),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.Y(n_251)
);

AND2x2_ASAP7_75t_SL g455 ( 
.A(n_252),
.B(n_456),
.Y(n_455)
);

BUFx4f_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_255),
.B(n_494),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_256),
.B(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_263),
.Y(n_441)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_264),
.Y(n_292)
);

NAND2x1_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_274),
.Y(n_264)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx4_ASAP7_75t_SL g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_275),
.B(n_277),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2x1p5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_403),
.Y(n_283)
);

OAI21x1_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_356),
.B(n_397),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_311),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_295),
.B2(n_310),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_288),
.B(n_295),
.Y(n_396)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_289),
.B(n_310),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_293),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_290),
.B(n_293),
.C(n_295),
.Y(n_399)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI22x1_ASAP7_75t_L g313 ( 
.A1(n_297),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_297),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_298),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_299),
.B(n_438),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_300),
.B(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_304),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_304),
.B(n_456),
.Y(n_502)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

AOI21x1_ASAP7_75t_L g394 ( 
.A1(n_311),
.A2(n_395),
.B(n_396),
.Y(n_394)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_317),
.C(n_320),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2x1_ASAP7_75t_L g360 ( 
.A(n_313),
.B(n_318),
.Y(n_360)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_315),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_320),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_321),
.A2(n_331),
.B(n_333),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_322),
.A2(n_332),
.B(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_323),
.A2(n_331),
.B1(n_332),
.B2(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_323),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_328),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_335),
.B(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

HAxp5_ASAP7_75t_SL g390 ( 
.A(n_336),
.B(n_337),
.CON(n_390),
.SN(n_390)
);

OAI31xp33_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_339),
.A3(n_342),
.B(n_346),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_351),
.B(n_355),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_352),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_372),
.B(n_394),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_361),
.Y(n_357)
);

NAND2x1p5_ASAP7_75t_L g373 ( 
.A(n_358),
.B(n_361),
.Y(n_373)
);

XNOR2x1_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_365),
.C(n_369),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_362),
.B(n_393),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_365),
.B(n_370),
.Y(n_393)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_366),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_367),
.B(n_441),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_368),
.B(n_377),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_373),
.B(n_520),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_392),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_375),
.B(n_392),
.Y(n_520)
);

OAI21xp33_ASAP7_75t_SL g375 ( 
.A1(n_376),
.A2(n_379),
.B(n_391),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_376),
.B(n_432),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_389),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_380),
.B(n_389),
.Y(n_391)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_381),
.B(n_390),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.C(n_385),
.Y(n_381)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_382),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_383),
.A2(n_384),
.B1(n_385),
.B2(n_386),
.Y(n_409)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

NOR2x1_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_387),
.Y(n_505)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

BUFx24_ASAP7_75t_SL g544 ( 
.A(n_390),
.Y(n_544)
);

NOR3xp33_ASAP7_75t_L g518 ( 
.A(n_394),
.B(n_398),
.C(n_519),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_398),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_399),
.B(n_400),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

AOI21x1_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_518),
.B(n_521),
.Y(n_403)
);

AO21x1_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_433),
.B(n_517),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_431),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_406),
.B(n_431),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_410),
.C(n_423),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_407),
.B(n_446),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_411),
.B(n_423),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_412),
.Y(n_444)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_434),
.A2(n_447),
.B(n_516),
.Y(n_433)
);

NOR2xp67_ASAP7_75t_SL g434 ( 
.A(n_435),
.B(n_445),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_435),
.B(n_445),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_439),
.C(n_442),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_436),
.A2(n_437),
.B1(n_439),
.B2(n_440),
.Y(n_464)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_443),
.B(n_464),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_465),
.B(n_515),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_463),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_L g515 ( 
.A(n_449),
.B(n_463),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_452),
.C(n_454),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_451),
.A2(n_452),
.B1(n_453),
.B2(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_451),
.Y(n_490)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_455),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_455),
.B(n_489),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_457),
.B(n_495),
.Y(n_494)
);

INVx6_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

BUFx12f_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_466),
.A2(n_491),
.B(n_514),
.Y(n_465)
);

NOR2x1_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_488),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_467),
.B(n_488),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_486),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_468),
.A2(n_469),
.B1(n_486),
.B2(n_487),
.Y(n_497)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_470),
.Y(n_507)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_472),
.Y(n_480)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_481),
.Y(n_479)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx4_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_492),
.A2(n_498),
.B(n_513),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_497),
.Y(n_492)
);

NOR2xp67_ASAP7_75t_SL g513 ( 
.A(n_493),
.B(n_497),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_505),
.Y(n_504)
);

INVx5_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_499),
.A2(n_503),
.B(n_512),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_502),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_502),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_504),
.B(n_506),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_508),
.Y(n_506)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_523),
.A2(n_524),
.B(n_525),
.Y(n_522)
);

NAND3xp33_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_532),
.C(n_533),
.Y(n_526)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_527),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_531),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_530),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_529),
.B(n_530),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_533),
.B(n_540),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_533),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_534),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_539),
.Y(n_537)
);


endmodule