module real_aes_11648_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_478;
wire n_356;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_693;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_936;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_142;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_756;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_498;
wire n_691;
wire n_481;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_928;
wire n_243;
wire n_899;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_926;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_166;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_888;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_0), .A2(n_105), .B1(n_937), .B2(n_944), .Y(n_104) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_1), .A2(n_85), .B1(n_600), .B2(n_601), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_2), .B(n_165), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_3), .B(n_206), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_4), .B(n_183), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g671 ( .A(n_5), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_6), .A2(n_40), .B1(n_155), .B2(n_598), .Y(n_627) );
NOR2xp67_ASAP7_75t_L g126 ( .A(n_7), .B(n_87), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_8), .B(n_157), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_9), .B(n_138), .Y(n_284) );
OAI22xp5_ASAP7_75t_SL g933 ( .A1(n_10), .A2(n_59), .B1(n_934), .B2(n_935), .Y(n_933) );
CKINVDCx5p33_ASAP7_75t_R g935 ( .A(n_10), .Y(n_935) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_11), .A2(n_66), .B1(n_155), .B2(n_235), .Y(n_651) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_12), .B(n_155), .C(n_158), .Y(n_592) );
NAND2x1p5_ASAP7_75t_L g219 ( .A(n_13), .B(n_138), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_14), .B(n_203), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g665 ( .A(n_15), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_16), .B(n_588), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_17), .B(n_145), .Y(n_635) );
AND2x2_ASAP7_75t_L g234 ( .A(n_18), .B(n_235), .Y(n_234) );
NAND3xp33_ASAP7_75t_L g589 ( .A(n_19), .B(n_151), .C(n_157), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_20), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_21), .A2(n_30), .B1(n_157), .B2(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_22), .B(n_588), .Y(n_614) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_23), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_24), .B(n_187), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_25), .A2(n_91), .B1(n_540), .B2(n_541), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_25), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_26), .A2(n_568), .B1(n_569), .B2(n_570), .Y(n_567) );
INVxp67_ASAP7_75t_SL g570 ( .A(n_26), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_26), .A2(n_570), .B1(n_573), .B2(n_574), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_27), .B(n_164), .Y(n_257) );
NAND2xp33_ASAP7_75t_L g214 ( .A(n_28), .B(n_215), .Y(n_214) );
NAND2xp33_ASAP7_75t_L g282 ( .A(n_29), .B(n_215), .Y(n_282) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_31), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_32), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_33), .B(n_693), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_34), .A2(n_55), .B1(n_215), .B2(n_235), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_35), .B(n_151), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_36), .B(n_182), .Y(n_218) );
INVx1_ASAP7_75t_L g125 ( .A(n_37), .Y(n_125) );
OAI21x1_ASAP7_75t_L g140 ( .A1(n_38), .A2(n_69), .B(n_141), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_39), .A2(n_150), .B(n_240), .C(n_242), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_41), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_42), .B(n_155), .Y(n_176) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_43), .Y(n_178) );
NAND2xp33_ASAP7_75t_L g207 ( .A(n_44), .B(n_201), .Y(n_207) );
AND2x6_ASAP7_75t_L g161 ( .A(n_45), .B(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g653 ( .A(n_46), .B(n_187), .Y(n_653) );
NAND2x1p5_ASAP7_75t_L g593 ( .A(n_47), .B(n_187), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_48), .B(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_49), .B(n_241), .Y(n_281) );
NAND2xp33_ASAP7_75t_L g256 ( .A(n_50), .B(n_201), .Y(n_256) );
XNOR2xp5_ASAP7_75t_L g568 ( .A(n_51), .B(n_128), .Y(n_568) );
XNOR2x1_ASAP7_75t_L g574 ( .A(n_51), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_52), .B(n_145), .Y(n_616) );
INVx1_ASAP7_75t_L g162 ( .A(n_53), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_54), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_56), .B(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_57), .B(n_187), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_58), .B(n_157), .Y(n_640) );
CKINVDCx5p33_ASAP7_75t_R g934 ( .A(n_59), .Y(n_934) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_60), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_61), .B(n_157), .Y(n_691) );
NAND2x1_ASAP7_75t_L g621 ( .A(n_62), .B(n_187), .Y(n_621) );
AND2x2_ASAP7_75t_L g244 ( .A(n_63), .B(n_164), .Y(n_244) );
AND2x2_ASAP7_75t_L g941 ( .A(n_64), .B(n_942), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_65), .B(n_158), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_67), .B(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_68), .B(n_685), .Y(n_684) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_70), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g688 ( .A(n_71), .Y(n_688) );
NAND2xp33_ASAP7_75t_L g144 ( .A(n_72), .B(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_73), .B(n_158), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_74), .A2(n_78), .B1(n_157), .B2(n_598), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_75), .B(n_206), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g675 ( .A(n_76), .Y(n_675) );
BUFx10_ASAP7_75t_L g117 ( .A(n_77), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_79), .B(n_175), .Y(n_279) );
INVx1_ASAP7_75t_SL g604 ( .A(n_80), .Y(n_604) );
NAND2xp33_ASAP7_75t_L g156 ( .A(n_81), .B(n_157), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_82), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_83), .B(n_215), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g620 ( .A(n_84), .Y(n_620) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_86), .Y(n_243) );
INVx2_ASAP7_75t_L g141 ( .A(n_88), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_89), .B(n_158), .Y(n_591) );
OR2x2_ASAP7_75t_L g122 ( .A(n_90), .B(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_90), .B(n_124), .Y(n_560) );
BUFx2_ASAP7_75t_L g566 ( .A(n_90), .Y(n_566) );
INVx1_ASAP7_75t_L g541 ( .A(n_91), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_92), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_93), .B(n_201), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_94), .B(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_95), .B(n_187), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_96), .Y(n_251) );
INVx1_ASAP7_75t_L g942 ( .A(n_97), .Y(n_942) );
INVx1_ASAP7_75t_L g233 ( .A(n_98), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_99), .Y(n_266) );
AND2x2_ASAP7_75t_L g274 ( .A(n_100), .B(n_138), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_101), .B(n_232), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_102), .B(n_164), .Y(n_163) );
OAI22xp5_ASAP7_75t_L g109 ( .A1(n_103), .A2(n_110), .B1(n_111), .B2(n_113), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_103), .Y(n_113) );
OR2x6_ASAP7_75t_L g105 ( .A(n_106), .B(n_561), .Y(n_105) );
OAI221xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_114), .B1(n_118), .B2(n_542), .C(n_553), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_114), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_109), .B(n_545), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_112), .B(n_603), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
BUFx12f_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_SL g559 ( .A(n_117), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_127), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx12f_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_122), .Y(n_547) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OR2x6_ASAP7_75t_L g931 ( .A(n_124), .B(n_559), .Y(n_931) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
OAI21xp33_ASAP7_75t_L g543 ( .A1(n_127), .A2(n_544), .B(n_548), .Y(n_543) );
XOR2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_539), .Y(n_127) );
NAND3x1_ASAP7_75t_L g128 ( .A(n_129), .B(n_402), .C(n_482), .Y(n_128) );
NOR4xp75_ASAP7_75t_L g129 ( .A(n_130), .B(n_323), .C(n_352), .D(n_378), .Y(n_129) );
NAND3x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_285), .C(n_307), .Y(n_130) );
OAI21xp5_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_189), .B(n_220), .Y(n_131) );
INVxp33_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_166), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_136), .B(n_312), .Y(n_342) );
OR2x2_ASAP7_75t_L g424 ( .A(n_136), .B(n_304), .Y(n_424) );
INVx2_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g299 ( .A(n_137), .Y(n_299) );
INVx1_ASAP7_75t_SL g384 ( .A(n_137), .Y(n_384) );
BUFx2_ASAP7_75t_L g449 ( .A(n_137), .Y(n_449) );
OA21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_142), .B(n_163), .Y(n_137) );
BUFx4f_ASAP7_75t_L g170 ( .A(n_138), .Y(n_170) );
OA21x2_ASAP7_75t_L g191 ( .A1(n_138), .A2(n_142), .B(n_163), .Y(n_191) );
INVx3_ASAP7_75t_L g197 ( .A(n_138), .Y(n_197) );
INVx4_ASAP7_75t_L g227 ( .A(n_138), .Y(n_227) );
OA21x2_ASAP7_75t_L g358 ( .A1(n_138), .A2(n_142), .B(n_163), .Y(n_358) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_138), .Y(n_707) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g188 ( .A(n_139), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_139), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g165 ( .A(n_140), .Y(n_165) );
OAI21x1_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_152), .B(n_159), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_147), .B(n_149), .Y(n_143) );
INVx2_ASAP7_75t_L g148 ( .A(n_145), .Y(n_148) );
INVx1_ASAP7_75t_L g175 ( .A(n_145), .Y(n_175) );
INVx2_ASAP7_75t_L g203 ( .A(n_145), .Y(n_203) );
INVx2_ASAP7_75t_L g600 ( .A(n_145), .Y(n_600) );
INVx1_ASAP7_75t_L g618 ( .A(n_145), .Y(n_618) );
INVx2_ASAP7_75t_L g673 ( .A(n_145), .Y(n_673) );
OR2x2_ASAP7_75t_L g674 ( .A(n_145), .B(n_675), .Y(n_674) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_146), .Y(n_155) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_146), .Y(n_157) );
INVx2_ASAP7_75t_L g183 ( .A(n_146), .Y(n_183) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_146), .Y(n_232) );
INVx1_ASAP7_75t_L g237 ( .A(n_146), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_149), .A2(n_213), .B(n_214), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_149), .A2(n_255), .B(n_256), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_149), .A2(n_184), .B1(n_597), .B2(n_599), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_149), .A2(n_273), .B1(n_627), .B2(n_628), .Y(n_626) );
OA22x2_ASAP7_75t_L g649 ( .A1(n_149), .A2(n_184), .B1(n_650), .B2(n_651), .Y(n_649) );
CKINVDCx6p67_ASAP7_75t_R g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_SL g267 ( .A(n_150), .Y(n_267) );
AOI21x1_ASAP7_75t_L g612 ( .A1(n_150), .A2(n_613), .B(n_614), .Y(n_612) );
AOI21x1_ASAP7_75t_L g634 ( .A1(n_150), .A2(n_635), .B(n_636), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g668 ( .A1(n_150), .A2(n_669), .B(n_674), .Y(n_668) );
INVx5_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx5_ASAP7_75t_L g158 ( .A(n_151), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_151), .A2(n_173), .B(n_174), .C(n_176), .Y(n_172) );
BUFx12f_ASAP7_75t_L g185 ( .A(n_151), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_151), .A2(n_638), .B1(n_639), .B2(n_640), .Y(n_637) );
OAI321xp33_ASAP7_75t_L g664 ( .A1(n_151), .A2(n_157), .A3(n_600), .B1(n_665), .B2(n_666), .C(n_667), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_156), .B(n_158), .Y(n_152) );
NOR2xp67_ASAP7_75t_L g265 ( .A(n_154), .B(n_266), .Y(n_265) );
INVx5_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g180 ( .A(n_157), .Y(n_180) );
INVx2_ASAP7_75t_L g206 ( .A(n_157), .Y(n_206) );
INVx2_ASAP7_75t_SL g241 ( .A(n_157), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_157), .B(n_264), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g687 ( .A1(n_157), .A2(n_158), .B(n_688), .C(n_689), .Y(n_687) );
AOI21x1_ASAP7_75t_L g199 ( .A1(n_158), .A2(n_200), .B(n_202), .Y(n_199) );
INVx1_ASAP7_75t_L g283 ( .A(n_158), .Y(n_283) );
OAI21x1_ASAP7_75t_L g171 ( .A1(n_159), .A2(n_172), .B(n_177), .Y(n_171) );
OAI21x1_ASAP7_75t_L g211 ( .A1(n_159), .A2(n_212), .B(n_216), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g249 ( .A1(n_159), .A2(n_250), .B(n_254), .Y(n_249) );
OAI21x1_ASAP7_75t_L g276 ( .A1(n_159), .A2(n_277), .B(n_280), .Y(n_276) );
AO31x2_ASAP7_75t_L g595 ( .A1(n_159), .A2(n_227), .A3(n_596), .B(n_602), .Y(n_595) );
AND2x2_ASAP7_75t_L g625 ( .A(n_159), .B(n_197), .Y(n_625) );
INVx8_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp67_ASAP7_75t_L g225 ( .A(n_160), .B(n_226), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_160), .A2(n_262), .B(n_268), .Y(n_261) );
INVx1_ASAP7_75t_L g648 ( .A(n_160), .Y(n_648) );
OAI21xp5_ASAP7_75t_L g676 ( .A1(n_160), .A2(n_667), .B(n_677), .Y(n_676) );
INVx8_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx2_ASAP7_75t_L g208 ( .A(n_161), .Y(n_208) );
OAI21x1_ASAP7_75t_L g584 ( .A1(n_161), .A2(n_585), .B(n_590), .Y(n_584) );
OAI21x1_ASAP7_75t_L g633 ( .A1(n_161), .A2(n_634), .B(n_637), .Y(n_633) );
INVx1_ASAP7_75t_L g695 ( .A(n_161), .Y(n_695) );
INVx2_ASAP7_75t_L g647 ( .A(n_164), .Y(n_647) );
BUFx5_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g603 ( .A(n_165), .Y(n_603) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_165), .Y(n_677) );
OR2x2_ASAP7_75t_L g437 ( .A(n_166), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_SL g401 ( .A(n_167), .B(n_367), .Y(n_401) );
NAND2xp33_ASAP7_75t_R g533 ( .A(n_167), .B(n_367), .Y(n_533) );
BUFx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_168), .B(n_358), .Y(n_364) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g351 ( .A(n_169), .B(n_313), .Y(n_351) );
OR2x2_ASAP7_75t_L g422 ( .A(n_169), .B(n_194), .Y(n_422) );
AND2x2_ASAP7_75t_L g471 ( .A(n_169), .B(n_304), .Y(n_471) );
OAI21x1_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_186), .Y(n_169) );
OA21x2_ASAP7_75t_L g210 ( .A1(n_170), .A2(n_211), .B(n_219), .Y(n_210) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_170), .A2(n_249), .B(n_257), .Y(n_248) );
OAI21x1_ASAP7_75t_L g302 ( .A1(n_170), .A2(n_171), .B(n_186), .Y(n_302) );
OAI21x1_ASAP7_75t_L g306 ( .A1(n_170), .A2(n_211), .B(n_219), .Y(n_306) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_181), .C(n_184), .Y(n_177) );
O2A1O1Ixp5_ASAP7_75t_L g216 ( .A1(n_179), .A2(n_184), .B(n_217), .C(n_218), .Y(n_216) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g201 ( .A(n_183), .Y(n_201) );
INVx2_ASAP7_75t_L g215 ( .A(n_183), .Y(n_215) );
O2A1O1Ixp5_ASAP7_75t_L g250 ( .A1(n_184), .A2(n_251), .B(n_252), .C(n_253), .Y(n_250) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_185), .A2(n_205), .B(n_207), .Y(n_204) );
BUFx2_ASAP7_75t_L g238 ( .A(n_185), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_185), .Y(n_273) );
AOI21x1_ASAP7_75t_L g615 ( .A1(n_185), .A2(n_616), .B(n_617), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_185), .A2(n_691), .B(n_692), .Y(n_690) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_189), .A2(n_473), .B1(n_478), .B2(n_480), .Y(n_472) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_192), .Y(n_189) );
AOI32xp33_ASAP7_75t_L g466 ( .A1(n_190), .A2(n_350), .A3(n_390), .B1(n_467), .B2(n_468), .Y(n_466) );
OAI322xp33_ASAP7_75t_L g483 ( .A1(n_190), .A2(n_484), .A3(n_485), .B1(n_486), .B2(n_489), .C1(n_492), .C2(n_494), .Y(n_483) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g311 ( .A(n_191), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g536 ( .A(n_191), .Y(n_536) );
INVx2_ASAP7_75t_L g438 ( .A(n_192), .Y(n_438) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_210), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_193), .B(n_304), .Y(n_345) );
INVx2_ASAP7_75t_L g416 ( .A(n_193), .Y(n_416) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g315 ( .A(n_194), .B(n_305), .Y(n_315) );
AND2x2_ASAP7_75t_L g367 ( .A(n_194), .B(n_306), .Y(n_367) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
OAI21x1_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_198), .B(n_209), .Y(n_195) );
OAI21x1_ASAP7_75t_L g275 ( .A1(n_196), .A2(n_276), .B(n_284), .Y(n_275) );
OAI21xp5_ASAP7_75t_L g313 ( .A1(n_196), .A2(n_198), .B(n_209), .Y(n_313) );
OAI21x1_ASAP7_75t_L g583 ( .A1(n_196), .A2(n_584), .B(n_593), .Y(n_583) );
OAI21x1_ASAP7_75t_L g656 ( .A1(n_196), .A2(n_584), .B(n_593), .Y(n_656) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OAI21x1_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_204), .B(n_208), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_201), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g252 ( .A(n_203), .Y(n_252) );
OAI21x1_ASAP7_75t_L g611 ( .A1(n_208), .A2(n_612), .B(n_615), .Y(n_611) );
INVx2_ASAP7_75t_L g341 ( .A(n_210), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_215), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_245), .Y(n_220) );
INVx2_ASAP7_75t_L g361 ( .A(n_221), .Y(n_361) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g293 ( .A(n_222), .B(n_260), .Y(n_293) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g330 ( .A(n_223), .B(n_260), .Y(n_330) );
AND2x2_ASAP7_75t_L g333 ( .A(n_223), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g370 ( .A(n_223), .Y(n_370) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g291 ( .A(n_224), .Y(n_291) );
AOI21x1_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_228), .B(n_244), .Y(n_224) );
OAI21x1_ASAP7_75t_L g610 ( .A1(n_226), .A2(n_611), .B(n_621), .Y(n_610) );
OAI21x1_ASAP7_75t_L g632 ( .A1(n_226), .A2(n_633), .B(n_641), .Y(n_632) );
OAI21x1_ASAP7_75t_L g701 ( .A1(n_226), .A2(n_633), .B(n_641), .Y(n_701) );
OAI21x1_ASAP7_75t_L g749 ( .A1(n_226), .A2(n_611), .B(n_621), .Y(n_749) );
INVx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_227), .A2(n_261), .B(n_274), .Y(n_260) );
AO21x2_ASAP7_75t_L g321 ( .A1(n_227), .A2(n_261), .B(n_274), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_239), .Y(n_228) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_234), .B(n_238), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_231), .B(n_233), .Y(n_230) );
NOR2xp33_ASAP7_75t_SL g271 ( .A(n_231), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g588 ( .A(n_232), .Y(n_588) );
INVx2_ASAP7_75t_L g598 ( .A(n_232), .Y(n_598) );
INVx2_ASAP7_75t_L g693 ( .A(n_232), .Y(n_693) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g601 ( .A(n_237), .Y(n_601) );
OAI21xp5_ASAP7_75t_L g590 ( .A1(n_240), .A2(n_591), .B(n_592), .Y(n_590) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx3_ASAP7_75t_L g518 ( .A(n_245), .Y(n_518) );
AND2x4_ASAP7_75t_L g245 ( .A(n_246), .B(n_258), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_247), .B(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g295 ( .A(n_247), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_247), .B(n_291), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_247), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_247), .B(n_258), .Y(n_400) );
AND2x2_ASAP7_75t_L g477 ( .A(n_247), .B(n_457), .Y(n_477) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g338 ( .A(n_248), .Y(n_338) );
AND2x2_ASAP7_75t_L g371 ( .A(n_248), .B(n_260), .Y(n_371) );
AND2x2_ASAP7_75t_L g308 ( .A(n_258), .B(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVxp67_ASAP7_75t_SL g287 ( .A(n_259), .Y(n_287) );
OR2x2_ASAP7_75t_L g347 ( .A(n_259), .B(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_275), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_265), .B(n_267), .Y(n_262) );
OAI21xp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_271), .B(n_273), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_273), .A2(n_278), .B(n_279), .Y(n_277) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_275), .Y(n_296) );
INVx1_ASAP7_75t_L g322 ( .A(n_275), .Y(n_322) );
INVx1_ASAP7_75t_L g337 ( .A(n_275), .Y(n_337) );
AND2x2_ASAP7_75t_L g369 ( .A(n_275), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g442 ( .A(n_275), .B(n_338), .Y(n_442) );
INVx1_ASAP7_75t_L g457 ( .A(n_275), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B(n_283), .Y(n_280) );
OAI21xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_292), .B(n_297), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_290), .B(n_427), .Y(n_481) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g348 ( .A(n_291), .Y(n_348) );
INVxp67_ASAP7_75t_SL g491 ( .A(n_291), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g343 ( .A1(n_292), .A2(n_344), .B1(n_346), .B2(n_349), .Y(n_343) );
AND2x4_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g381 ( .A(n_293), .Y(n_381) );
AND2x2_ASAP7_75t_L g467 ( .A(n_293), .B(n_434), .Y(n_467) );
NAND2xp67_ASAP7_75t_L g538 ( .A(n_293), .B(n_442), .Y(n_538) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g511 ( .A(n_295), .Y(n_511) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
OR2x2_ASAP7_75t_L g374 ( .A(n_299), .B(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g498 ( .A(n_299), .B(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_300), .B(n_464), .Y(n_463) );
NAND2x1_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx1_ASAP7_75t_L g317 ( .A(n_301), .Y(n_317) );
AND2x4_ASAP7_75t_SL g415 ( .A(n_301), .B(n_416), .Y(n_415) );
BUFx2_ASAP7_75t_L g485 ( .A(n_301), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_301), .B(n_341), .Y(n_499) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g388 ( .A(n_302), .Y(n_388) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_302), .Y(n_431) );
INVx1_ASAP7_75t_L g517 ( .A(n_303), .Y(n_517) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g414 ( .A(n_304), .B(n_358), .Y(n_414) );
AND2x2_ASAP7_75t_L g460 ( .A(n_304), .B(n_358), .Y(n_460) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_311), .B1(n_314), .B2(n_318), .Y(n_307) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_309), .Y(n_520) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g319 ( .A(n_310), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g464 ( .A(n_312), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_312), .B(n_396), .Y(n_503) );
BUFx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g375 ( .A(n_315), .Y(n_375) );
AND2x4_ASAP7_75t_L g386 ( .A(n_315), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g447 ( .A(n_315), .B(n_448), .Y(n_447) );
O2A1O1Ixp5_ASAP7_75t_L g516 ( .A1(n_316), .A2(n_374), .B(n_517), .C(n_518), .Y(n_516) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_319), .B(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx2_ASAP7_75t_SL g334 ( .A(n_321), .Y(n_334) );
INVx1_ASAP7_75t_L g393 ( .A(n_321), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_321), .B(n_338), .Y(n_427) );
INVx1_ASAP7_75t_L g329 ( .A(n_322), .Y(n_329) );
OAI21xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_339), .B(n_343), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2x1_ASAP7_75t_SL g325 ( .A(n_326), .B(n_331), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_328), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g529 ( .A(n_329), .B(n_333), .Y(n_529) );
AND2x2_ASAP7_75t_L g376 ( .A(n_330), .B(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g418 ( .A(n_330), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_330), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_330), .B(n_435), .Y(n_446) );
AND2x2_ASAP7_75t_L g461 ( .A(n_330), .B(n_442), .Y(n_461) );
OAI221xp5_ASAP7_75t_L g495 ( .A1(n_331), .A2(n_347), .B1(n_496), .B2(n_498), .C(n_500), .Y(n_495) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
AND2x4_ASAP7_75t_L g441 ( .A(n_333), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g493 ( .A(n_333), .B(n_435), .Y(n_493) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_334), .Y(n_409) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g377 ( .A(n_336), .Y(n_377) );
INVx1_ASAP7_75t_L g410 ( .A(n_336), .Y(n_410) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
BUFx3_ASAP7_75t_L g435 ( .A(n_338), .Y(n_435) );
OR2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
AND2x2_ASAP7_75t_L g349 ( .A(n_340), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2x1p5_ASAP7_75t_L g356 ( .A(n_341), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_344), .B(n_363), .Y(n_479) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g444 ( .A(n_345), .B(n_431), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_346), .A2(n_443), .B1(n_532), .B2(n_537), .Y(n_531) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g475 ( .A(n_348), .Y(n_475) );
AND2x2_ASAP7_75t_L g487 ( .A(n_350), .B(n_488), .Y(n_487) );
BUFx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_351), .B(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g398 ( .A(n_351), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_372), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_359), .B1(n_362), .B2(n_368), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g515 ( .A(n_356), .Y(n_515) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVxp67_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
INVxp67_ASAP7_75t_L g451 ( .A(n_363), .Y(n_451) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g469 ( .A(n_365), .Y(n_469) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g526 ( .A(n_367), .B(n_387), .Y(n_526) );
AND2x2_ASAP7_75t_L g530 ( .A(n_367), .B(n_449), .Y(n_530) );
AND2x4_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
INVx1_ASAP7_75t_L g394 ( .A(n_369), .Y(n_394) );
AND2x2_ASAP7_75t_L g523 ( .A(n_369), .B(n_393), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_376), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI32xp33_ASAP7_75t_L g458 ( .A1(n_376), .A2(n_459), .A3(n_460), .B1(n_461), .B2(n_462), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_382), .B(n_389), .Y(n_378) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR2x1p5_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_L g396 ( .A(n_384), .Y(n_396) );
INVx3_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g514 ( .A(n_387), .Y(n_514) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_395), .B1(n_399), .B2(n_401), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_392), .Y(n_452) );
INVx1_ASAP7_75t_L g512 ( .A(n_393), .Y(n_512) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NOR3xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_439), .C(n_465), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_404), .B(n_425), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_411), .B1(n_417), .B2(n_419), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_407), .B(n_410), .Y(n_406) );
INVxp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g506 ( .A(n_408), .Y(n_506) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVxp67_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_413), .B(n_415), .Y(n_412) );
AND2x4_ASAP7_75t_L g501 ( .A(n_413), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g488 ( .A(n_414), .Y(n_488) );
INVx2_ASAP7_75t_L g459 ( .A(n_415), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_415), .B(n_535), .Y(n_534) );
BUFx2_ASAP7_75t_L g454 ( .A(n_416), .Y(n_454) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NAND2x1_ASAP7_75t_SL g420 ( .A(n_421), .B(n_423), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g429 ( .A(n_424), .B(n_430), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_428), .B1(n_432), .B2(n_436), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_431), .Y(n_502) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g535 ( .A(n_435), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_458), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_443), .B1(n_445), .B2(n_447), .C(n_450), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_442), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g505 ( .A(n_442), .Y(n_505) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NOR4xp25_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .C(n_453), .D(n_455), .Y(n_450) );
INVxp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g484 ( .A(n_456), .B(n_481), .Y(n_484) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g494 ( .A(n_460), .Y(n_494) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_472), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NOR3xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_495), .C(n_507), .Y(n_482) );
AND2x2_ASAP7_75t_L g497 ( .A(n_485), .B(n_488), .Y(n_497) );
INVxp67_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OAI21xp33_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_503), .B(n_504), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
NAND3xp33_ASAP7_75t_SL g507 ( .A(n_508), .B(n_519), .C(n_531), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_513), .B(n_516), .Y(n_508) );
INVxp67_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_511), .B(n_512), .Y(n_510) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
O2A1O1Ixp5_ASAP7_75t_SL g519 ( .A1(n_520), .A2(n_521), .B(n_524), .C(n_527), .Y(n_519) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2x1p5_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
INVxp67_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx6_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx5_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx4_ASAP7_75t_L g552 ( .A(n_547), .Y(n_552) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NOR2xp33_ASAP7_75t_SL g553 ( .A(n_549), .B(n_554), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
INVx5_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NOR2xp33_ASAP7_75t_R g554 ( .A(n_555), .B(n_556), .Y(n_554) );
BUFx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx12f_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx1_ASAP7_75t_L g943 ( .A(n_560), .Y(n_943) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B1(n_928), .B2(n_936), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OAI21x1_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_567), .B(n_571), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_564), .B(n_572), .Y(n_571) );
BUFx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
BUFx8_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g569 ( .A(n_568), .Y(n_569) );
INVx2_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
NAND2x1p5_ASAP7_75t_L g575 ( .A(n_576), .B(n_851), .Y(n_575) );
NOR2x1_ASAP7_75t_L g576 ( .A(n_577), .B(n_777), .Y(n_576) );
NAND3xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_713), .C(n_751), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_579), .B(n_678), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_605), .B1(n_642), .B2(n_657), .Y(n_579) );
OR2x2_ASAP7_75t_L g736 ( .A(n_580), .B(n_715), .Y(n_736) );
NOR2x1p5_ASAP7_75t_L g876 ( .A(n_580), .B(n_841), .Y(n_876) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_594), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_582), .B(n_682), .Y(n_704) );
AND2x2_ASAP7_75t_L g760 ( .A(n_582), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g819 ( .A(n_582), .Y(n_819) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g816 ( .A(n_583), .B(n_706), .Y(n_816) );
OAI21xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B(n_589), .Y(n_585) );
INVxp67_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x4_ASAP7_75t_L g681 ( .A(n_594), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g839 ( .A(n_594), .Y(n_839) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_595), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g705 ( .A(n_595), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g718 ( .A(n_595), .Y(n_718) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_595), .Y(n_743) );
INVx1_ASAP7_75t_L g765 ( .A(n_595), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g685 ( .A(n_603), .Y(n_685) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_630), .Y(n_607) );
INVx2_ASAP7_75t_L g919 ( .A(n_608), .Y(n_919) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_622), .Y(n_608) );
INVx2_ASAP7_75t_L g797 ( .A(n_609), .Y(n_797) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g884 ( .A(n_610), .B(n_712), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g639 ( .A(n_618), .Y(n_639) );
INVx4_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_622), .B(n_660), .Y(n_659) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_622), .Y(n_699) );
INVx1_ASAP7_75t_L g757 ( .A(n_622), .Y(n_757) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g776 ( .A(n_623), .B(n_748), .Y(n_776) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_623), .Y(n_787) );
AND2x2_ASAP7_75t_L g790 ( .A(n_623), .B(n_663), .Y(n_790) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g711 ( .A(n_624), .Y(n_711) );
AOI21x1_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B(n_629), .Y(n_624) );
AND2x2_ASAP7_75t_L g859 ( .A(n_630), .B(n_803), .Y(n_859) );
INVx2_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g750 ( .A(n_631), .Y(n_750) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g660 ( .A(n_632), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_654), .Y(n_642) );
AND2x2_ASAP7_75t_L g863 ( .A(n_643), .B(n_864), .Y(n_863) );
AND2x2_ASAP7_75t_L g887 ( .A(n_643), .B(n_888), .Y(n_887) );
NAND2xp33_ASAP7_75t_SL g896 ( .A(n_643), .B(n_655), .Y(n_896) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVxp67_ASAP7_75t_L g759 ( .A(n_644), .Y(n_759) );
INVx1_ASAP7_75t_L g696 ( .A(n_645), .Y(n_696) );
INVx1_ASAP7_75t_L g716 ( .A(n_645), .Y(n_716) );
INVxp67_ASAP7_75t_SL g769 ( .A(n_645), .Y(n_769) );
INVx1_ASAP7_75t_L g810 ( .A(n_645), .Y(n_810) );
HB1xp67_ASAP7_75t_L g820 ( .A(n_645), .Y(n_820) );
OAI21x1_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_649), .B(n_652), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
OA21x2_ASAP7_75t_L g706 ( .A1(n_649), .A2(n_707), .B(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVxp67_ASAP7_75t_L g708 ( .A(n_653), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_654), .B(n_705), .Y(n_771) );
OR2x2_ASAP7_75t_L g847 ( .A(n_654), .B(n_848), .Y(n_847) );
AND2x4_ASAP7_75t_L g856 ( .A(n_654), .B(n_681), .Y(n_856) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_655), .B(n_718), .Y(n_794) );
NOR2xp67_ASAP7_75t_L g837 ( .A(n_655), .B(n_838), .Y(n_837) );
BUFx3_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g720 ( .A(n_656), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g744 ( .A(n_656), .B(n_683), .Y(n_744) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .Y(n_658) );
OR2x2_ASAP7_75t_L g874 ( .A(n_659), .B(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g785 ( .A(n_660), .Y(n_785) );
AND2x2_ASAP7_75t_L g905 ( .A(n_660), .B(n_739), .Y(n_905) );
INVxp67_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g700 ( .A(n_662), .B(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g725 ( .A(n_662), .B(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g732 ( .A(n_662), .B(n_711), .Y(n_732) );
OR2x2_ASAP7_75t_L g753 ( .A(n_662), .B(n_750), .Y(n_753) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g712 ( .A(n_663), .Y(n_712) );
OAI21x1_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_668), .B(n_676), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_697), .B1(n_702), .B2(n_709), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g846 ( .A1(n_679), .A2(n_847), .B(n_849), .Y(n_846) );
INVx3_ASAP7_75t_L g910 ( .A(n_679), .Y(n_910) );
OR2x6_ASAP7_75t_L g679 ( .A(n_680), .B(n_696), .Y(n_679) );
OR2x2_ASAP7_75t_L g927 ( .A(n_680), .B(n_818), .Y(n_927) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g848 ( .A(n_681), .Y(n_848) );
BUFx2_ASAP7_75t_L g872 ( .A(n_681), .Y(n_872) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g721 ( .A(n_683), .Y(n_721) );
NAND2x1p5_ASAP7_75t_L g683 ( .A(n_684), .B(n_686), .Y(n_683) );
OAI21x1_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_690), .B(n_694), .Y(n_686) );
AND2x2_ASAP7_75t_L g842 ( .A(n_696), .B(n_815), .Y(n_842) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
AND2x2_ASAP7_75t_L g883 ( .A(n_699), .B(n_884), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_700), .B(n_773), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_700), .B(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_700), .B(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g844 ( .A(n_700), .Y(n_844) );
INVx1_ASAP7_75t_L g726 ( .A(n_701), .Y(n_726) );
INVx2_ASAP7_75t_L g731 ( .A(n_701), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_702), .A2(n_874), .B1(n_925), .B2(n_927), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_705), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_703), .B(n_827), .Y(n_920) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AOI222xp33_ASAP7_75t_L g853 ( .A1(n_705), .A2(n_754), .B1(n_854), .B2(n_856), .C1(n_857), .C2(n_860), .Y(n_853) );
AND2x2_ASAP7_75t_L g793 ( .A(n_706), .B(n_761), .Y(n_793) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_710), .Y(n_735) );
AND2x4_ASAP7_75t_L g801 ( .A(n_710), .B(n_802), .Y(n_801) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_711), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_711), .B(n_731), .Y(n_909) );
INVx2_ASAP7_75t_L g739 ( .A(n_712), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_712), .B(n_756), .Y(n_926) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_722), .B1(n_733), .B2(n_745), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_717), .Y(n_714) );
AND2x2_ASAP7_75t_L g901 ( .A(n_715), .B(n_902), .Y(n_901) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NOR2x1_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
HB1xp67_ASAP7_75t_L g807 ( .A(n_718), .Y(n_807) );
INVx1_ASAP7_75t_L g827 ( .A(n_718), .Y(n_827) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g878 ( .A(n_720), .B(n_810), .Y(n_878) );
INVx2_ASAP7_75t_L g761 ( .A(n_721), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_728), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_723), .A2(n_812), .B1(n_817), .B2(n_821), .Y(n_811) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AOI321xp33_ASAP7_75t_L g751 ( .A1(n_724), .A2(n_752), .A3(n_754), .B1(n_758), .B2(n_762), .C(n_770), .Y(n_751) );
AND2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_727), .Y(n_724) );
INVx2_ASAP7_75t_L g918 ( .A(n_725), .Y(n_918) );
INVx1_ASAP7_75t_L g830 ( .A(n_727), .Y(n_830) );
INVxp67_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
NOR2xp67_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .Y(n_729) );
AND2x2_ASAP7_75t_L g822 ( .A(n_730), .B(n_790), .Y(n_822) );
AND2x2_ASAP7_75t_L g829 ( .A(n_730), .B(n_830), .Y(n_829) );
AND2x4_ASAP7_75t_L g870 ( .A(n_730), .B(n_739), .Y(n_870) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g850 ( .A(n_731), .B(n_790), .Y(n_850) );
OR2x2_ASAP7_75t_L g796 ( .A(n_732), .B(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g858 ( .A(n_732), .Y(n_858) );
OR2x2_ASAP7_75t_L g895 ( .A(n_732), .B(n_781), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_736), .B1(n_737), .B2(n_740), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
O2A1O1Ixp5_ASAP7_75t_L g828 ( .A1(n_738), .A2(n_807), .B(n_829), .C(n_831), .Y(n_828) );
BUFx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_744), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND2x1p5_ASAP7_75t_L g767 ( .A(n_744), .B(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g833 ( .A(n_744), .Y(n_833) );
INVx2_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
OR2x2_ASAP7_75t_L g840 ( .A(n_746), .B(n_789), .Y(n_840) );
OR2x2_ASAP7_75t_L g746 ( .A(n_747), .B(n_750), .Y(n_746) );
INVx1_ASAP7_75t_L g781 ( .A(n_747), .Y(n_781) );
BUFx2_ASAP7_75t_L g875 ( .A(n_747), .Y(n_875) );
AND2x2_ASAP7_75t_L g906 ( .A(n_747), .B(n_819), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_747), .B(n_750), .Y(n_913) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_748), .Y(n_832) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g756 ( .A(n_749), .Y(n_756) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
OR2x2_ASAP7_75t_L g891 ( .A(n_753), .B(n_776), .Y(n_891) );
BUFx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
INVxp67_ASAP7_75t_SL g773 ( .A(n_756), .Y(n_773) );
BUFx2_ASAP7_75t_L g900 ( .A(n_756), .Y(n_900) );
AND2x2_ASAP7_75t_L g845 ( .A(n_757), .B(n_797), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_758), .A2(n_779), .B1(n_791), .B2(n_795), .Y(n_778) );
AND2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
BUFx2_ASAP7_75t_L g916 ( .A(n_759), .Y(n_916) );
AND2x2_ASAP7_75t_L g808 ( .A(n_760), .B(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g894 ( .A(n_760), .Y(n_894) );
INVx2_ASAP7_75t_L g815 ( .A(n_761), .Y(n_815) );
AND2x2_ASAP7_75t_L g902 ( .A(n_761), .B(n_765), .Y(n_902) );
AND2x4_ASAP7_75t_L g762 ( .A(n_763), .B(n_766), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NOR2xp67_ASAP7_75t_L g814 ( .A(n_765), .B(n_815), .Y(n_814) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_767), .A2(n_771), .B1(n_772), .B2(n_774), .Y(n_770) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_775), .B(n_784), .Y(n_805) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
NAND3xp33_ASAP7_75t_L g777 ( .A(n_778), .B(n_798), .C(n_823), .Y(n_777) );
NAND3xp33_ASAP7_75t_SL g779 ( .A(n_780), .B(n_782), .C(n_788), .Y(n_779) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
NOR2xp67_ASAP7_75t_L g783 ( .A(n_784), .B(n_786), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g867 ( .A(n_789), .Y(n_867) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
AND2x2_ASAP7_75t_L g899 ( .A(n_790), .B(n_900), .Y(n_899) );
NOR2x1p5_ASAP7_75t_SL g791 ( .A(n_792), .B(n_794), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g825 ( .A(n_793), .Y(n_825) );
AND2x4_ASAP7_75t_L g836 ( .A(n_793), .B(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_796), .B(n_855), .Y(n_854) );
INVx2_ASAP7_75t_L g803 ( .A(n_797), .Y(n_803) );
AND2x2_ASAP7_75t_L g922 ( .A(n_797), .B(n_923), .Y(n_922) );
O2A1O1Ixp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_804), .B(n_806), .C(n_811), .Y(n_798) );
AOI21xp5_ASAP7_75t_L g886 ( .A1(n_799), .A2(n_887), .B(n_890), .Y(n_886) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
OR2x2_ASAP7_75t_L g908 ( .A(n_802), .B(n_909), .Y(n_908) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
AND2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_807), .B(n_893), .Y(n_892) );
INVx2_ASAP7_75t_L g882 ( .A(n_809), .Y(n_882) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
AND2x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_816), .Y(n_813) );
INVx1_ASAP7_75t_L g889 ( .A(n_815), .Y(n_889) );
AND2x2_ASAP7_75t_L g871 ( .A(n_816), .B(n_872), .Y(n_871) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
OR2x2_ASAP7_75t_L g861 ( .A(n_818), .B(n_827), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
O2A1O1Ixp5_ASAP7_75t_L g824 ( .A1(n_821), .A2(n_825), .B(n_826), .C(n_828), .Y(n_824) );
INVx2_ASAP7_75t_SL g821 ( .A(n_822), .Y(n_821) );
NOR3xp33_ASAP7_75t_L g823 ( .A(n_824), .B(n_834), .C(n_846), .Y(n_823) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g855 ( .A(n_829), .Y(n_855) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_833), .Y(n_831) );
INVx1_ASAP7_75t_L g864 ( .A(n_833), .Y(n_864) );
OAI22xp5_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_840), .B1(n_841), .B2(n_843), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVxp67_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_844), .B(n_845), .Y(n_843) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
NOR2x1_ASAP7_75t_L g851 ( .A(n_852), .B(n_885), .Y(n_851) );
NAND3xp33_ASAP7_75t_L g852 ( .A(n_853), .B(n_862), .C(n_877), .Y(n_852) );
NAND2x1p5_ASAP7_75t_L g880 ( .A(n_856), .B(n_881), .Y(n_880) );
AND2x2_ASAP7_75t_L g857 ( .A(n_858), .B(n_859), .Y(n_857) );
AOI222xp33_ASAP7_75t_L g862 ( .A1(n_859), .A2(n_863), .B1(n_865), .B2(n_871), .C1(n_873), .C2(n_876), .Y(n_862) );
INVx2_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
NOR2x1_ASAP7_75t_L g866 ( .A(n_867), .B(n_868), .Y(n_866) );
INVx2_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx4_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx2_ASAP7_75t_SL g873 ( .A(n_874), .Y(n_873) );
OAI21xp33_ASAP7_75t_L g877 ( .A1(n_878), .A2(n_879), .B(n_883), .Y(n_877) );
AOI211xp5_ASAP7_75t_L g911 ( .A1(n_879), .A2(n_912), .B(n_914), .C(n_924), .Y(n_911) );
INVx2_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx2_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
NAND3xp33_ASAP7_75t_L g885 ( .A(n_886), .B(n_897), .C(n_911), .Y(n_885) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_891), .A2(n_892), .B1(n_895), .B2(n_896), .Y(n_890) );
INVx2_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
AND2x2_ASAP7_75t_L g897 ( .A(n_898), .B(n_903), .Y(n_897) );
NAND2x1p5_ASAP7_75t_L g898 ( .A(n_899), .B(n_901), .Y(n_898) );
OAI21xp5_ASAP7_75t_L g903 ( .A1(n_904), .A2(n_907), .B(n_910), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_905), .B(n_906), .Y(n_904) );
INVx2_ASAP7_75t_SL g907 ( .A(n_908), .Y(n_907) );
INVx1_ASAP7_75t_SL g923 ( .A(n_909), .Y(n_923) );
INVxp67_ASAP7_75t_SL g912 ( .A(n_913), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g914 ( .A1(n_915), .A2(n_917), .B1(n_920), .B2(n_921), .Y(n_914) );
INVx2_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
OR2x2_ASAP7_75t_L g917 ( .A(n_918), .B(n_919), .Y(n_917) );
INVx2_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
HB1xp67_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_929), .B(n_932), .Y(n_928) );
NAND2xp5_ASAP7_75t_SL g936 ( .A(n_929), .B(n_933), .Y(n_936) );
INVxp33_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
BUFx2_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
CKINVDCx5p33_ASAP7_75t_R g932 ( .A(n_933), .Y(n_932) );
INVx2_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
BUFx12f_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
BUFx12f_ASAP7_75t_L g948 ( .A(n_940), .Y(n_948) );
AND2x4_ASAP7_75t_L g940 ( .A(n_941), .B(n_943), .Y(n_940) );
HB1xp67_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx2_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
endmodule