module fake_netlist_1_11119_n_45 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_45);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_30;
wire n_16;
wire n_26;
wire n_25;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
BUFx6f_ASAP7_75t_L g16 ( .A(n_12), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_4), .Y(n_17) );
INVx3_ASAP7_75t_L g18 ( .A(n_3), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_7), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_3), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_8), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_11), .Y(n_22) );
BUFx6f_ASAP7_75t_L g23 ( .A(n_14), .Y(n_23) );
INVx1_ASAP7_75t_SL g24 ( .A(n_19), .Y(n_24) );
BUFx4f_ASAP7_75t_L g25 ( .A(n_16), .Y(n_25) );
AND2x4_ASAP7_75t_L g26 ( .A(n_18), .B(n_0), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_18), .Y(n_27) );
BUFx2_ASAP7_75t_L g28 ( .A(n_24), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
INVx2_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
OAI33xp33_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_27), .A3(n_20), .B1(n_17), .B2(n_19), .B3(n_22), .Y(n_32) );
OR2x2_ASAP7_75t_L g33 ( .A(n_31), .B(n_28), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_33), .Y(n_34) );
AOI22xp33_ASAP7_75t_SL g35 ( .A1(n_32), .A2(n_26), .B1(n_17), .B2(n_22), .Y(n_35) );
AOI22xp5_ASAP7_75t_L g36 ( .A1(n_34), .A2(n_26), .B1(n_21), .B2(n_23), .Y(n_36) );
NOR2xp67_ASAP7_75t_L g37 ( .A(n_34), .B(n_0), .Y(n_37) );
AOI211xp5_ASAP7_75t_L g38 ( .A1(n_35), .A2(n_23), .B(n_16), .C(n_4), .Y(n_38) );
AOI21xp33_ASAP7_75t_SL g39 ( .A1(n_36), .A2(n_1), .B(n_2), .Y(n_39) );
NAND3x1_ASAP7_75t_L g40 ( .A(n_37), .B(n_1), .C(n_2), .Y(n_40) );
AOI211x1_ASAP7_75t_SL g41 ( .A1(n_38), .A2(n_23), .B(n_16), .C(n_5), .Y(n_41) );
NOR3xp33_ASAP7_75t_L g42 ( .A(n_39), .B(n_5), .C(n_25), .Y(n_42) );
AOI221xp5_ASAP7_75t_L g43 ( .A1(n_41), .A2(n_25), .B1(n_9), .B2(n_10), .C(n_13), .Y(n_43) );
OAI21xp5_ASAP7_75t_SL g44 ( .A1(n_42), .A2(n_43), .B(n_40), .Y(n_44) );
AOI22x1_ASAP7_75t_L g45 ( .A1(n_44), .A2(n_6), .B1(n_15), .B2(n_25), .Y(n_45) );
endmodule