module fake_jpeg_3677_n_108 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_33),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_44),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_38),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_30),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_30),
.B(n_34),
.C(n_29),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_51),
.A2(n_49),
.B(n_39),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_1),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_60),
.B(n_47),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_31),
.B1(n_39),
.B2(n_34),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_61),
.A2(n_64),
.B1(n_0),
.B2(n_1),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_39),
.B1(n_29),
.B2(n_2),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_63),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_57),
.B1(n_55),
.B2(n_58),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_3),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_2),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_73),
.B(n_7),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_3),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_21),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_81),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_75),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_79),
.B(n_82),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_7),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_69),
.B(n_67),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_86),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_93),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_83),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_71),
.C(n_11),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_85),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_22),
.B(n_16),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_25),
.C(n_17),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_97),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_99),
.A2(n_98),
.B(n_95),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_94),
.C(n_92),
.Y(n_102)
);

INVxp67_ASAP7_75t_SL g103 ( 
.A(n_102),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_101),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_104),
.B(n_89),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_88),
.B(n_97),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_84),
.B1(n_90),
.B2(n_20),
.Y(n_107)
);

A2O1A1O1Ixp25_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_18),
.B(n_24),
.C(n_26),
.D(n_27),
.Y(n_108)
);


endmodule