module fake_jpeg_29293_n_133 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_133);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_9),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_24),
.Y(n_30)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_30),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_32),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_37),
.Y(n_41)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_15),
.B(n_27),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_45),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_27),
.C(n_14),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_32),
.B(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_48),
.B(n_54),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_20),
.B(n_25),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_22),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_SL g51 ( 
.A(n_30),
.B(n_23),
.C(n_25),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_30),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_22),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_58),
.B(n_65),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_50),
.A2(n_33),
.B1(n_39),
.B2(n_40),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_59),
.A2(n_53),
.B1(n_56),
.B2(n_49),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_35),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_33),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_68),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_26),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_66),
.B(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_29),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_44),
.B(n_21),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_29),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_26),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_26),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_39),
.B1(n_46),
.B2(n_42),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_73),
.A2(n_46),
.B1(n_42),
.B2(n_49),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_81),
.B1(n_61),
.B2(n_75),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_38),
.C(n_43),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_69),
.C(n_73),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_17),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_88),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_26),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_62),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_17),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_70),
.B1(n_60),
.B2(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_78),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_91),
.B(n_92),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_83),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_98),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_57),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_97),
.C(n_100),
.Y(n_104)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_84),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_64),
.Y(n_100)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_87),
.C(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_103),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_80),
.C(n_77),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_96),
.C(n_90),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_106),
.B(n_28),
.Y(n_116)
);

A2O1A1O1Ixp25_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_75),
.B(n_28),
.C(n_7),
.D(n_8),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_101),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_111),
.Y(n_121)
);

INVxp67_ASAP7_75t_SL g112 ( 
.A(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_95),
.B(n_96),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_116),
.C(n_107),
.Y(n_119)
);

OA21x2_ASAP7_75t_SL g123 ( 
.A1(n_119),
.A2(n_111),
.B(n_115),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_L g120 ( 
.A1(n_114),
.A2(n_104),
.A3(n_16),
.B1(n_76),
.B2(n_11),
.C1(n_3),
.C2(n_10),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_16),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_110),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_123),
.C(n_124),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_21),
.C(n_5),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

AOI322xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_118),
.A3(n_119),
.B1(n_11),
.B2(n_13),
.C1(n_3),
.C2(n_10),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_129),
.C(n_127),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_13),
.Y(n_133)
);


endmodule