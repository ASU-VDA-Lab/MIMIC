module fake_jpeg_18238_n_90 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_90);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_90;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx10_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_0),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_19),
.A2(n_26),
.B1(n_16),
.B2(n_14),
.Y(n_29)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

INVx5_ASAP7_75t_SL g33 ( 
.A(n_21),
.Y(n_33)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_21),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_20),
.A2(n_16),
.B1(n_14),
.B2(n_17),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_21),
.B1(n_23),
.B2(n_22),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_24),
.C(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_26),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_10),
.B(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_15),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_36),
.B1(n_37),
.B2(n_27),
.Y(n_48)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_51),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_30),
.B1(n_44),
.B2(n_28),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_12),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_10),
.B(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_52),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_56),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_32),
.B1(n_22),
.B2(n_27),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_39),
.B1(n_40),
.B2(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_59),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_24),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_50),
.C(n_52),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_24),
.Y(n_60)
);

OAI21x1_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_46),
.B(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_61),
.B(n_12),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_63),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_46),
.C(n_50),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_58),
.C(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_8),
.Y(n_69)
);

OAI322xp33_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_4),
.A3(n_9),
.B1(n_2),
.B2(n_3),
.C1(n_7),
.C2(n_0),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_73),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_2),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_56),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_79),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_66),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_75),
.C(n_70),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_80),
.A2(n_45),
.B(n_34),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_76),
.B(n_3),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_81),
.A2(n_64),
.B1(n_4),
.B2(n_1),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_83),
.A2(n_73),
.B(n_45),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_84),
.B(n_25),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_85),
.A2(n_86),
.B(n_82),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_87),
.A2(n_88),
.B(n_28),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_30),
.Y(n_90)
);


endmodule