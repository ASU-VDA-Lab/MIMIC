module fake_jpeg_9546_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_38),
.Y(n_66)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_42),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_44),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_0),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_17),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_33),
.B1(n_19),
.B2(n_29),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_24),
.B(n_2),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_30),
.B(n_29),
.C(n_27),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_2),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

CKINVDCx9p33_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_51),
.A2(n_58),
.B1(n_25),
.B2(n_23),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_33),
.B1(n_26),
.B2(n_35),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_56),
.B1(n_59),
.B2(n_63),
.Y(n_82)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_65),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_26),
.B1(n_34),
.B2(n_31),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_18),
.B1(n_29),
.B2(n_27),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_68),
.B1(n_44),
.B2(n_46),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_35),
.B1(n_34),
.B2(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_67),
.Y(n_92)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_39),
.A2(n_31),
.B1(n_30),
.B2(n_24),
.Y(n_68)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_18),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_25),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_48),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_42),
.A2(n_45),
.B1(n_41),
.B2(n_43),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_75),
.A2(n_42),
.B1(n_45),
.B2(n_43),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_70),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_77),
.B(n_83),
.Y(n_116)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_80),
.Y(n_119)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_87),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_85),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_41),
.B1(n_38),
.B2(n_37),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_86),
.A2(n_90),
.B1(n_102),
.B2(n_106),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_88),
.B(n_91),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_89),
.B(n_94),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_38),
.B1(n_37),
.B2(n_45),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_66),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_93),
.A2(n_98),
.B1(n_104),
.B2(n_20),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_69),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_95),
.B(n_97),
.Y(n_142)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_57),
.A2(n_43),
.B1(n_38),
.B2(n_37),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_67),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_99),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_105),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_56),
.A2(n_38),
.B1(n_19),
.B2(n_23),
.Y(n_102)
);

AOI31xp33_ASAP7_75t_L g103 ( 
.A1(n_55),
.A2(n_36),
.A3(n_43),
.B(n_21),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_103),
.A2(n_109),
.B1(n_81),
.B2(n_20),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_55),
.A2(n_44),
.B1(n_30),
.B2(n_19),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_48),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_53),
.A2(n_36),
.B1(n_22),
.B2(n_28),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_15),
.C(n_14),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_25),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_113),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_73),
.B1(n_22),
.B2(n_74),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_59),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_76),
.B(n_23),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_3),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_117),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_139),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_3),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_120),
.A2(n_131),
.B(n_111),
.Y(n_167)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_122),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_73),
.B1(n_53),
.B2(n_20),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_124),
.A2(n_133),
.B1(n_137),
.B2(n_138),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_129),
.B(n_130),
.Y(n_175)
);

MAJx2_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_36),
.C(n_73),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_86),
.A2(n_74),
.B1(n_50),
.B2(n_60),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_93),
.A2(n_60),
.B1(n_50),
.B2(n_22),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_135),
.A2(n_136),
.B1(n_141),
.B2(n_85),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_95),
.A2(n_50),
.B1(n_28),
.B2(n_17),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_81),
.A2(n_28),
.B1(n_17),
.B2(n_36),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_87),
.A2(n_90),
.B1(n_102),
.B2(n_103),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_140),
.B(n_4),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_92),
.A2(n_28),
.B1(n_72),
.B2(n_15),
.Y(n_141)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_144),
.Y(n_159)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_92),
.B(n_72),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_82),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_127),
.A2(n_98),
.B(n_89),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_147),
.A2(n_152),
.B(n_120),
.Y(n_191)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_148),
.B(n_157),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_149),
.B(n_166),
.C(n_138),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_101),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_155),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_91),
.B(n_110),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_151),
.A2(n_154),
.B(n_167),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_142),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_82),
.B1(n_104),
.B2(n_83),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_153),
.A2(n_160),
.B1(n_5),
.B2(n_6),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_79),
.B(n_106),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_3),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_128),
.A2(n_111),
.B1(n_107),
.B2(n_96),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_162),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_163),
.B(n_169),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_4),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_174),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_14),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_107),
.B(n_84),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_168),
.A2(n_137),
.B(n_132),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g170 ( 
.A(n_121),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_170),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_122),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_172),
.Y(n_196)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_125),
.A2(n_80),
.B1(n_78),
.B2(n_85),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_173),
.A2(n_136),
.B1(n_143),
.B2(n_139),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_121),
.B(n_5),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_133),
.B1(n_141),
.B2(n_135),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_13),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_178),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_13),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_5),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_180),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_13),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_181),
.A2(n_156),
.B1(n_157),
.B2(n_179),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_118),
.B(n_130),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_183),
.A2(n_191),
.B(n_201),
.Y(n_224)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_184),
.B(n_186),
.Y(n_221)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_166),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_192),
.A2(n_193),
.B1(n_11),
.B2(n_12),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_160),
.A2(n_130),
.B1(n_134),
.B2(n_144),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_195),
.A2(n_204),
.B1(n_206),
.B2(n_211),
.Y(n_231)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_198),
.B(n_209),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_165),
.B(n_120),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_200),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_155),
.B(n_140),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_5),
.B(n_6),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_172),
.A2(n_132),
.B1(n_117),
.B2(n_7),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_134),
.B1(n_117),
.B2(n_7),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_178),
.B1(n_180),
.B2(n_174),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_175),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_151),
.B(n_8),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_210),
.Y(n_233)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_147),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_150),
.B(n_9),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_167),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_164),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_148),
.B(n_9),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_175),
.C(n_149),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_215),
.C(n_219),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_175),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_218),
.A2(n_238),
.B1(n_199),
.B2(n_202),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_152),
.C(n_153),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_194),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_226),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_152),
.C(n_154),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_227),
.C(n_229),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_225),
.A2(n_236),
.B1(n_241),
.B2(n_200),
.Y(n_247)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_185),
.B(n_152),
.C(n_156),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_164),
.Y(n_230)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_196),
.Y(n_232)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_171),
.C(n_161),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_237),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_198),
.A2(n_161),
.B1(n_164),
.B2(n_169),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_202),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_204),
.A2(n_162),
.B1(n_12),
.B2(n_13),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_183),
.B(n_162),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_11),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_240),
.B(n_203),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_181),
.A2(n_11),
.B1(n_12),
.B2(n_183),
.Y(n_241)
);

MAJx2_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_188),
.C(n_206),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_242),
.B(n_264),
.Y(n_273)
);

AOI22x1_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_195),
.B1(n_193),
.B2(n_205),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_SL g274 ( 
.A1(n_244),
.A2(n_235),
.B(n_224),
.C(n_234),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_214),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_248),
.C(n_256),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_247),
.A2(n_250),
.B1(n_255),
.B2(n_258),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_231),
.A2(n_184),
.B1(n_186),
.B2(n_207),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_252),
.B(n_253),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_221),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_212),
.B1(n_187),
.B2(n_182),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_259),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_222),
.B1(n_239),
.B2(n_232),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_220),
.B(n_208),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_226),
.A2(n_187),
.B1(n_182),
.B2(n_192),
.Y(n_260)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_260),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_219),
.B(n_223),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_262),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_188),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_237),
.A2(n_211),
.B1(n_213),
.B2(n_201),
.Y(n_263)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_263),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_216),
.Y(n_265)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_265),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_276),
.C(n_269),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_260),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_272),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_243),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_279),
.Y(n_285)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_274),
.A2(n_270),
.B1(n_271),
.B2(n_263),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_224),
.C(n_217),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_277),
.A2(n_281),
.B(n_265),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_264),
.B(n_217),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_278),
.B(n_242),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_250),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_247),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_216),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_244),
.A2(n_233),
.B(n_197),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_282),
.A2(n_233),
.B(n_218),
.Y(n_295)
);

BUFx12_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_282),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_289),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_SL g286 ( 
.A(n_276),
.B(n_261),
.C(n_256),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_286),
.A2(n_288),
.B(n_296),
.Y(n_309)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_257),
.B1(n_251),
.B2(n_249),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_281),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_290),
.B(n_291),
.Y(n_304)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_295),
.C(n_297),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_267),
.C(n_271),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_SL g296 ( 
.A(n_274),
.B(n_243),
.C(n_262),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_273),
.B(n_190),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_273),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_301),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_275),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_288),
.B(n_266),
.Y(n_302)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_302),
.Y(n_318)
);

AOI21x1_ASAP7_75t_SL g303 ( 
.A1(n_295),
.A2(n_290),
.B(n_274),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_303),
.A2(n_284),
.B(n_12),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_298),
.B(n_283),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_310),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_311),
.B(n_284),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_292),
.C(n_293),
.Y(n_310)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_312),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_303),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_309),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_307),
.A2(n_270),
.B1(n_274),
.B2(n_278),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_315),
.B(n_299),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_304),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_316),
.B(n_313),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_305),
.A2(n_190),
.B1(n_197),
.B2(n_210),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_317),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_320),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_322),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_318),
.B(n_208),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_326),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_319),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_329),
.B(n_330),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_323),
.A2(n_320),
.B(n_315),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_308),
.C(n_310),
.Y(n_332)
);

NOR2x1_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_331),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_333),
.B(n_325),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_335),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_325),
.B1(n_305),
.B2(n_299),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_300),
.Y(n_338)
);


endmodule