module real_jpeg_16331_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_455;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_458),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_0),
.B(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_1),
.A2(n_67),
.B1(n_131),
.B2(n_135),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_1),
.A2(n_66),
.B1(n_351),
.B2(n_355),
.Y(n_350)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_3),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_3),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_3),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_3),
.Y(n_127)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_4),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_4),
.A2(n_100),
.B1(n_180),
.B2(n_183),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_4),
.A2(n_100),
.B1(n_199),
.B2(n_202),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_4),
.A2(n_100),
.B1(n_251),
.B2(n_253),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_5),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_5),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_5),
.B(n_28),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_5),
.A2(n_80),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_5),
.B(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_5),
.A2(n_80),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_5),
.B(n_139),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_5),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_5),
.B(n_284),
.Y(n_322)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_6),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_6),
.Y(n_208)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_6),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_7),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_7),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_7),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g252 ( 
.A(n_7),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_7),
.Y(n_373)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_8),
.Y(n_92)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_8),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_9),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_11),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_11),
.Y(n_201)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_11),
.Y(n_211)
);

BUFx4f_ASAP7_75t_L g362 ( 
.A(n_11),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_12),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_12),
.A2(n_22),
.B1(n_105),
.B2(n_109),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_12),
.A2(n_22),
.B1(n_358),
.B2(n_363),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_13),
.Y(n_83)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_13),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_161),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_160),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_140),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_19),
.B(n_140),
.Y(n_160)
);

BUFx24_ASAP7_75t_SL g460 ( 
.A(n_19),
.Y(n_460)
);

FAx1_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_60),
.CI(n_95),
.CON(n_19),
.SN(n_19)
);

NAND2xp33_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_21),
.A2(n_35),
.B1(n_130),
.B2(n_139),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_25),
.Y(n_138)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_25),
.Y(n_159)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_30),
.Y(n_257)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

NAND2xp33_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_53),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_34),
.A2(n_53),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_35),
.A2(n_130),
.B1(n_139),
.B2(n_153),
.Y(n_152)
);

AOI22x1_ASAP7_75t_L g178 ( 
.A1(n_35),
.A2(n_139),
.B1(n_153),
.B2(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_35),
.A2(n_139),
.B(n_153),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_53),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_42),
.B1(n_46),
.B2(n_50),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_45),
.Y(n_182)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_47),
.Y(n_261)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_71),
.B1(n_72),
.B2(n_74),
.Y(n_70)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_53),
.Y(n_139)
);

OA22x2_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_55),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g297 ( 
.A(n_55),
.Y(n_297)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_55),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_70),
.B(n_76),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_65),
.A2(n_66),
.B1(n_370),
.B2(n_374),
.Y(n_369)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_68),
.B(n_80),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_94),
.Y(n_93)
);

OAI21x1_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_87),
.B(n_93),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_78),
.B1(n_86),
.B2(n_98),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_70),
.A2(n_78),
.B1(n_86),
.B2(n_98),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_70),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_70),
.B(n_86),
.Y(n_401)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_71),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_71),
.Y(n_230)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_84),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_77),
.B(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_80),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_80),
.B(n_307),
.Y(n_306)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_87),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_103),
.C(n_129),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_97),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_97),
.A2(n_143),
.B1(n_177),
.B2(n_178),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_97),
.B(n_348),
.C(n_391),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_97),
.B(n_247),
.C(n_413),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_97),
.A2(n_143),
.B1(n_187),
.B2(n_248),
.Y(n_423)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_103),
.B(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_103),
.B(n_152),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_111),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_104),
.A2(n_283),
.B1(n_284),
.B2(n_369),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_107),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_109),
.Y(n_253)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_121),
.Y(n_111)
);

NAND2x1p5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_112),
.A2(n_121),
.B(n_171),
.Y(n_170)
);

OA22x2_ASAP7_75t_L g249 ( 
.A1(n_112),
.A2(n_121),
.B1(n_171),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_112),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_112),
.A2(n_368),
.B(n_377),
.Y(n_367)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_115),
.Y(n_320)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_119),
.Y(n_303)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_121),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_126),
.B2(n_128),
.Y(n_122)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_125),
.Y(n_173)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_125),
.Y(n_268)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_146),
.C(n_150),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_141),
.A2(n_142),
.B1(n_146),
.B2(n_147),
.Y(n_443)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_151),
.C(n_152),
.Y(n_150)
);

XOR2x1_ASAP7_75t_SL g167 ( 
.A(n_146),
.B(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_147),
.B(n_382),
.C(n_387),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_147),
.B(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_148),
.A2(n_149),
.B1(n_388),
.B2(n_409),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_148),
.B(n_170),
.C(n_177),
.Y(n_427)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_150),
.B(n_443),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g189 ( 
.A(n_153),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g255 ( 
.A1(n_155),
.A2(n_256),
.A3(n_258),
.B1(n_259),
.B2(n_262),
.Y(n_255)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVxp67_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_440),
.B(n_455),
.Y(n_162)
);

AO221x1_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_344),
.B1(n_433),
.B2(n_438),
.C(n_439),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_275),
.B(n_343),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_240),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_166),
.B(n_240),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_185),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_167),
.B(n_186),
.C(n_218),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_177),
.B2(n_178),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_171),
.Y(n_282)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_177),
.A2(n_178),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_177),
.Y(n_337)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_218),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_186)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_187),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_187),
.B(n_395),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_190),
.A2(n_192),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_190),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_192),
.Y(n_246)
);

NOR2xp67_ASAP7_75t_SL g310 ( 
.A(n_192),
.B(n_311),
.Y(n_310)
);

OA21x2_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_197),
.B(n_205),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_198),
.A2(n_206),
.B1(n_212),
.B2(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_201),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_201),
.Y(n_363)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_205),
.A2(n_350),
.B(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_212),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_206),
.B(n_272),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_206),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g386 ( 
.A(n_208),
.Y(n_386)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_210),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVxp33_ASAP7_75t_L g270 ( 
.A(n_212),
.Y(n_270)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_214),
.Y(n_305)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_234),
.B2(n_235),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_220),
.B(n_234),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_231),
.B2(n_233),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_228),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_234),
.A2(n_235),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_235),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_235),
.B(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_235),
.B(n_322),
.Y(n_323)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_238),
.Y(n_274)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_249),
.C(n_254),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_241),
.A2(n_242),
.B1(n_339),
.B2(n_341),
.Y(n_338)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_247),
.B2(n_248),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NOR2xp67_ASAP7_75t_SL g292 ( 
.A(n_246),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_246),
.B(n_293),
.Y(n_324)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

AOI21x1_ASAP7_75t_L g393 ( 
.A1(n_248),
.A2(n_394),
.B(n_396),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_249),
.B(n_288),
.C(n_289),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_249),
.A2(n_289),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_249),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_249),
.A2(n_254),
.B1(n_330),
.B2(n_340),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_249),
.A2(n_330),
.B1(n_349),
.B2(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_250),
.Y(n_285)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_254),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_269),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_269),
.Y(n_286)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_261),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp67_ASAP7_75t_SL g379 ( 
.A(n_271),
.B(n_357),
.Y(n_379)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_274),
.Y(n_315)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_274),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_334),
.B(n_342),
.Y(n_275)
);

OAI21x1_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_290),
.B(n_333),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_287),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_278),
.B(n_287),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_286),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_280),
.A2(n_281),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_280),
.A2(n_281),
.B1(n_384),
.B2(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp33_ASAP7_75t_R g326 ( 
.A(n_281),
.B(n_295),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_281),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_281),
.B(n_384),
.Y(n_383)
);

AO22x2_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_282),
.B(n_283),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_286),
.B(n_336),
.C(n_337),
.Y(n_335)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_289),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_325),
.B(n_332),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_309),
.B(n_324),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

OAI32xp33_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_298),
.A3(n_302),
.B1(n_304),
.B2(n_306),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_321),
.B(n_323),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_316),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_319),
.Y(n_355)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_320),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_327),
.Y(n_332)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_330),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_338),
.Y(n_334)
);

NOR2x1_ASAP7_75t_L g342 ( 
.A(n_335),
.B(n_338),
.Y(n_342)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_337),
.Y(n_391)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_339),
.Y(n_341)
);

NOR3xp33_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_403),
.C(n_416),
.Y(n_344)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_345),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_389),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_346),
.B(n_389),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_366),
.C(n_381),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_347),
.B(n_366),
.Y(n_415)
);

XNOR2x1_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_365),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_349),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_350),
.A2(n_356),
.B1(n_357),
.B2(n_364),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_367),
.A2(n_378),
.B1(n_379),
.B2(n_380),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_367),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_367),
.B(n_379),
.Y(n_398)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_378),
.A2(n_379),
.B1(n_400),
.B2(n_402),
.Y(n_399)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

AOI21xp33_ASAP7_75t_L g448 ( 
.A1(n_379),
.A2(n_398),
.B(n_400),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_381),
.B(n_415),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

XNOR2x1_ASAP7_75t_L g407 ( 
.A(n_383),
.B(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_384),
.Y(n_425)
);

INVx6_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_388),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_392),
.Y(n_389)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_390),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_397),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_393),
.B(n_397),
.C(n_454),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_396),
.B(n_445),
.C(n_447),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_396),
.B(n_445),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_400),
.Y(n_402)
);

A2O1A1Ixp33_ASAP7_75t_L g433 ( 
.A1(n_403),
.A2(n_434),
.B(n_435),
.C(n_437),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_414),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_404),
.B(n_414),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_410),
.C(n_412),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_406),
.A2(n_407),
.B1(n_410),
.B2(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_410),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_412),
.B(n_419),
.Y(n_418)
);

XNOR2x1_ASAP7_75t_L g422 ( 
.A(n_413),
.B(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_417),
.B(n_428),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_417),
.B(n_436),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_418),
.B(n_421),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_421),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_424),
.C(n_426),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_422),
.B(n_431),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_424),
.A2(n_426),
.B1(n_427),
.B2(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_424),
.Y(n_432)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

NOR2x1_ASAP7_75t_L g436 ( 
.A(n_429),
.B(n_430),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_449),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_441),
.A2(n_456),
.B(n_457),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_444),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_442),
.B(n_444),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_447),
.A2(n_448),
.B1(n_451),
.B2(n_452),
.Y(n_450)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_450),
.B(n_453),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_450),
.B(n_453),
.Y(n_456)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_451),
.Y(n_452)
);


endmodule