module real_aes_1341_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g549 ( .A(n_0), .B(n_189), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_1), .B(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g120 ( .A(n_2), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_3), .B(n_481), .Y(n_480) );
NAND2xp33_ASAP7_75t_SL g535 ( .A(n_4), .B(n_149), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_5), .B(n_129), .Y(n_180) );
INVx1_ASAP7_75t_L g528 ( .A(n_6), .Y(n_528) );
INVx1_ASAP7_75t_L g226 ( .A(n_7), .Y(n_226) );
CKINVDCx16_ASAP7_75t_R g763 ( .A(n_8), .Y(n_763) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_9), .Y(n_240) );
AND2x2_ASAP7_75t_L g478 ( .A(n_10), .B(n_168), .Y(n_478) );
INVx2_ASAP7_75t_L g128 ( .A(n_11), .Y(n_128) );
CKINVDCx16_ASAP7_75t_R g462 ( .A(n_12), .Y(n_462) );
INVx1_ASAP7_75t_L g190 ( .A(n_13), .Y(n_190) );
AOI221x1_ASAP7_75t_L g531 ( .A1(n_14), .A2(n_154), .B1(n_483), .B2(n_532), .C(n_534), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_15), .B(n_481), .Y(n_518) );
INVx1_ASAP7_75t_L g465 ( .A(n_16), .Y(n_465) );
INVx1_ASAP7_75t_L g187 ( .A(n_17), .Y(n_187) );
INVx1_ASAP7_75t_SL g173 ( .A(n_18), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_19), .B(n_140), .Y(n_139) );
AOI33xp33_ASAP7_75t_L g206 ( .A1(n_20), .A2(n_50), .A3(n_117), .B1(n_135), .B2(n_207), .B3(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_21), .A2(n_483), .B(n_484), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_22), .B(n_189), .Y(n_485) );
AOI221xp5_ASAP7_75t_SL g539 ( .A1(n_23), .A2(n_39), .B1(n_481), .B2(n_483), .C(n_540), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_24), .Y(n_101) );
INVx1_ASAP7_75t_L g234 ( .A(n_25), .Y(n_234) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_26), .A2(n_88), .B(n_128), .Y(n_127) );
OR2x2_ASAP7_75t_L g130 ( .A(n_26), .B(n_88), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_27), .B(n_192), .Y(n_522) );
INVxp67_ASAP7_75t_L g530 ( .A(n_28), .Y(n_530) );
AND2x2_ASAP7_75t_L g504 ( .A(n_29), .B(n_167), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_30), .B(n_161), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_31), .A2(n_483), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_32), .B(n_192), .Y(n_541) );
AND2x2_ASAP7_75t_L g123 ( .A(n_33), .B(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g134 ( .A(n_33), .Y(n_134) );
AND2x2_ASAP7_75t_L g149 ( .A(n_33), .B(n_120), .Y(n_149) );
OR2x6_ASAP7_75t_L g463 ( .A(n_34), .B(n_464), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_35), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_36), .B(n_161), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g113 ( .A1(n_37), .A2(n_114), .B1(n_126), .B2(n_129), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_38), .B(n_146), .Y(n_145) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_40), .A2(n_80), .B1(n_132), .B2(n_483), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_41), .B(n_140), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_42), .Y(n_776) );
XOR2xp5_ASAP7_75t_L g104 ( .A(n_43), .B(n_105), .Y(n_104) );
AOI22x1_ASAP7_75t_SL g779 ( .A1(n_43), .A2(n_65), .B1(n_780), .B2(n_781), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_43), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_44), .B(n_189), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_45), .B(n_151), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_46), .B(n_140), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_47), .Y(n_125) );
AND2x2_ASAP7_75t_L g552 ( .A(n_48), .B(n_167), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_49), .B(n_167), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_51), .B(n_140), .Y(n_218) );
INVx1_ASAP7_75t_L g118 ( .A(n_52), .Y(n_118) );
INVx1_ASAP7_75t_L g142 ( .A(n_52), .Y(n_142) );
AND2x2_ASAP7_75t_L g219 ( .A(n_53), .B(n_167), .Y(n_219) );
AOI221xp5_ASAP7_75t_L g224 ( .A1(n_54), .A2(n_72), .B1(n_132), .B2(n_161), .C(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_55), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_56), .B(n_481), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_57), .B(n_126), .Y(n_242) );
AOI21xp5_ASAP7_75t_SL g156 ( .A1(n_58), .A2(n_132), .B(n_157), .Y(n_156) );
AND2x2_ASAP7_75t_L g495 ( .A(n_59), .B(n_167), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_60), .B(n_192), .Y(n_550) );
INVx1_ASAP7_75t_L g183 ( .A(n_61), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_62), .B(n_189), .Y(n_493) );
AND2x2_ASAP7_75t_SL g523 ( .A(n_63), .B(n_168), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_64), .A2(n_483), .B(n_500), .Y(n_499) );
AOI222xp33_ASAP7_75t_L g99 ( .A1(n_65), .A2(n_100), .B1(n_756), .B2(n_767), .C1(n_790), .C2(n_794), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_65), .Y(n_781) );
INVx1_ASAP7_75t_L g217 ( .A(n_66), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_67), .B(n_192), .Y(n_486) );
AND2x2_ASAP7_75t_SL g513 ( .A(n_68), .B(n_151), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_69), .A2(n_132), .B(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g124 ( .A(n_70), .Y(n_124) );
INVx1_ASAP7_75t_L g144 ( .A(n_70), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_71), .B(n_161), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_73), .Y(n_753) );
AND2x2_ASAP7_75t_L g175 ( .A(n_74), .B(n_154), .Y(n_175) );
INVx1_ASAP7_75t_L g184 ( .A(n_75), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_76), .A2(n_132), .B(n_172), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g131 ( .A1(n_77), .A2(n_132), .B(n_138), .C(n_150), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_78), .B(n_481), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_79), .A2(n_83), .B1(n_161), .B2(n_481), .Y(n_511) );
INVx1_ASAP7_75t_L g466 ( .A(n_81), .Y(n_466) );
AND2x2_ASAP7_75t_SL g153 ( .A(n_82), .B(n_154), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_84), .A2(n_132), .B1(n_204), .B2(n_205), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_85), .B(n_189), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_86), .B(n_189), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_87), .A2(n_483), .B(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g158 ( .A(n_89), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_90), .B(n_192), .Y(n_492) );
AND2x2_ASAP7_75t_L g210 ( .A(n_91), .B(n_154), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_92), .A2(n_232), .B(n_233), .C(n_235), .Y(n_231) );
INVxp67_ASAP7_75t_L g533 ( .A(n_93), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_94), .B(n_481), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_95), .B(n_192), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_96), .A2(n_483), .B(n_520), .Y(n_519) );
BUFx2_ASAP7_75t_L g764 ( .A(n_97), .Y(n_764) );
BUFx2_ASAP7_75t_SL g798 ( .A(n_97), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_98), .B(n_140), .Y(n_159) );
OAI21xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_102), .B(n_746), .Y(n_100) );
AOI21xp33_ASAP7_75t_L g746 ( .A1(n_101), .A2(n_747), .B(n_752), .Y(n_746) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OAI22xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_460), .B1(n_467), .B2(n_469), .Y(n_103) );
INVx1_ASAP7_75t_L g751 ( .A(n_104), .Y(n_751) );
INVx1_ASAP7_75t_L g785 ( .A(n_105), .Y(n_785) );
NAND4xp75_ASAP7_75t_L g105 ( .A(n_106), .B(n_311), .C(n_377), .D(n_440), .Y(n_105) );
NOR2x1_ASAP7_75t_L g106 ( .A(n_107), .B(n_274), .Y(n_106) );
OR3x1_ASAP7_75t_L g107 ( .A(n_108), .B(n_244), .C(n_271), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_176), .B(n_199), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_162), .Y(n_110) );
AND2x2_ASAP7_75t_L g374 ( .A(n_111), .B(n_344), .Y(n_374) );
INVx1_ASAP7_75t_L g447 ( .A(n_111), .Y(n_447) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_152), .Y(n_111) );
INVx2_ASAP7_75t_L g198 ( .A(n_112), .Y(n_198) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_112), .Y(n_262) );
AND2x2_ASAP7_75t_L g266 ( .A(n_112), .B(n_179), .Y(n_266) );
AND2x4_ASAP7_75t_L g282 ( .A(n_112), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g286 ( .A(n_112), .Y(n_286) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_131), .Y(n_112) );
NOR3xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_121), .C(n_125), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x4_ASAP7_75t_L g161 ( .A(n_116), .B(n_122), .Y(n_161) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_119), .Y(n_116) );
OR2x6_ASAP7_75t_L g147 ( .A(n_117), .B(n_136), .Y(n_147) );
INVxp33_ASAP7_75t_L g207 ( .A(n_117), .Y(n_207) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g137 ( .A(n_118), .B(n_120), .Y(n_137) );
AND2x4_ASAP7_75t_L g192 ( .A(n_118), .B(n_143), .Y(n_192) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x6_ASAP7_75t_L g483 ( .A(n_123), .B(n_137), .Y(n_483) );
INVx2_ASAP7_75t_L g136 ( .A(n_124), .Y(n_136) );
AND2x6_ASAP7_75t_L g189 ( .A(n_124), .B(n_141), .Y(n_189) );
INVx4_ASAP7_75t_L g154 ( .A(n_126), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_126), .B(n_239), .Y(n_238) );
AOI21x1_ASAP7_75t_L g545 ( .A1(n_126), .A2(n_546), .B(n_552), .Y(n_545) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx4f_ASAP7_75t_L g151 ( .A(n_127), .Y(n_151) );
AND2x4_ASAP7_75t_L g129 ( .A(n_128), .B(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_SL g168 ( .A(n_128), .B(n_130), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_129), .A2(n_156), .B(n_160), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_129), .B(n_148), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_129), .A2(n_480), .B(n_482), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_129), .B(n_528), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_129), .B(n_530), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_129), .B(n_533), .Y(n_532) );
NOR3xp33_ASAP7_75t_L g534 ( .A(n_129), .B(n_185), .C(n_535), .Y(n_534) );
INVxp67_ASAP7_75t_L g241 ( .A(n_132), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_132), .A2(n_161), .B1(n_527), .B2(n_529), .Y(n_526) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_137), .Y(n_132) );
NOR2x1p5_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
INVx1_ASAP7_75t_L g208 ( .A(n_135), .Y(n_208) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_145), .B(n_148), .Y(n_138) );
INVx1_ASAP7_75t_L g185 ( .A(n_140), .Y(n_185) );
AND2x4_ASAP7_75t_L g481 ( .A(n_140), .B(n_149), .Y(n_481) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_L g157 ( .A1(n_147), .A2(n_148), .B(n_158), .C(n_159), .Y(n_157) );
O2A1O1Ixp33_ASAP7_75t_SL g172 ( .A1(n_147), .A2(n_148), .B(n_173), .C(n_174), .Y(n_172) );
OAI22xp5_ASAP7_75t_L g182 ( .A1(n_147), .A2(n_183), .B1(n_184), .B2(n_185), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_147), .A2(n_148), .B(n_217), .C(n_218), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_SL g225 ( .A1(n_147), .A2(n_148), .B(n_226), .C(n_227), .Y(n_225) );
INVxp67_ASAP7_75t_L g232 ( .A(n_147), .Y(n_232) );
INVx1_ASAP7_75t_L g204 ( .A(n_148), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_148), .A2(n_485), .B(n_486), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_148), .A2(n_492), .B(n_493), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_148), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_148), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_148), .A2(n_541), .B(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_148), .A2(n_549), .B(n_550), .Y(n_548) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_149), .Y(n_235) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_150), .A2(n_202), .B(n_210), .Y(n_201) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_150), .A2(n_202), .B(n_210), .Y(n_250) );
AOI21x1_ASAP7_75t_L g509 ( .A1(n_150), .A2(n_510), .B(n_513), .Y(n_509) );
INVx2_ASAP7_75t_SL g150 ( .A(n_151), .Y(n_150) );
OA21x2_ASAP7_75t_L g223 ( .A1(n_151), .A2(n_224), .B(n_228), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_151), .A2(n_518), .B(n_519), .Y(n_517) );
AND2x2_ASAP7_75t_L g177 ( .A(n_152), .B(n_178), .Y(n_177) );
INVx4_ASAP7_75t_L g263 ( .A(n_152), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_152), .B(n_253), .Y(n_267) );
INVx2_ASAP7_75t_L g281 ( .A(n_152), .Y(n_281) );
AND2x4_ASAP7_75t_L g285 ( .A(n_152), .B(n_286), .Y(n_285) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_152), .Y(n_320) );
OR2x2_ASAP7_75t_L g326 ( .A(n_152), .B(n_165), .Y(n_326) );
NOR2x1_ASAP7_75t_SL g355 ( .A(n_152), .B(n_179), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_152), .B(n_429), .Y(n_457) );
OR2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_155), .Y(n_152) );
INVx3_ASAP7_75t_L g212 ( .A(n_154), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_154), .A2(n_212), .B1(n_231), .B2(n_236), .Y(n_230) );
INVx1_ASAP7_75t_L g243 ( .A(n_161), .Y(n_243) );
AND2x2_ASAP7_75t_L g354 ( .A(n_162), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NAND2x1_ASAP7_75t_L g388 ( .A(n_163), .B(n_178), .Y(n_388) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g195 ( .A(n_165), .Y(n_195) );
INVx2_ASAP7_75t_L g254 ( .A(n_165), .Y(n_254) );
AND2x2_ASAP7_75t_L g277 ( .A(n_165), .B(n_179), .Y(n_277) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_165), .Y(n_304) );
INVx1_ASAP7_75t_L g345 ( .A(n_165), .Y(n_345) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_169), .B(n_175), .Y(n_165) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_166), .A2(n_489), .B(n_495), .Y(n_488) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_166), .A2(n_498), .B(n_504), .Y(n_497) );
AO21x2_ASAP7_75t_L g570 ( .A1(n_166), .A2(n_498), .B(n_504), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_167), .Y(n_166) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_167), .A2(n_539), .B(n_543), .Y(n_538) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_177), .B(n_194), .Y(n_176) );
AND2x2_ASAP7_75t_L g357 ( .A(n_177), .B(n_252), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_178), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g424 ( .A(n_178), .Y(n_424) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx3_ASAP7_75t_L g283 ( .A(n_179), .Y(n_283) );
AND2x4_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_186), .B(n_193), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_185), .B(n_234), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B1(n_190), .B2(n_191), .Y(n_186) );
INVxp67_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVxp67_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
OAI211xp5_ASAP7_75t_SL g360 ( .A1(n_194), .A2(n_361), .B(n_365), .C(n_371), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_195), .B(n_196), .Y(n_194) );
AND2x2_ASAP7_75t_SL g276 ( .A(n_196), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_SL g407 ( .A(n_196), .Y(n_407) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g329 ( .A(n_198), .B(n_283), .Y(n_329) );
OR2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_220), .Y(n_199) );
AOI32xp33_ASAP7_75t_L g365 ( .A1(n_200), .A2(n_349), .A3(n_366), .B1(n_367), .B2(n_369), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_201), .B(n_211), .Y(n_200) );
INVx2_ASAP7_75t_L g291 ( .A(n_201), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_201), .B(n_223), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_203), .B(n_209), .Y(n_202) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx3_ASAP7_75t_L g303 ( .A(n_211), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_211), .B(n_229), .Y(n_334) );
AND2x2_ASAP7_75t_L g339 ( .A(n_211), .B(n_340), .Y(n_339) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_211), .Y(n_421) );
AO21x2_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_219), .Y(n_211) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_212), .A2(n_213), .B(n_219), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
OR2x2_ASAP7_75t_L g322 ( .A(n_220), .B(n_323), .Y(n_322) );
INVx3_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g273 ( .A(n_221), .B(n_247), .Y(n_273) );
AND2x2_ASAP7_75t_L g422 ( .A(n_221), .B(n_420), .Y(n_422) );
AND2x4_ASAP7_75t_L g221 ( .A(n_222), .B(n_229), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g259 ( .A(n_223), .Y(n_259) );
AND2x4_ASAP7_75t_L g298 ( .A(n_223), .B(n_299), .Y(n_298) );
INVxp67_ASAP7_75t_L g332 ( .A(n_223), .Y(n_332) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_223), .Y(n_340) );
AND2x2_ASAP7_75t_L g349 ( .A(n_223), .B(n_229), .Y(n_349) );
INVx1_ASAP7_75t_L g433 ( .A(n_223), .Y(n_433) );
INVx2_ASAP7_75t_L g270 ( .A(n_229), .Y(n_270) );
INVx1_ASAP7_75t_L g297 ( .A(n_229), .Y(n_297) );
INVx1_ASAP7_75t_L g364 ( .A(n_229), .Y(n_364) );
OR2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_237), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_241), .B1(n_242), .B2(n_243), .Y(n_237) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
OAI32xp33_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_255), .A3(n_260), .B1(n_264), .B2(n_268), .Y(n_244) );
INVx1_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_246), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_251), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_247), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g348 ( .A(n_247), .B(n_349), .Y(n_348) );
INVxp67_ASAP7_75t_L g373 ( .A(n_247), .Y(n_373) );
AND2x2_ASAP7_75t_L g454 ( .A(n_247), .B(n_296), .Y(n_454) );
AND2x4_ASAP7_75t_L g247 ( .A(n_248), .B(n_250), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g269 ( .A(n_249), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g368 ( .A(n_249), .B(n_291), .Y(n_368) );
NOR2xp67_ASAP7_75t_L g390 ( .A(n_249), .B(n_270), .Y(n_390) );
NOR2x1_ASAP7_75t_L g432 ( .A(n_249), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g299 ( .A(n_250), .Y(n_299) );
INVx1_ASAP7_75t_L g323 ( .A(n_250), .Y(n_323) );
AND2x2_ASAP7_75t_L g338 ( .A(n_250), .B(n_270), .Y(n_338) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g366 ( .A(n_252), .B(n_355), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_252), .B(n_285), .Y(n_436) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_253), .Y(n_405) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_254), .Y(n_387) );
INVxp67_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g288 ( .A(n_257), .B(n_289), .Y(n_288) );
NOR2xp67_ASAP7_75t_L g372 ( .A(n_257), .B(n_373), .Y(n_372) );
NOR2xp67_ASAP7_75t_SL g459 ( .A(n_257), .B(n_397), .Y(n_459) );
INVx3_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g316 ( .A(n_259), .B(n_270), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_260), .B(n_326), .Y(n_384) );
INVx2_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_SL g350 ( .A(n_261), .B(n_277), .Y(n_350) );
AND2x4_ASAP7_75t_SL g261 ( .A(n_262), .B(n_263), .Y(n_261) );
NOR2x1_ASAP7_75t_L g309 ( .A(n_263), .B(n_310), .Y(n_309) );
AND2x4_ASAP7_75t_L g415 ( .A(n_263), .B(n_286), .Y(n_415) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_263), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_264), .B(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
OR2x2_ASAP7_75t_L g386 ( .A(n_265), .B(n_387), .Y(n_386) );
NOR2x1_ASAP7_75t_L g451 ( .A(n_265), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g375 ( .A(n_266), .B(n_320), .Y(n_375) );
INVxp33_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2x1p5_ASAP7_75t_L g289 ( .A(n_269), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g449 ( .A(n_269), .B(n_331), .Y(n_449) );
INVx2_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_292), .Y(n_274) );
OAI21xp33_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_278), .B(n_287), .Y(n_275) );
AND2x2_ASAP7_75t_L g410 ( .A(n_277), .B(n_285), .Y(n_410) );
NAND2xp33_ASAP7_75t_R g278 ( .A(n_279), .B(n_284), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx1_ASAP7_75t_L g452 ( .A(n_281), .Y(n_452) );
INVx4_ASAP7_75t_L g310 ( .A(n_282), .Y(n_310) );
INVx1_ASAP7_75t_L g429 ( .A(n_283), .Y(n_429) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g423 ( .A(n_285), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_SL g427 ( .A(n_285), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_288), .A2(n_353), .B1(n_457), .B2(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x4_ASAP7_75t_L g317 ( .A(n_291), .B(n_303), .Y(n_317) );
AND2x2_ASAP7_75t_L g331 ( .A(n_291), .B(n_332), .Y(n_331) );
A2O1A1Ixp33_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_300), .B(n_305), .C(n_308), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx3_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g379 ( .A(n_295), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx1_ASAP7_75t_L g307 ( .A(n_296), .Y(n_307) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g367 ( .A(n_297), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g376 ( .A(n_297), .B(n_298), .Y(n_376) );
INVx1_ASAP7_75t_L g408 ( .A(n_297), .Y(n_408) );
AND2x4_ASAP7_75t_L g389 ( .A(n_298), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g411 ( .A(n_298), .B(n_302), .Y(n_411) );
AND2x2_ASAP7_75t_L g419 ( .A(n_298), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_L g394 ( .A(n_302), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_302), .B(n_316), .Y(n_396) );
AND2x2_ASAP7_75t_L g399 ( .A(n_302), .B(n_349), .Y(n_399) );
INVx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_303), .B(n_364), .Y(n_413) );
AND2x2_ASAP7_75t_L g341 ( .A(n_304), .B(n_329), .Y(n_341) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g437 ( .A(n_307), .B(n_317), .Y(n_437) );
BUFx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_309), .B(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g321 ( .A(n_310), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_310), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_351), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_335), .Y(n_312) );
OAI222xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_318), .B1(n_322), .B2(n_324), .C1(n_327), .C2(n_330), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_SL g328 ( .A(n_320), .B(n_329), .Y(n_328) );
OR2x6_ASAP7_75t_L g400 ( .A(n_320), .B(n_370), .Y(n_400) );
NAND5xp2_ASAP7_75t_L g403 ( .A(n_320), .B(n_323), .C(n_339), .D(n_404), .E(n_406), .Y(n_403) );
NAND2x1_ASAP7_75t_L g439 ( .A(n_321), .B(n_325), .Y(n_439) );
INVx2_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
NOR2x1_ASAP7_75t_L g369 ( .A(n_326), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_328), .A2(n_419), .B1(n_422), .B2(n_423), .Y(n_418) );
INVx2_ASAP7_75t_L g370 ( .A(n_329), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_329), .B(n_345), .Y(n_382) );
INVx3_ASAP7_75t_L g417 ( .A(n_330), .Y(n_417) );
NAND2x1p5_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
AND2x2_ASAP7_75t_L g362 ( .A(n_331), .B(n_363), .Y(n_362) );
BUFx2_ASAP7_75t_L g395 ( .A(n_331), .Y(n_395) );
INVx2_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g358 ( .A(n_334), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g335 ( .A(n_336), .B(n_347), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_341), .B(n_342), .Y(n_336) );
AND2x4_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g346 ( .A(n_338), .Y(n_346) );
AOI22xp5_ASAP7_75t_L g347 ( .A1(n_341), .A2(n_348), .B1(n_349), .B2(n_350), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_346), .Y(n_342) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_SL g428 ( .A(n_345), .B(n_429), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_360), .Y(n_351) );
AOI21xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_356), .B(n_358), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g397 ( .A(n_368), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_374), .B1(n_375), .B2(n_376), .Y(n_371) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_401), .Y(n_377) );
NOR3xp33_ASAP7_75t_L g378 ( .A(n_379), .B(n_383), .C(n_391), .Y(n_378) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OA21x2_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_385), .B(n_389), .Y(n_383) );
NAND2xp33_ASAP7_75t_SL g385 ( .A(n_386), .B(n_388), .Y(n_385) );
AOI21xp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_398), .B(n_400), .Y(n_391) );
OAI211xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_395), .B(n_396), .C(n_397), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_395), .A2(n_435), .B1(n_437), .B2(n_438), .Y(n_434) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_402), .B(n_425), .Y(n_401) );
NAND4xp25_ASAP7_75t_L g402 ( .A(n_403), .B(n_409), .C(n_416), .D(n_418), .Y(n_402) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g414 ( .A(n_405), .B(n_415), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVx1_ASAP7_75t_L g445 ( .A(n_408), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B1(n_412), .B2(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_414), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OAI21xp5_ASAP7_75t_SL g425 ( .A1(n_426), .A2(n_430), .B(n_434), .Y(n_425) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_455), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_445), .B(n_446), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B1(n_450), .B2(n_453), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OAI22x1_ASAP7_75t_L g747 ( .A1(n_460), .A2(n_748), .B1(n_749), .B2(n_751), .Y(n_747) );
CKINVDCx11_ASAP7_75t_R g460 ( .A(n_461), .Y(n_460) );
AND2x6_ASAP7_75t_SL g461 ( .A(n_462), .B(n_463), .Y(n_461) );
OR2x6_ASAP7_75t_SL g467 ( .A(n_462), .B(n_468), .Y(n_467) );
OR2x2_ASAP7_75t_L g755 ( .A(n_462), .B(n_463), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_462), .B(n_468), .Y(n_766) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_463), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
CKINVDCx11_ASAP7_75t_R g750 ( .A(n_467), .Y(n_750) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_470), .Y(n_748) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_668), .Y(n_470) );
NOR3xp33_ASAP7_75t_SL g471 ( .A(n_472), .B(n_592), .C(n_642), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_572), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_514), .B(n_553), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_505), .Y(n_475) );
INVx1_ASAP7_75t_SL g678 ( .A(n_476), .Y(n_678) );
AOI32xp33_ASAP7_75t_L g709 ( .A1(n_476), .A2(n_691), .A3(n_710), .B1(n_711), .B2(n_712), .Y(n_709) );
AND2x2_ASAP7_75t_L g711 ( .A(n_476), .B(n_568), .Y(n_711) );
AND2x4_ASAP7_75t_SL g476 ( .A(n_477), .B(n_487), .Y(n_476) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_477), .Y(n_506) );
INVx5_ASAP7_75t_L g571 ( .A(n_477), .Y(n_571) );
OR2x2_ASAP7_75t_L g578 ( .A(n_477), .B(n_570), .Y(n_578) );
INVx2_ASAP7_75t_L g583 ( .A(n_477), .Y(n_583) );
AND2x2_ASAP7_75t_L g595 ( .A(n_477), .B(n_488), .Y(n_595) );
AND2x2_ASAP7_75t_L g600 ( .A(n_477), .B(n_496), .Y(n_600) );
OR2x2_ASAP7_75t_L g607 ( .A(n_477), .B(n_508), .Y(n_607) );
AND2x4_ASAP7_75t_L g616 ( .A(n_477), .B(n_497), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_SL g658 ( .A1(n_477), .A2(n_574), .B(n_609), .C(n_647), .Y(n_658) );
OR2x6_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
INVx3_ASAP7_75t_SL g608 ( .A(n_487), .Y(n_608) );
AND2x2_ASAP7_75t_L g654 ( .A(n_487), .B(n_571), .Y(n_654) );
AND2x4_ASAP7_75t_L g487 ( .A(n_488), .B(n_496), .Y(n_487) );
AND2x2_ASAP7_75t_L g507 ( .A(n_488), .B(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g585 ( .A(n_488), .B(n_497), .Y(n_585) );
AND2x2_ASAP7_75t_L g589 ( .A(n_488), .B(n_568), .Y(n_589) );
INVx1_ASAP7_75t_L g615 ( .A(n_488), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_488), .B(n_497), .Y(n_637) );
INVx2_ASAP7_75t_L g641 ( .A(n_488), .Y(n_641) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_488), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_488), .B(n_571), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_494), .Y(n_489) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g652 ( .A(n_497), .B(n_508), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_503), .Y(n_498) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g662 ( .A(n_506), .Y(n_662) );
NAND2xp33_ASAP7_75t_SL g687 ( .A(n_506), .B(n_579), .Y(n_687) );
AND2x2_ASAP7_75t_L g729 ( .A(n_507), .B(n_571), .Y(n_729) );
AND2x2_ASAP7_75t_L g640 ( .A(n_508), .B(n_641), .Y(n_640) );
BUFx2_ASAP7_75t_L g703 ( .A(n_508), .Y(n_703) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_509), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_514), .A2(n_594), .B1(n_696), .B2(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_536), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_515), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_515), .B(n_619), .Y(n_618) );
AND2x4_ASAP7_75t_L g515 ( .A(n_516), .B(n_524), .Y(n_515) );
INVx2_ASAP7_75t_L g559 ( .A(n_516), .Y(n_559) );
OR2x2_ASAP7_75t_L g563 ( .A(n_516), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_516), .B(n_576), .Y(n_581) );
AND2x4_ASAP7_75t_SL g591 ( .A(n_516), .B(n_525), .Y(n_591) );
OR2x2_ASAP7_75t_L g598 ( .A(n_516), .B(n_538), .Y(n_598) );
OR2x2_ASAP7_75t_L g610 ( .A(n_516), .B(n_525), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_516), .B(n_538), .Y(n_624) );
INVx1_ASAP7_75t_L g629 ( .A(n_516), .Y(n_629) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_516), .Y(n_647) );
AND2x2_ASAP7_75t_L g710 ( .A(n_516), .B(n_630), .Y(n_710) );
INVx2_ASAP7_75t_L g714 ( .A(n_516), .Y(n_714) );
OR2x2_ASAP7_75t_L g721 ( .A(n_516), .B(n_611), .Y(n_721) );
OR2x2_ASAP7_75t_L g743 ( .A(n_516), .B(n_744), .Y(n_743) );
OR2x6_ASAP7_75t_L g516 ( .A(n_517), .B(n_523), .Y(n_516) );
AND2x2_ASAP7_75t_L g560 ( .A(n_524), .B(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_524), .B(n_544), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_524), .B(n_620), .Y(n_682) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g579 ( .A(n_525), .Y(n_579) );
AND2x4_ASAP7_75t_L g630 ( .A(n_525), .B(n_631), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_525), .B(n_575), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_525), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_525), .B(n_564), .Y(n_723) );
AND2x4_ASAP7_75t_L g525 ( .A(n_526), .B(n_531), .Y(n_525) );
AND2x2_ASAP7_75t_L g590 ( .A(n_536), .B(n_591), .Y(n_590) );
AO221x1_ASAP7_75t_L g664 ( .A1(n_536), .A2(n_579), .B1(n_610), .B2(n_665), .C(n_666), .Y(n_664) );
OAI322xp33_ASAP7_75t_L g716 ( .A1(n_536), .A2(n_636), .A3(n_717), .B1(n_719), .B2(n_720), .C1(n_721), .C2(n_722), .Y(n_716) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_544), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx3_ASAP7_75t_L g558 ( .A(n_538), .Y(n_558) );
INVx2_ASAP7_75t_L g564 ( .A(n_538), .Y(n_564) );
AND2x2_ASAP7_75t_L g576 ( .A(n_538), .B(n_544), .Y(n_576) );
INVx1_ASAP7_75t_L g621 ( .A(n_538), .Y(n_621) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_538), .Y(n_677) );
INVx1_ASAP7_75t_L g561 ( .A(n_544), .Y(n_561) );
OR2x2_ASAP7_75t_L g611 ( .A(n_544), .B(n_564), .Y(n_611) );
INVx2_ASAP7_75t_L g631 ( .A(n_544), .Y(n_631) );
INVx1_ASAP7_75t_L g684 ( .A(n_544), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_544), .B(n_714), .Y(n_713) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_551), .Y(n_546) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OAI21xp33_ASAP7_75t_SL g554 ( .A1(n_555), .A2(n_562), .B(n_565), .Y(n_554) );
AOI221xp5_ASAP7_75t_L g593 ( .A1(n_555), .A2(n_594), .B1(n_596), .B2(n_600), .C(n_601), .Y(n_593) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_560), .Y(n_556) );
NOR2x1p5_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g680 ( .A(n_559), .Y(n_680) );
INVx1_ASAP7_75t_SL g599 ( .A(n_560), .Y(n_599) );
OAI21xp5_ASAP7_75t_L g704 ( .A1(n_560), .A2(n_705), .B(n_707), .Y(n_704) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_561), .Y(n_604) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_564), .Y(n_667) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
OAI211xp5_ASAP7_75t_L g642 ( .A1(n_567), .A2(n_643), .B(n_648), .C(n_659), .Y(n_642) );
OR2x2_ASAP7_75t_L g732 ( .A(n_567), .B(n_637), .Y(n_732) );
AND2x2_ASAP7_75t_L g734 ( .A(n_567), .B(n_600), .Y(n_734) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g574 ( .A(n_568), .B(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g636 ( .A(n_568), .B(n_637), .Y(n_636) );
AND2x4_ASAP7_75t_L g674 ( .A(n_568), .B(n_641), .Y(n_674) );
OA33x2_ASAP7_75t_L g681 ( .A1(n_568), .A2(n_598), .A3(n_682), .B1(n_683), .B2(n_685), .B3(n_687), .Y(n_681) );
OR2x2_ASAP7_75t_L g692 ( .A(n_568), .B(n_677), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_568), .B(n_616), .Y(n_706) );
AND2x4_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
AND2x2_ASAP7_75t_L g594 ( .A(n_570), .B(n_595), .Y(n_594) );
AOI22xp33_ASAP7_75t_SL g643 ( .A1(n_570), .A2(n_600), .B1(n_644), .B2(n_645), .Y(n_643) );
NAND3xp33_ASAP7_75t_L g683 ( .A(n_571), .B(n_651), .C(n_684), .Y(n_683) );
AOI322xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_577), .A3(n_579), .B1(n_580), .B2(n_582), .C1(n_586), .C2(n_590), .Y(n_572) );
INVx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g679 ( .A(n_575), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_576), .A2(n_591), .B(n_635), .C(n_638), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_577), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
NAND4xp25_ASAP7_75t_SL g698 ( .A(n_578), .B(n_607), .C(n_699), .D(n_701), .Y(n_698) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx2_ASAP7_75t_L g588 ( .A(n_583), .Y(n_588) );
OR2x2_ASAP7_75t_L g633 ( .A(n_583), .B(n_585), .Y(n_633) );
AND2x2_ASAP7_75t_L g702 ( .A(n_584), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
AND2x2_ASAP7_75t_L g707 ( .A(n_588), .B(n_702), .Y(n_707) );
BUFx2_ASAP7_75t_L g700 ( .A(n_589), .Y(n_700) );
INVx1_ASAP7_75t_SL g730 ( .A(n_590), .Y(n_730) );
AND2x4_ASAP7_75t_L g666 ( .A(n_591), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g719 ( .A(n_591), .Y(n_719) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_612), .C(n_634), .Y(n_592) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx1_ASAP7_75t_SL g656 ( .A(n_598), .Y(n_656) );
OAI211xp5_ASAP7_75t_L g724 ( .A1(n_598), .A2(n_725), .B(n_726), .C(n_735), .Y(n_724) );
OR2x2_ASAP7_75t_L g646 ( .A(n_599), .B(n_647), .Y(n_646) );
OAI22xp33_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_605), .B1(n_608), .B2(n_609), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_603), .B(n_686), .Y(n_685) );
INVxp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_606), .B(n_663), .Y(n_745) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g720 ( .A(n_607), .B(n_608), .Y(n_720) );
OR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g665 ( .A(n_611), .Y(n_665) );
AOI222xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_617), .B1(n_622), .B2(n_626), .C1(n_627), .C2(n_632), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_615), .Y(n_626) );
AND2x2_ASAP7_75t_L g673 ( .A(n_616), .B(n_674), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_616), .A2(n_689), .B1(n_694), .B2(n_698), .Y(n_688) );
INVx2_ASAP7_75t_SL g741 ( .A(n_616), .Y(n_741) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVxp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g697 ( .A(n_621), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_621), .B(n_684), .Y(n_744) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx1_ASAP7_75t_L g657 ( .A(n_625), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_627), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g695 ( .A(n_629), .Y(n_695) );
AND2x2_ASAP7_75t_SL g696 ( .A(n_630), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g738 ( .A(n_630), .B(n_667), .Y(n_738) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g663 ( .A(n_637), .Y(n_663) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g742 ( .A(n_640), .Y(n_742) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_641), .Y(n_686) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
O2A1O1Ixp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_653), .B(n_655), .C(n_658), .Y(n_648) );
AND2x2_ASAP7_75t_SL g649 ( .A(n_650), .B(n_652), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g693 ( .A(n_655), .Y(n_693) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_664), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NOR3xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_708), .C(n_724), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_688), .C(n_704), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI221xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_675), .B1(n_678), .B2(n_679), .C(n_681), .Y(n_671) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_690), .B(n_693), .Y(n_689) );
INVx1_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OR2x2_ASAP7_75t_L g717 ( .A(n_703), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g725 ( .A(n_707), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_715), .Y(n_708) );
INVx2_ASAP7_75t_L g731 ( .A(n_710), .Y(n_731) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
OR2x2_ASAP7_75t_L g722 ( .A(n_713), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI221xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_730), .B1(n_731), .B2(n_732), .C(n_733), .Y(n_727) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_739), .B1(n_743), .B2(n_745), .Y(n_736) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_750), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
BUFx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_765), .Y(n_758) );
INVxp67_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NAND2xp5_ASAP7_75t_SL g760 ( .A(n_761), .B(n_764), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
OR2x2_ASAP7_75t_SL g793 ( .A(n_762), .B(n_764), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g795 ( .A1(n_762), .A2(n_796), .B(n_799), .Y(n_795) );
INVx1_ASAP7_75t_SL g777 ( .A(n_765), .Y(n_777) );
BUFx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
BUFx3_ASAP7_75t_L g775 ( .A(n_766), .Y(n_775) );
BUFx2_ASAP7_75t_L g800 ( .A(n_766), .Y(n_800) );
INVxp67_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_778), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_777), .Y(n_769) );
INVxp67_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
AOI21xp5_ASAP7_75t_L g786 ( .A1(n_771), .A2(n_787), .B(n_788), .Y(n_786) );
NOR2xp33_ASAP7_75t_SL g771 ( .A(n_772), .B(n_776), .Y(n_771) );
INVx1_ASAP7_75t_SL g772 ( .A(n_773), .Y(n_772) );
BUFx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_775), .Y(n_774) );
OAI21xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_782), .B(n_786), .Y(n_778) );
CKINVDCx16_ASAP7_75t_R g789 ( .A(n_779), .Y(n_789) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g787 ( .A(n_783), .Y(n_787) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_SL g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_SL g794 ( .A(n_795), .Y(n_794) );
CKINVDCx11_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
CKINVDCx8_ASAP7_75t_R g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
endmodule