module real_aes_7654_n_8 (n_4, n_0, n_3, n_5, n_2, n_7, n_6, n_1, n_8);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_6;
input n_1;
output n_8;
wire n_17;
wire n_28;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_27;
wire n_9;
wire n_23;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_10;
wire n_33;
INVx1_ASAP7_75t_L g28 ( .A(n_0), .Y(n_28) );
AND2x6_ASAP7_75t_L g11 ( .A(n_1), .B(n_12), .Y(n_11) );
HB1xp67_ASAP7_75t_L g32 ( .A(n_1), .Y(n_32) );
CKINVDCx20_ASAP7_75t_R g25 ( .A(n_2), .Y(n_25) );
INVx2_ASAP7_75t_L g16 ( .A(n_3), .Y(n_16) );
INVx1_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
AOI221xp5_ASAP7_75t_L g8 ( .A1(n_5), .A2(n_9), .B1(n_17), .B2(n_21), .C(n_22), .Y(n_8) );
INVx1_ASAP7_75t_L g20 ( .A(n_5), .Y(n_20) );
INVx1_ASAP7_75t_L g19 ( .A(n_6), .Y(n_19) );
INVx1_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_9), .B(n_19), .Y(n_21) );
INVx1_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
NAND2xp5_ASAP7_75t_SL g10 ( .A(n_11), .B(n_13), .Y(n_10) );
HB1xp67_ASAP7_75t_L g33 ( .A(n_12), .Y(n_33) );
NOR2xp33_ASAP7_75t_L g13 ( .A(n_14), .B(n_16), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_15), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_18), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_19), .B(n_20), .Y(n_18) );
INVx1_ASAP7_75t_L g22 ( .A(n_23), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_24), .B(n_29), .Y(n_23) );
NOR2xp33_ASAP7_75t_L g24 ( .A(n_25), .B(n_26), .Y(n_24) );
HB1xp67_ASAP7_75t_L g26 ( .A(n_27), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_28), .Y(n_27) );
CKINVDCx20_ASAP7_75t_R g29 ( .A(n_30), .Y(n_29) );
NAND2xp5_ASAP7_75t_L g30 ( .A(n_31), .B(n_33), .Y(n_30) );
CKINVDCx16_ASAP7_75t_R g31 ( .A(n_32), .Y(n_31) );
endmodule