module fake_jpeg_15367_n_311 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_6),
.B(n_11),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_9),
.B(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_33),
.Y(n_48)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_31),
.B(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_38),
.Y(n_52)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_50),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

HAxp5_ASAP7_75t_SL g46 ( 
.A(n_32),
.B(n_29),
.CON(n_46),
.SN(n_46)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_39),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_32),
.Y(n_58)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_31),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_58),
.B(n_62),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_17),
.B1(n_19),
.B2(n_33),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_59),
.A2(n_16),
.B1(n_54),
.B2(n_18),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_53),
.B(n_32),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_16),
.C(n_27),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_17),
.B1(n_19),
.B2(n_33),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_78),
.B1(n_28),
.B2(n_25),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_31),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_70),
.Y(n_85)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_35),
.B(n_36),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVxp67_ASAP7_75t_SL g97 ( 
.A(n_69),
.Y(n_97)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_74),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_73),
.A2(n_15),
.B1(n_16),
.B2(n_21),
.Y(n_104)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_76),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_43),
.A2(n_19),
.B1(n_17),
.B2(n_25),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_77),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_33),
.B1(n_29),
.B2(n_28),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_39),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_82),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_84),
.A2(n_95),
.B1(n_98),
.B2(n_101),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_33),
.B1(n_38),
.B2(n_42),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_89),
.B1(n_93),
.B2(n_94),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_38),
.B1(n_50),
.B2(n_40),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_38),
.B1(n_40),
.B2(n_34),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_40),
.B1(n_34),
.B2(n_54),
.Y(n_94)
);

AOI22x1_ASAP7_75t_L g95 ( 
.A1(n_68),
.A2(n_40),
.B1(n_34),
.B2(n_54),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_34),
.B1(n_18),
.B2(n_23),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_59),
.A2(n_74),
.B1(n_71),
.B2(n_18),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_15),
.Y(n_103)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_21),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_60),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_106),
.A2(n_95),
.B1(n_100),
.B2(n_82),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_36),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_61),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_67),
.A2(n_36),
.B1(n_35),
.B2(n_30),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_70),
.B1(n_69),
.B2(n_36),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_16),
.Y(n_131)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_64),
.C(n_55),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_131),
.C(n_135),
.Y(n_163)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_120),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_85),
.C(n_100),
.Y(n_140)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_95),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_122),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_132),
.Y(n_142)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_72),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_127),
.Y(n_154)
);

BUFx12_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_83),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_128),
.B(n_134),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_103),
.B(n_27),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_130),
.B(n_24),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_36),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_36),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_132),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_55),
.C(n_36),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_94),
.B1(n_90),
.B2(n_88),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_91),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_91),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_86),
.A2(n_30),
.B1(n_23),
.B2(n_27),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_30),
.B1(n_23),
.B2(n_27),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_140),
.B(n_149),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_120),
.A2(n_86),
.B1(n_89),
.B2(n_84),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_143),
.A2(n_148),
.B1(n_150),
.B2(n_157),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_93),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_144),
.A2(n_152),
.B(n_136),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_146),
.A2(n_155),
.B1(n_161),
.B2(n_169),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_117),
.A2(n_96),
.B1(n_85),
.B2(n_88),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_108),
.B1(n_109),
.B2(n_105),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_159),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_114),
.A2(n_60),
.B(n_16),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_118),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_24),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_119),
.A2(n_27),
.B1(n_22),
.B2(n_24),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_4),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_113),
.B(n_55),
.Y(n_167)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_55),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_0),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_118),
.A2(n_22),
.B1(n_8),
.B2(n_13),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_135),
.A2(n_22),
.B1(n_7),
.B2(n_12),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_170),
.A2(n_9),
.B1(n_8),
.B2(n_7),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_174),
.Y(n_215)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_149),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_131),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_175),
.B(n_184),
.C(n_199),
.Y(n_220)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_153),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_178),
.B(n_179),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_153),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_181),
.Y(n_210)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_138),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_183),
.A2(n_189),
.B(n_196),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_127),
.C(n_122),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_185),
.A2(n_152),
.B(n_144),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_139),
.A2(n_124),
.B1(n_121),
.B2(n_126),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_186),
.A2(n_190),
.B1(n_201),
.B2(n_157),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_193),
.Y(n_211)
);

OA21x2_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_126),
.B(n_60),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_139),
.A2(n_55),
.B1(n_1),
.B2(n_2),
.Y(n_190)
);

NAND3xp33_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_202),
.C(n_1),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_147),
.Y(n_195)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_147),
.B(n_4),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_6),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_198),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_142),
.B(n_8),
.C(n_1),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_0),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_200),
.Y(n_225)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_160),
.Y(n_219)
);

O2A1O1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_203),
.A2(n_213),
.B(n_185),
.C(n_140),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_208),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_193),
.A2(n_144),
.B1(n_148),
.B2(n_141),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_143),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_183),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_172),
.A2(n_159),
.B(n_151),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_142),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_184),
.C(n_194),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_218),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_194),
.A2(n_188),
.B1(n_171),
.B2(n_176),
.Y(n_222)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_223),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_224),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_201),
.Y(n_229)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_172),
.Y(n_232)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_220),
.C(n_213),
.Y(n_252)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_237),
.Y(n_257)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_238),
.A2(n_245),
.B1(n_187),
.B2(n_141),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_187),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_239),
.B(n_241),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_243),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_206),
.B(n_197),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_181),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_242),
.B(n_204),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_215),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_214),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_247),
.C(n_252),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_220),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_228),
.A2(n_218),
.B1(n_211),
.B2(n_216),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_248),
.A2(n_249),
.B1(n_260),
.B2(n_227),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_208),
.B1(n_219),
.B2(n_203),
.Y(n_249)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_254),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_230),
.A2(n_245),
.B1(n_233),
.B2(n_192),
.Y(n_255)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_207),
.C(n_204),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_231),
.Y(n_262)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_230),
.A2(n_233),
.B1(n_227),
.B2(n_244),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_264),
.C(n_266),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_252),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_235),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_271),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_231),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_199),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_269),
.C(n_162),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_239),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_240),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_274),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_257),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_258),
.B(n_209),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_275),
.B(n_196),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_249),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_281),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_266),
.A2(n_261),
.B(n_251),
.Y(n_279)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_248),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_282),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_236),
.C(n_237),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_268),
.A2(n_205),
.B(n_244),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_189),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_284),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_221),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_276),
.A2(n_270),
.B1(n_269),
.B2(n_273),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_289),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_285),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_155),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_277),
.B(n_166),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_293),
.A2(n_295),
.B(n_189),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_192),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_297),
.Y(n_303)
);

AO21x1_ASAP7_75t_L g297 ( 
.A1(n_292),
.A2(n_283),
.B(n_276),
.Y(n_297)
);

AOI322xp5_ASAP7_75t_L g304 ( 
.A1(n_298),
.A2(n_299),
.A3(n_301),
.B1(n_287),
.B2(n_288),
.C1(n_290),
.C2(n_294),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_190),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_301),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_302),
.A2(n_304),
.B(n_300),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_303),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_0),
.B(n_2),
.Y(n_307)
);

OA21x2_ASAP7_75t_SL g308 ( 
.A1(n_307),
.A2(n_3),
.B(n_0),
.Y(n_308)
);

NAND2xp33_ASAP7_75t_R g309 ( 
.A(n_308),
.B(n_2),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_3),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_3),
.B(n_307),
.Y(n_311)
);


endmodule