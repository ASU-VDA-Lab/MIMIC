module real_jpeg_20903_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_244;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_0),
.A2(n_75),
.B1(n_80),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_0),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_0),
.A2(n_46),
.B1(n_47),
.B2(n_153),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_0),
.A2(n_27),
.B1(n_30),
.B2(n_153),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_153),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_1),
.A2(n_75),
.B1(n_80),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_1),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_131),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_131),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_1),
.A2(n_27),
.B1(n_30),
.B2(n_131),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_2),
.A2(n_75),
.B1(n_80),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_2),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_99),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_99),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_99),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_3),
.A2(n_27),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_3),
.A2(n_38),
.B1(n_75),
.B2(n_80),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_3),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_4),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_4),
.B(n_77),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g199 ( 
.A1(n_4),
.A2(n_14),
.B(n_34),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_4),
.A2(n_27),
.B1(n_30),
.B2(n_151),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_4),
.A2(n_60),
.B1(n_61),
.B2(n_208),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_4),
.B(n_182),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_4),
.B(n_46),
.Y(n_232)
);

AOI21xp33_ASAP7_75t_L g236 ( 
.A1(n_4),
.A2(n_46),
.B(n_232),
.Y(n_236)
);

BUFx16f_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_6),
.Y(n_93)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_8),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_8),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_8),
.A2(n_29),
.B1(n_75),
.B2(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_8),
.A2(n_29),
.B1(n_46),
.B2(n_47),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_54),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_9),
.A2(n_27),
.B1(n_30),
.B2(n_54),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_54),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_11),
.A2(n_27),
.B1(n_30),
.B2(n_52),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_52),
.Y(n_159)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_13),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_74),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_32)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_14),
.A2(n_30),
.B(n_32),
.C(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_30),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_15),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_134),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_133),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_108),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_20),
.B(n_108),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_85),
.B2(n_107),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_56),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_42),
.B(n_55),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_24),
.B(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_25),
.A2(n_40),
.B(n_239),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_26),
.Y(n_144)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_27),
.A2(n_30),
.B1(n_44),
.B2(n_50),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_27),
.A2(n_35),
.B(n_151),
.C(n_199),
.Y(n_198)
);

NAND2xp33_ASAP7_75t_SL g233 ( 
.A(n_27),
.B(n_44),
.Y(n_233)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g231 ( 
.A1(n_30),
.A2(n_47),
.A3(n_50),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_31),
.B(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_32),
.A2(n_40),
.B1(n_67),
.B2(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_32),
.A2(n_36),
.B(n_95),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_32),
.A2(n_40),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_32),
.B(n_151),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_32),
.A2(n_40),
.B1(n_203),
.B2(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_32),
.A2(n_40),
.B1(n_223),
.B2(n_239),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_33),
.B(n_212),
.Y(n_211)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_67),
.B(n_68),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_40),
.A2(n_68),
.B(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.Y(n_42)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_43),
.A2(n_49),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_43),
.A2(n_49),
.B1(n_181),
.B2(n_236),
.Y(n_235)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B(n_48),
.C(n_49),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_46),
.Y(n_48)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_46),
.B(n_74),
.Y(n_157)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_47),
.A2(n_76),
.B1(n_150),
.B2(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_49),
.A2(n_51),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_49),
.B(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_49),
.B(n_126),
.Y(n_167)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_49),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_69),
.B2(n_70),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_66),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_71),
.B1(n_83),
.B2(n_84),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_59),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_59),
.A2(n_66),
.B1(n_84),
.B2(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B(n_64),
.Y(n_59)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_60),
.A2(n_61),
.B1(n_121),
.B2(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_60),
.A2(n_88),
.B(n_159),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_60),
.B(n_151),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_61),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_61),
.A2(n_93),
.B1(n_193),
.B2(n_208),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_61),
.A2(n_91),
.B(n_195),
.Y(n_224)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_62),
.B(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_62),
.A2(n_63),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_62),
.A2(n_65),
.B(n_123),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_71),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_78),
.B(n_81),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_98),
.B(n_100),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_72),
.A2(n_98),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_72),
.A2(n_130),
.B1(n_132),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_73),
.A2(n_77),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B(n_76),
.C(n_77),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_75),
.Y(n_76)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

HAxp5_ASAP7_75t_SL g150 ( 
.A(n_75),
.B(n_151),
.CON(n_150),
.SN(n_150)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_77),
.B(n_79),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_77),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_85),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_96),
.C(n_101),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_94),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_87),
.B(n_94),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_93),
.Y(n_123)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_96),
.A2(n_97),
.B1(n_101),
.B2(n_102),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_125),
.B(n_127),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_104),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_104),
.A2(n_180),
.B1(n_182),
.B2(n_183),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.C(n_114),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_112),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_114),
.B(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_124),
.C(n_128),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_115),
.A2(n_116),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_119),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_124),
.A2(n_128),
.B1(n_129),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_124),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_277),
.B(n_282),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_184),
.B(n_262),
.C(n_276),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_169),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_137),
.B(n_169),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_154),
.B2(n_168),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_140),
.B(n_141),
.C(n_168),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.C(n_149),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_147),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_148),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_149),
.B(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_152),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_160),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_155),
.B(n_161),
.C(n_165),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_158),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_164),
.B2(n_165),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.C(n_174),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_170),
.B(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_179),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_178),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_179),
.B(n_249),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_261),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_256),
.B(n_260),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_244),
.B(n_255),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_226),
.B(n_243),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_215),
.B(n_225),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_204),
.B(n_214),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_196),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_198),
.B(n_200),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_209),
.B(n_213),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_207),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_216),
.B(n_217),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_224),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_222),
.C(n_224),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_228),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_234),
.B1(n_241),
.B2(n_242),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_229),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_231),
.Y(n_254)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_234),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_237),
.B1(n_238),
.B2(n_240),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_235),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_240),
.C(n_241),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_245),
.B(n_246),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_251),
.B2(n_252),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_253),
.C(n_254),
.Y(n_257)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_257),
.B(n_258),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_263),
.B(n_264),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_274),
.B2(n_275),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_270),
.C(n_275),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_274),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_278),
.B(n_279),
.Y(n_282)
);


endmodule