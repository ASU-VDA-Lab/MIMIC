module fake_jpeg_29200_n_142 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx5p33_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_30),
.Y(n_44)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_37),
.Y(n_48)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_42),
.Y(n_51)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_30),
.A2(n_21),
.B1(n_16),
.B2(n_27),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_30),
.A2(n_21),
.B1(n_16),
.B2(n_27),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_16),
.B1(n_27),
.B2(n_15),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_13),
.B1(n_24),
.B2(n_15),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_24),
.B1(n_13),
.B2(n_25),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_60),
.B1(n_33),
.B2(n_36),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_31),
.A2(n_22),
.B1(n_18),
.B2(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_51),
.B(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_64),
.Y(n_85)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_44),
.B(n_17),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_68),
.Y(n_95)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVxp67_ASAP7_75t_SL g94 ( 
.A(n_70),
.Y(n_94)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_38),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_54),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_79),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_55),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_77),
.B1(n_29),
.B2(n_47),
.Y(n_82)
);

NOR2xp67_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_54),
.B(n_57),
.Y(n_88)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_60),
.B1(n_57),
.B2(n_61),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_91),
.B1(n_57),
.B2(n_65),
.Y(n_101)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_79),
.B1(n_71),
.B2(n_48),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_59),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_99),
.B(n_100),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_67),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_12),
.B(n_11),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_105),
.B(n_5),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_89),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_84),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_88),
.B(n_93),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_112),
.B(n_105),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_86),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_105),
.C(n_90),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_107),
.C(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_117),
.B(n_121),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

AOI221xp5_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_69),
.B1(n_66),
.B2(n_80),
.C(n_94),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_122),
.B(n_123),
.Y(n_128)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_63),
.C(n_102),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_121),
.C(n_119),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_129),
.C(n_126),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_113),
.C(n_108),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_127),
.A2(n_108),
.B(n_10),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_132),
.Y(n_135)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_133),
.A2(n_134),
.B(n_127),
.C(n_70),
.Y(n_136)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_136),
.A2(n_61),
.B1(n_34),
.B2(n_4),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_135),
.A2(n_8),
.B(n_10),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_5),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_2),
.B1(n_7),
.B2(n_119),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_2),
.Y(n_142)
);


endmodule