module fake_jpeg_16604_n_324 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_23),
.B1(n_26),
.B2(n_32),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_63),
.B1(n_31),
.B2(n_27),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_23),
.B1(n_26),
.B2(n_25),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_46),
.A2(n_53),
.B1(n_29),
.B2(n_30),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_17),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_54),
.Y(n_77)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_24),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_52),
.A2(n_29),
.B1(n_34),
.B2(n_30),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_23),
.B1(n_26),
.B2(n_22),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_17),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_59),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_26),
.B1(n_22),
.B2(n_33),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_57),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_18),
.C(n_34),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_44),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_61),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_33),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_32),
.B1(n_22),
.B2(n_33),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_32),
.Y(n_69)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_42),
.B1(n_36),
.B2(n_24),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_70),
.A2(n_78),
.B1(n_90),
.B2(n_91),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_SL g71 ( 
.A1(n_60),
.A2(n_36),
.B(n_42),
.C(n_44),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_71),
.A2(n_65),
.B(n_64),
.C(n_47),
.Y(n_111)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_75),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_52),
.B(n_59),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_31),
.B1(n_27),
.B2(n_34),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_87),
.Y(n_120)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_82),
.A2(n_84),
.B1(n_85),
.B2(n_20),
.Y(n_122)
);

HAxp5_ASAP7_75t_SL g87 ( 
.A(n_52),
.B(n_34),
.CON(n_87),
.SN(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_18),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_68),
.Y(n_102)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_58),
.A2(n_46),
.B1(n_55),
.B2(n_49),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_56),
.A2(n_29),
.B1(n_1),
.B2(n_2),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_20),
.Y(n_117)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_56),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_95),
.B(n_49),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_71),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_101),
.Y(n_135)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_75),
.B(n_61),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_99),
.B(n_86),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_102),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_93),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_90),
.A2(n_65),
.B1(n_64),
.B2(n_47),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_103),
.A2(n_111),
.B1(n_112),
.B2(n_116),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_83),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_110),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_80),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_80),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_90),
.A2(n_65),
.B1(n_64),
.B2(n_47),
.Y(n_112)
);

OR2x2_ASAP7_75t_SL g113 ( 
.A(n_79),
.B(n_29),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_78),
.Y(n_115)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_82),
.A2(n_62),
.B1(n_34),
.B2(n_20),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_122),
.B1(n_91),
.B2(n_94),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_88),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_121),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_74),
.B(n_62),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_68),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_119),
.C(n_102),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_134),
.C(n_137),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_151),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_73),
.B1(n_71),
.B2(n_85),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_146),
.B1(n_150),
.B2(n_152),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_132),
.B(n_109),
.Y(n_156)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_73),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_142),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_107),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_143),
.B(n_145),
.Y(n_155)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_101),
.A2(n_71),
.B1(n_85),
.B2(n_86),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_114),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_148),
.B(n_149),
.Y(n_162)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_95),
.B1(n_84),
.B2(n_76),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_115),
.A2(n_93),
.B1(n_70),
.B2(n_76),
.Y(n_152)
);

AND2x6_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_96),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_154),
.A2(n_165),
.B(n_179),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_156),
.B(n_168),
.Y(n_209)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_110),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_171),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_104),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_167),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_130),
.A2(n_108),
.B1(n_103),
.B2(n_112),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_163),
.A2(n_176),
.B1(n_139),
.B2(n_124),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_126),
.A2(n_117),
.B(n_99),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_103),
.Y(n_166)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_104),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_147),
.B(n_77),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_112),
.Y(n_171)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_181),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_126),
.A2(n_117),
.B(n_111),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_173),
.A2(n_141),
.B(n_133),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_150),
.A2(n_111),
.B1(n_116),
.B2(n_106),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_116),
.C(n_113),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_131),
.C(n_133),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_135),
.A2(n_97),
.B(n_113),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_146),
.A2(n_72),
.B1(n_89),
.B2(n_118),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_180),
.A2(n_124),
.B1(n_129),
.B2(n_131),
.Y(n_188)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

AND2x6_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_151),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_182),
.A2(n_28),
.B(n_21),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_77),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_186),
.A2(n_210),
.B(n_175),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_188),
.A2(n_192),
.B1(n_195),
.B2(n_196),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_199),
.C(n_200),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_155),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_191),
.B(n_201),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_SL g193 ( 
.A1(n_165),
.A2(n_139),
.B(n_152),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_193),
.A2(n_176),
.B1(n_163),
.B2(n_154),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_160),
.A2(n_118),
.B1(n_72),
.B2(n_140),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_157),
.A2(n_118),
.B1(n_92),
.B2(n_2),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_92),
.C(n_28),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_28),
.C(n_21),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_162),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_180),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_160),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_207),
.B1(n_178),
.B2(n_5),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_21),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_153),
.C(n_178),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_0),
.Y(n_206)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_157),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_156),
.B(n_3),
.Y(n_208)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_179),
.A2(n_173),
.B(n_159),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_220),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_194),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_221),
.Y(n_246)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_189),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_181),
.Y(n_217)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_223),
.C(n_234),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_205),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_182),
.C(n_171),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_224),
.B(n_232),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_159),
.Y(n_225)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_226),
.B(n_210),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_184),
.B(n_175),
.Y(n_227)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_187),
.A2(n_170),
.B1(n_174),
.B2(n_172),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_228),
.A2(n_195),
.B1(n_192),
.B2(n_188),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_170),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_230),
.B(n_229),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_174),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_231),
.A2(n_198),
.B(n_206),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_233),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_158),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_169),
.C(n_30),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_200),
.C(n_185),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_201),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_236),
.A2(n_208),
.B1(n_207),
.B2(n_11),
.Y(n_240)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_240),
.A2(n_252),
.B1(n_256),
.B2(n_236),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_245),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_250),
.C(n_257),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_223),
.C(n_234),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_251),
.B(n_225),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_185),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_251),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_231),
.A2(n_202),
.B1(n_186),
.B2(n_203),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_211),
.B(n_209),
.C(n_196),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_246),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_258),
.B(n_241),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_218),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_262),
.C(n_270),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_220),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_248),
.A2(n_212),
.B(n_215),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_240),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_255),
.A2(n_228),
.B(n_231),
.Y(n_264)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_267),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_235),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_252),
.Y(n_279)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_269),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_222),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_222),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_272),
.C(n_274),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_224),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_219),
.C(n_209),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_254),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_276),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_287),
.C(n_272),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_274),
.B(n_253),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_281),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_242),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_273),
.B(n_244),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_284),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_288),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_247),
.C(n_238),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_291),
.C(n_295),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_261),
.C(n_259),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_266),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_237),
.Y(n_296)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_296),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_277),
.A2(n_271),
.B1(n_270),
.B2(n_267),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_283),
.Y(n_302)
);

NOR2xp67_ASAP7_75t_SL g298 ( 
.A(n_283),
.B(n_10),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_10),
.A3(n_16),
.B1(n_15),
.B2(n_14),
.C1(n_12),
.C2(n_4),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_30),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_285),
.Y(n_301)
);

NOR2x1_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_9),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_300),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_303),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_304),
.Y(n_311)
);

A2O1A1Ixp33_ASAP7_75t_L g304 ( 
.A1(n_300),
.A2(n_278),
.B(n_12),
.C(n_6),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_292),
.A2(n_12),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_4),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_308),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_293),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_8),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_291),
.C(n_289),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_313),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_307),
.A2(n_290),
.B(n_294),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_304),
.A2(n_295),
.B1(n_5),
.B2(n_7),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_316),
.Y(n_320)
);

NAND2xp33_ASAP7_75t_SL g318 ( 
.A(n_311),
.B(n_4),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_319),
.Y(n_321)
);

AOI21x1_ASAP7_75t_L g319 ( 
.A1(n_310),
.A2(n_7),
.B(n_8),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_317),
.B(n_320),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_315),
.C(n_316),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_8),
.Y(n_324)
);


endmodule