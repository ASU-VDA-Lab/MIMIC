module fake_jpeg_25975_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx14_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_25),
.Y(n_40)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_10),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_9),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_12),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_25),
.A2(n_22),
.B1(n_16),
.B2(n_21),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_32),
.A2(n_37),
.B1(n_20),
.B2(n_29),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_21),
.B(n_13),
.C(n_15),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_20),
.B(n_14),
.C(n_29),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_23),
.A2(n_22),
.B1(n_19),
.B2(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_15),
.Y(n_46)
);

O2A1O1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_23),
.B(n_27),
.C(n_24),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_36),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_28),
.C(n_27),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_43),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_19),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_50),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_46),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_18),
.B1(n_20),
.B2(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_51),
.B1(n_39),
.B2(n_1),
.Y(n_58)
);

NOR3xp33_ASAP7_75t_SL g53 ( 
.A(n_48),
.B(n_20),
.C(n_29),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_49),
.Y(n_64)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

NOR3xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_57),
.C(n_49),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_0),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_43),
.B(n_45),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_58),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_35),
.B1(n_1),
.B2(n_2),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_62),
.A2(n_52),
.B1(n_44),
.B2(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_0),
.Y(n_73)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_71),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_46),
.B(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_68),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_70),
.A2(n_73),
.B(n_60),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_0),
.Y(n_74)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_8),
.Y(n_79)
);

NOR3xp33_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_8),
.C(n_2),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_57),
.B1(n_63),
.B2(n_55),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_74),
.C(n_71),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_81),
.C(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_77),
.Y(n_89)
);

AO21x2_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_69),
.B(n_61),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_88),
.A2(n_69),
.B1(n_67),
.B2(n_55),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_80),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_91),
.B(n_93),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_92),
.B(n_84),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_81),
.B(n_3),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

AOI322xp5_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_88),
.A3(n_87),
.B1(n_86),
.B2(n_61),
.C1(n_6),
.C2(n_5),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_97),
.B(n_1),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_88),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_95),
.B(n_4),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_98),
.C(n_4),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_102),
.Y(n_104)
);


endmodule