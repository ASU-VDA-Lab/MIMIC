module fake_netlist_5_37_n_47 (n_8, n_10, n_4, n_5, n_7, n_0, n_9, n_2, n_3, n_11, n_6, n_1, n_47);

input n_8;
input n_10;
input n_4;
input n_5;
input n_7;
input n_0;
input n_9;
input n_2;
input n_3;
input n_11;
input n_6;
input n_1;

output n_47;

wire n_29;
wire n_16;
wire n_43;
wire n_12;
wire n_36;
wire n_25;
wire n_18;
wire n_27;
wire n_42;
wire n_22;
wire n_45;
wire n_24;
wire n_28;
wire n_46;
wire n_21;
wire n_44;
wire n_40;
wire n_34;
wire n_38;
wire n_32;
wire n_35;
wire n_41;
wire n_17;
wire n_19;
wire n_37;
wire n_26;
wire n_15;
wire n_30;
wire n_20;
wire n_33;
wire n_14;
wire n_31;
wire n_23;
wire n_13;
wire n_39;

AND2x4_ASAP7_75t_L g12 ( 
.A(n_11),
.B(n_9),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

OAI21x1_ASAP7_75t_L g17 ( 
.A1(n_6),
.A2(n_1),
.B(n_7),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

AND2x6_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

AND2x4_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_4),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_4),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_15),
.B(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_16),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_18),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_24),
.B(n_22),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NOR3xp33_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_19),
.C(n_15),
.Y(n_30)
);

AOI21x1_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_12),
.B(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

OAI21x1_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_26),
.B(n_20),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

OAI222xp33_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_32),
.B1(n_31),
.B2(n_33),
.C1(n_12),
.C2(n_19),
.Y(n_37)
);

NOR3xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_32),
.C(n_31),
.Y(n_38)
);

AOI21xp33_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_35),
.B(n_34),
.Y(n_39)
);

NAND3xp33_ASAP7_75t_SL g40 ( 
.A(n_39),
.B(n_20),
.C(n_14),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_14),
.B1(n_16),
.B2(n_20),
.Y(n_41)
);

NOR3xp33_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_20),
.C(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

NAND3xp33_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_44),
.C(n_16),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_16),
.Y(n_47)
);


endmodule