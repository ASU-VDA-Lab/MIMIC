module fake_netlist_1_11434_n_655 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_655);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_655;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_490;
wire n_247;
wire n_393;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_446;
wire n_342;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_582;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_49), .Y(n_86) );
INVxp33_ASAP7_75t_L g87 ( .A(n_65), .Y(n_87) );
INVxp67_ASAP7_75t_L g88 ( .A(n_59), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_58), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_7), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_84), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_24), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_2), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_70), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_2), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_66), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_25), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_19), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_42), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_53), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_85), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_5), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_71), .Y(n_103) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_45), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_27), .Y(n_105) );
BUFx3_ASAP7_75t_L g106 ( .A(n_23), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_43), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_56), .Y(n_108) );
BUFx2_ASAP7_75t_L g109 ( .A(n_21), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_54), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_22), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_69), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_64), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_26), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_20), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_28), .Y(n_116) );
BUFx10_ASAP7_75t_L g117 ( .A(n_17), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_73), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_16), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_78), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_44), .Y(n_121) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_68), .B(n_83), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_62), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_36), .Y(n_124) );
INVx5_ASAP7_75t_L g125 ( .A(n_104), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_90), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_94), .Y(n_127) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_119), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_92), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_104), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_119), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_86), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_109), .B(n_4), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_92), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_106), .B(n_6), .Y(n_135) );
OAI21x1_ASAP7_75t_L g136 ( .A1(n_100), .A2(n_40), .B(n_81), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_104), .Y(n_137) );
AOI22xp5_ASAP7_75t_L g138 ( .A1(n_86), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_138) );
OAI22xp5_ASAP7_75t_SL g139 ( .A1(n_89), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_139) );
BUFx8_ASAP7_75t_L g140 ( .A(n_100), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_104), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_93), .B(n_10), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_95), .B(n_11), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_108), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_97), .Y(n_145) );
OA21x2_ASAP7_75t_L g146 ( .A1(n_108), .A2(n_46), .B(n_80), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_106), .B(n_11), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_117), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_123), .Y(n_149) );
AOI22xp5_ASAP7_75t_L g150 ( .A1(n_89), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_114), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_98), .B(n_12), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_114), .B(n_13), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_130), .Y(n_154) );
BUFx3_ASAP7_75t_L g155 ( .A(n_135), .Y(n_155) );
BUFx10_ASAP7_75t_L g156 ( .A(n_135), .Y(n_156) );
OR2x2_ASAP7_75t_L g157 ( .A(n_148), .B(n_102), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_130), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_148), .B(n_87), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_130), .Y(n_160) );
INVx5_ASAP7_75t_L g161 ( .A(n_125), .Y(n_161) );
NAND3xp33_ASAP7_75t_L g162 ( .A(n_127), .B(n_124), .C(n_99), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_148), .B(n_112), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_127), .B(n_88), .Y(n_164) );
INVx5_ASAP7_75t_L g165 ( .A(n_125), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_133), .B(n_117), .Y(n_166) );
AOI22xp33_ASAP7_75t_L g167 ( .A1(n_153), .A2(n_117), .B1(n_105), .B2(n_121), .Y(n_167) );
INVx4_ASAP7_75t_L g168 ( .A(n_135), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_153), .Y(n_169) );
XNOR2x2_ASAP7_75t_SL g170 ( .A(n_132), .B(n_113), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_153), .Y(n_171) );
INVx6_ASAP7_75t_L g172 ( .A(n_140), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_130), .Y(n_173) );
BUFx4f_ASAP7_75t_L g174 ( .A(n_147), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_129), .Y(n_175) );
AOI22xp33_ASAP7_75t_L g176 ( .A1(n_133), .A2(n_103), .B1(n_110), .B2(n_120), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_145), .B(n_112), .Y(n_177) );
AND2x6_ASAP7_75t_L g178 ( .A(n_147), .B(n_101), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_145), .B(n_107), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_130), .Y(n_180) );
OAI22xp5_ASAP7_75t_SL g181 ( .A1(n_139), .A2(n_113), .B1(n_96), .B2(n_115), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_137), .Y(n_182) );
INVx1_ASAP7_75t_SL g183 ( .A(n_133), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_129), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_134), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_137), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_147), .A2(n_116), .B1(n_118), .B2(n_107), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_134), .Y(n_188) );
INVxp67_ASAP7_75t_SL g189 ( .A(n_140), .Y(n_189) );
INVx2_ASAP7_75t_SL g190 ( .A(n_157), .Y(n_190) );
NOR2x1_ASAP7_75t_L g191 ( .A(n_162), .B(n_142), .Y(n_191) );
NOR2x1p5_ASAP7_75t_L g192 ( .A(n_189), .B(n_126), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_175), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_166), .B(n_126), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_166), .A2(n_183), .B1(n_178), .B2(n_167), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_175), .Y(n_196) );
INVxp67_ASAP7_75t_SL g197 ( .A(n_155), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_163), .B(n_140), .Y(n_198) );
INVx1_ASAP7_75t_SL g199 ( .A(n_157), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_177), .B(n_179), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_178), .A2(n_132), .B1(n_96), .B2(n_115), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_174), .B(n_136), .Y(n_202) );
INVxp67_ASAP7_75t_SL g203 ( .A(n_155), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_159), .B(n_126), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_169), .A2(n_144), .B1(n_151), .B2(n_143), .Y(n_205) );
BUFx6f_ASAP7_75t_SL g206 ( .A(n_178), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_168), .B(n_131), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_164), .B(n_152), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_172), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_184), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_184), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_176), .B(n_111), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_187), .B(n_111), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_168), .B(n_118), .Y(n_214) );
AO22x1_ASAP7_75t_L g215 ( .A1(n_178), .A2(n_150), .B1(n_138), .B2(n_128), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_178), .A2(n_128), .B1(n_131), .B2(n_151), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_168), .B(n_91), .Y(n_217) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_169), .A2(n_144), .B1(n_146), .B2(n_136), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_185), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_185), .Y(n_220) );
INVx4_ASAP7_75t_L g221 ( .A(n_172), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_178), .A2(n_146), .B1(n_122), .B2(n_123), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_188), .Y(n_223) );
BUFx3_ASAP7_75t_L g224 ( .A(n_172), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_168), .B(n_146), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_171), .B(n_146), .Y(n_226) );
OAI221xp5_ASAP7_75t_L g227 ( .A1(n_171), .A2(n_123), .B1(n_125), .B2(n_137), .C(n_141), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_178), .A2(n_123), .B1(n_125), .B2(n_137), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_172), .B(n_125), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_174), .B(n_155), .Y(n_230) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_174), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_156), .B(n_141), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_156), .B(n_141), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_156), .B(n_141), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_156), .B(n_141), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_204), .A2(n_162), .B(n_188), .C(n_137), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_225), .A2(n_180), .B(n_160), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_226), .A2(n_180), .B(n_160), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_226), .A2(n_186), .B(n_182), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_199), .B(n_14), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_223), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_190), .B(n_181), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_193), .Y(n_243) );
NOR2xp33_ASAP7_75t_SL g244 ( .A(n_206), .B(n_181), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_192), .Y(n_245) );
INVxp67_ASAP7_75t_SL g246 ( .A(n_209), .Y(n_246) );
OAI21x1_ASAP7_75t_L g247 ( .A1(n_202), .A2(n_186), .B(n_182), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_221), .B(n_165), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_207), .B(n_15), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_204), .B(n_15), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_207), .B(n_16), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_202), .A2(n_186), .B(n_182), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_196), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_194), .B(n_17), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_194), .B(n_18), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_216), .A2(n_149), .B1(n_170), .B2(n_165), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_210), .Y(n_257) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_231), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_221), .B(n_165), .Y(n_259) );
INVx3_ASAP7_75t_L g260 ( .A(n_206), .Y(n_260) );
BUFx2_ASAP7_75t_L g261 ( .A(n_209), .Y(n_261) );
NAND2xp33_ASAP7_75t_SL g262 ( .A(n_200), .B(n_149), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_233), .A2(n_154), .B(n_158), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_224), .B(n_165), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_201), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_195), .A2(n_149), .B1(n_154), .B2(n_161), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_234), .A2(n_154), .B(n_158), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_205), .A2(n_149), .B1(n_165), .B2(n_161), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_213), .B(n_18), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_205), .A2(n_149), .B1(n_165), .B2(n_161), .Y(n_270) );
BUFx3_ASAP7_75t_L g271 ( .A(n_224), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_230), .A2(n_161), .B1(n_173), .B2(n_158), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_L g273 ( .A1(n_208), .A2(n_161), .B(n_30), .C(n_31), .Y(n_273) );
OAI21x1_ASAP7_75t_L g274 ( .A1(n_218), .A2(n_173), .B(n_158), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_230), .B(n_29), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_212), .B(n_161), .Y(n_276) );
BUFx2_ASAP7_75t_L g277 ( .A(n_197), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g278 ( .A1(n_198), .A2(n_173), .B(n_158), .C(n_34), .Y(n_278) );
O2A1O1Ixp33_ASAP7_75t_L g279 ( .A1(n_211), .A2(n_32), .B(n_33), .C(n_35), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_219), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_243), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_240), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_245), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_242), .B(n_215), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_258), .B(n_198), .Y(n_285) );
OAI21xp5_ASAP7_75t_L g286 ( .A1(n_236), .A2(n_222), .B(n_238), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_260), .B(n_203), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_239), .A2(n_235), .B(n_232), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_260), .B(n_220), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_256), .B(n_214), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g291 ( .A1(n_249), .A2(n_191), .B1(n_217), .B2(n_218), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_240), .B(n_228), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_277), .B(n_232), .Y(n_293) );
INVxp67_ASAP7_75t_L g294 ( .A(n_251), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_277), .A2(n_227), .B1(n_235), .B2(n_229), .Y(n_295) );
OAI22xp33_ASAP7_75t_L g296 ( .A1(n_265), .A2(n_173), .B1(n_38), .B2(n_39), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_243), .A2(n_173), .B1(n_41), .B2(n_47), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_L g298 ( .A1(n_269), .A2(n_37), .B(n_48), .C(n_50), .Y(n_298) );
CKINVDCx20_ASAP7_75t_R g299 ( .A(n_265), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_254), .Y(n_300) );
AO21x2_ASAP7_75t_L g301 ( .A1(n_274), .A2(n_51), .B(n_52), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_237), .A2(n_55), .B(n_57), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_253), .Y(n_303) );
INVx5_ASAP7_75t_L g304 ( .A(n_260), .Y(n_304) );
OAI22xp5_ASAP7_75t_SL g305 ( .A1(n_244), .A2(n_60), .B1(n_61), .B2(n_63), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_244), .B(n_67), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_275), .B(n_82), .Y(n_307) );
NAND3xp33_ASAP7_75t_L g308 ( .A(n_262), .B(n_72), .C(n_74), .Y(n_308) );
O2A1O1Ixp33_ASAP7_75t_L g309 ( .A1(n_250), .A2(n_75), .B(n_76), .C(n_77), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_253), .B(n_79), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_255), .Y(n_311) );
AOI31xp67_ASAP7_75t_L g312 ( .A1(n_257), .A2(n_280), .A3(n_241), .B(n_275), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_257), .B(n_280), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_SL g314 ( .A1(n_278), .A2(n_279), .B(n_273), .C(n_266), .Y(n_314) );
INVxp67_ASAP7_75t_L g315 ( .A(n_275), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_284), .B(n_241), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_284), .B(n_261), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_294), .B(n_261), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_315), .A2(n_266), .B1(n_246), .B2(n_271), .Y(n_319) );
OA21x2_ASAP7_75t_L g320 ( .A1(n_286), .A2(n_274), .B(n_247), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_313), .Y(n_321) );
OAI21xp5_ASAP7_75t_L g322 ( .A1(n_291), .A2(n_276), .B(n_270), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_314), .A2(n_262), .B(n_252), .Y(n_323) );
AO21x2_ASAP7_75t_L g324 ( .A1(n_301), .A2(n_247), .B(n_268), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_281), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_303), .Y(n_326) );
INVx1_ASAP7_75t_SL g327 ( .A(n_307), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_290), .B(n_271), .Y(n_328) );
OAI21x1_ASAP7_75t_L g329 ( .A1(n_302), .A2(n_263), .B(n_267), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_293), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_285), .B(n_264), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_312), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_285), .B(n_248), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_314), .A2(n_272), .B(n_259), .Y(n_334) );
INVx5_ASAP7_75t_L g335 ( .A(n_307), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_289), .Y(n_336) );
OA21x2_ASAP7_75t_L g337 ( .A1(n_291), .A2(n_298), .B(n_288), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_282), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_300), .B(n_311), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_310), .A2(n_296), .B(n_301), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_289), .B(n_287), .Y(n_341) );
A2O1A1Ixp33_ASAP7_75t_L g342 ( .A1(n_306), .A2(n_309), .B(n_292), .C(n_287), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_304), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_339), .B(n_299), .Y(n_344) );
NOR2x1_ASAP7_75t_SL g345 ( .A(n_335), .B(n_304), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_336), .Y(n_346) );
BUFx5_ASAP7_75t_L g347 ( .A(n_321), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_336), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_321), .B(n_306), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_330), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_330), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_325), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_325), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_332), .Y(n_354) );
AO21x2_ASAP7_75t_L g355 ( .A1(n_340), .A2(n_296), .B(n_308), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_325), .B(n_304), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_335), .B(n_304), .Y(n_357) );
INVxp67_ASAP7_75t_L g358 ( .A(n_318), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_332), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_326), .Y(n_360) );
OA21x2_ASAP7_75t_L g361 ( .A1(n_323), .A2(n_297), .B(n_295), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_320), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_320), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_326), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_326), .B(n_297), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_335), .A2(n_283), .B1(n_305), .B2(n_327), .Y(n_366) );
BUFx2_ASAP7_75t_L g367 ( .A(n_335), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_320), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_320), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_338), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_338), .B(n_316), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_354), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_352), .B(n_335), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_354), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_352), .B(n_353), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_347), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_354), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_353), .B(n_335), .Y(n_378) );
BUFx2_ASAP7_75t_L g379 ( .A(n_347), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_360), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_359), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_359), .Y(n_382) );
INVx3_ASAP7_75t_L g383 ( .A(n_347), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_350), .B(n_328), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_359), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_350), .B(n_328), .Y(n_386) );
AOI22xp33_ASAP7_75t_SL g387 ( .A1(n_347), .A2(n_327), .B1(n_317), .B2(n_319), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_362), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_360), .B(n_316), .Y(n_389) );
BUFx2_ASAP7_75t_L g390 ( .A(n_347), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_364), .B(n_337), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_364), .B(n_337), .Y(n_392) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_361), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_362), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_362), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_370), .B(n_337), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_370), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_363), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_351), .B(n_343), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_371), .B(n_337), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_363), .B(n_343), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_363), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_351), .Y(n_403) );
INVx2_ASAP7_75t_SL g404 ( .A(n_347), .Y(n_404) );
INVx2_ASAP7_75t_SL g405 ( .A(n_347), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_356), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_368), .B(n_324), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_368), .B(n_324), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_400), .B(n_369), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_380), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_397), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_400), .B(n_369), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_397), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_404), .B(n_369), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_388), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_380), .B(n_368), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_396), .B(n_347), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_403), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_403), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_404), .B(n_405), .Y(n_420) );
NAND3xp33_ASAP7_75t_SL g421 ( .A(n_387), .B(n_344), .C(n_366), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_388), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_374), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_396), .B(n_347), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_374), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_406), .B(n_371), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_389), .B(n_349), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_381), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_389), .B(n_386), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_381), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_388), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_382), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_382), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_401), .B(n_349), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_401), .B(n_365), .Y(n_435) );
AND2x2_ASAP7_75t_SL g436 ( .A(n_376), .B(n_367), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_384), .B(n_358), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_375), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_401), .B(n_365), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_406), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_401), .B(n_356), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_394), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_391), .B(n_361), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_375), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_391), .B(n_361), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_384), .B(n_348), .Y(n_446) );
AND2x6_ASAP7_75t_SL g447 ( .A(n_373), .B(n_357), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_404), .B(n_357), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_391), .B(n_361), .Y(n_449) );
INVx1_ASAP7_75t_SL g450 ( .A(n_376), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_399), .B(n_405), .Y(n_451) );
INVx1_ASAP7_75t_SL g452 ( .A(n_379), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_392), .B(n_367), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_386), .B(n_346), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_372), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_399), .B(n_343), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_394), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_405), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_372), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_394), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_426), .B(n_390), .Y(n_461) );
INVxp67_ASAP7_75t_SL g462 ( .A(n_440), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_411), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_438), .B(n_392), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_438), .B(n_392), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_435), .B(n_408), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_436), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_426), .B(n_390), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_411), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_413), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_441), .B(n_379), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_413), .Y(n_472) );
INVx2_ASAP7_75t_SL g473 ( .A(n_436), .Y(n_473) );
AND2x4_ASAP7_75t_L g474 ( .A(n_444), .B(n_383), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_435), .B(n_408), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_444), .B(n_407), .Y(n_476) );
OR2x6_ASAP7_75t_L g477 ( .A(n_448), .B(n_383), .Y(n_477) );
NAND2x1p5_ASAP7_75t_L g478 ( .A(n_436), .B(n_357), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_451), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_418), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_410), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_415), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_458), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_418), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_429), .B(n_407), .Y(n_485) );
NAND2x1_ASAP7_75t_L g486 ( .A(n_414), .B(n_383), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_437), .B(n_407), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_451), .B(n_402), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_416), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_419), .Y(n_490) );
INVxp67_ASAP7_75t_L g491 ( .A(n_420), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_439), .B(n_408), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_439), .B(n_385), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_419), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_423), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_415), .Y(n_496) );
INVxp67_ASAP7_75t_SL g497 ( .A(n_416), .Y(n_497) );
BUFx2_ASAP7_75t_L g498 ( .A(n_447), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_409), .B(n_385), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_427), .B(n_456), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_423), .Y(n_501) );
NOR2x1p5_ASAP7_75t_SL g502 ( .A(n_415), .B(n_398), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_454), .B(n_387), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_409), .B(n_412), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_425), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_454), .B(n_372), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_453), .B(n_398), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_446), .B(n_377), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_412), .B(n_385), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_425), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_450), .B(n_383), .Y(n_511) );
AND2x4_ASAP7_75t_L g512 ( .A(n_441), .B(n_377), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_428), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_434), .B(n_377), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_434), .B(n_402), .Y(n_515) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_422), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_422), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_453), .B(n_402), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_447), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_443), .B(n_398), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_504), .B(n_449), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_481), .Y(n_522) );
OR2x6_ASAP7_75t_L g523 ( .A(n_478), .B(n_414), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_481), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_504), .B(n_417), .Y(n_525) );
INVx1_ASAP7_75t_SL g526 ( .A(n_479), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_497), .B(n_445), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_489), .Y(n_528) );
OAI21xp5_ASAP7_75t_SL g529 ( .A1(n_519), .A2(n_421), .B(n_450), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_489), .B(n_452), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_503), .B(n_443), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_491), .B(n_452), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_466), .B(n_417), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_487), .B(n_449), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_466), .B(n_445), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_475), .B(n_428), .Y(n_536) );
AOI221xp5_ASAP7_75t_L g537 ( .A1(n_498), .A2(n_430), .B1(n_433), .B2(n_432), .C(n_414), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_475), .B(n_432), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_461), .Y(n_539) );
INVxp67_ASAP7_75t_L g540 ( .A(n_462), .Y(n_540) );
INVx1_ASAP7_75t_SL g541 ( .A(n_468), .Y(n_541) );
INVx3_ASAP7_75t_L g542 ( .A(n_478), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_499), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_482), .Y(n_544) );
NAND3xp33_ASAP7_75t_L g545 ( .A(n_483), .B(n_430), .C(n_433), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_500), .B(n_424), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_499), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_492), .B(n_459), .Y(n_548) );
OAI21xp33_ASAP7_75t_L g549 ( .A1(n_502), .A2(n_483), .B(n_485), .Y(n_549) );
INVx1_ASAP7_75t_SL g550 ( .A(n_509), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_464), .B(n_414), .Y(n_551) );
NOR3xp33_ASAP7_75t_L g552 ( .A(n_511), .B(n_333), .C(n_331), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_463), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_469), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_516), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_492), .B(n_424), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_493), .B(n_455), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_467), .B(n_460), .Y(n_558) );
INVx2_ASAP7_75t_SL g559 ( .A(n_486), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_470), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_520), .B(n_515), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_472), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_515), .B(n_460), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_493), .B(n_455), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_480), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_471), .B(n_460), .Y(n_566) );
OAI221xp5_ASAP7_75t_L g567 ( .A1(n_467), .A2(n_342), .B1(n_341), .B2(n_459), .C(n_442), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_512), .B(n_457), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_512), .B(n_457), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_465), .B(n_457), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_507), .B(n_442), .Y(n_571) );
INVx2_ASAP7_75t_SL g572 ( .A(n_530), .Y(n_572) );
NOR2xp33_ASAP7_75t_R g573 ( .A(n_542), .B(n_473), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_526), .Y(n_574) );
OAI21xp33_ASAP7_75t_SL g575 ( .A1(n_559), .A2(n_473), .B(n_511), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_544), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_521), .B(n_512), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_521), .B(n_520), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_531), .B(n_476), .Y(n_579) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_540), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_522), .Y(n_581) );
OAI21xp33_ASAP7_75t_SL g582 ( .A1(n_559), .A2(n_523), .B(n_537), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_524), .B(n_514), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_528), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_561), .B(n_509), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_553), .Y(n_586) );
AOI211xp5_ASAP7_75t_L g587 ( .A1(n_529), .A2(n_474), .B(n_508), .C(n_506), .Y(n_587) );
OAI22xp33_ASAP7_75t_L g588 ( .A1(n_523), .A2(n_542), .B1(n_477), .B2(n_545), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_523), .A2(n_477), .B1(n_474), .B2(n_488), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_540), .B(n_518), .Y(n_590) );
NAND2x1_ASAP7_75t_L g591 ( .A(n_542), .B(n_477), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_554), .Y(n_592) );
INVxp33_ASAP7_75t_L g593 ( .A(n_558), .Y(n_593) );
OAI221xp5_ASAP7_75t_SL g594 ( .A1(n_549), .A2(n_518), .B1(n_484), .B2(n_494), .C(n_490), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_561), .B(n_474), .Y(n_595) );
OAI21xp33_ASAP7_75t_SL g596 ( .A1(n_558), .A2(n_501), .B(n_495), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_551), .A2(n_505), .B1(n_513), .B2(n_510), .Y(n_597) );
OAI21xp5_ASAP7_75t_SL g598 ( .A1(n_567), .A2(n_357), .B(n_516), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_533), .B(n_517), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_539), .B(n_517), .Y(n_600) );
OAI221xp5_ASAP7_75t_L g601 ( .A1(n_532), .A2(n_496), .B1(n_482), .B2(n_431), .C(n_442), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_560), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_525), .B(n_496), .Y(n_603) );
OA21x2_ASAP7_75t_L g604 ( .A1(n_555), .A2(n_431), .B(n_422), .Y(n_604) );
INVxp67_ASAP7_75t_L g605 ( .A(n_532), .Y(n_605) );
OAI21xp5_ASAP7_75t_L g606 ( .A1(n_582), .A2(n_555), .B(n_552), .Y(n_606) );
OAI211xp5_ASAP7_75t_L g607 ( .A1(n_575), .A2(n_527), .B(n_552), .C(n_551), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g608 ( .A1(n_588), .A2(n_541), .B1(n_538), .B2(n_536), .C(n_547), .Y(n_608) );
AOI322xp5_ASAP7_75t_L g609 ( .A1(n_588), .A2(n_535), .A3(n_543), .B1(n_550), .B2(n_556), .C1(n_534), .C2(n_548), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_580), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_586), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_597), .B(n_565), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_578), .B(n_563), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_584), .B(n_562), .Y(n_614) );
OAI221xp5_ASAP7_75t_L g615 ( .A1(n_598), .A2(n_570), .B1(n_546), .B2(n_564), .C(n_557), .Y(n_615) );
OAI21xp33_ASAP7_75t_L g616 ( .A1(n_596), .A2(n_569), .B(n_568), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_587), .A2(n_571), .B1(n_566), .B2(n_544), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_581), .B(n_393), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_592), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_602), .Y(n_620) );
NAND2x1p5_ASAP7_75t_L g621 ( .A(n_591), .B(n_378), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_574), .B(n_431), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_578), .B(n_393), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_590), .Y(n_624) );
INVxp67_ASAP7_75t_SL g625 ( .A(n_600), .Y(n_625) );
AOI211xp5_ASAP7_75t_L g626 ( .A1(n_606), .A2(n_594), .B(n_589), .C(n_593), .Y(n_626) );
NOR4xp25_ASAP7_75t_L g627 ( .A(n_606), .B(n_605), .C(n_572), .D(n_601), .Y(n_627) );
NAND3xp33_ASAP7_75t_SL g628 ( .A(n_608), .B(n_573), .C(n_593), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_607), .A2(n_572), .B1(n_600), .B2(n_579), .Y(n_629) );
NAND4xp25_ASAP7_75t_L g630 ( .A(n_609), .B(n_595), .C(n_583), .D(n_577), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_625), .A2(n_604), .B(n_576), .Y(n_631) );
AOI211xp5_ASAP7_75t_L g632 ( .A1(n_615), .A2(n_573), .B(n_603), .C(n_585), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_612), .B(n_610), .Y(n_633) );
NAND3xp33_ASAP7_75t_L g634 ( .A(n_617), .B(n_604), .C(n_576), .Y(n_634) );
NOR3xp33_ASAP7_75t_SL g635 ( .A(n_616), .B(n_319), .C(n_322), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_621), .B(n_603), .Y(n_636) );
AOI322xp5_ASAP7_75t_L g637 ( .A1(n_628), .A2(n_624), .A3(n_613), .B1(n_623), .B2(n_622), .C1(n_599), .C2(n_620), .Y(n_637) );
AOI211xp5_ASAP7_75t_L g638 ( .A1(n_627), .A2(n_619), .B(n_611), .C(n_618), .Y(n_638) );
AOI211xp5_ASAP7_75t_L g639 ( .A1(n_626), .A2(n_614), .B(n_621), .C(n_393), .Y(n_639) );
OAI21xp5_ASAP7_75t_L g640 ( .A1(n_635), .A2(n_604), .B(n_378), .Y(n_640) );
AOI211xp5_ASAP7_75t_L g641 ( .A1(n_634), .A2(n_393), .B(n_373), .C(n_322), .Y(n_641) );
OAI321xp33_ASAP7_75t_L g642 ( .A1(n_632), .A2(n_393), .A3(n_395), .B1(n_334), .B2(n_345), .C(n_355), .Y(n_642) );
OR5x1_ASAP7_75t_L g643 ( .A(n_637), .B(n_630), .C(n_633), .D(n_629), .E(n_631), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_638), .Y(n_644) );
NOR3xp33_ASAP7_75t_L g645 ( .A(n_642), .B(n_636), .C(n_329), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_640), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_646), .Y(n_647) );
AND2x4_ASAP7_75t_L g648 ( .A(n_644), .B(n_639), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_648), .A2(n_641), .B1(n_643), .B2(n_645), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_648), .B(n_393), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_649), .B(n_647), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_651), .A2(n_650), .B1(n_355), .B2(n_395), .Y(n_652) );
AOI21xp5_ASAP7_75t_SL g653 ( .A1(n_652), .A2(n_345), .B(n_355), .Y(n_653) );
OA21x2_ASAP7_75t_L g654 ( .A1(n_653), .A2(n_329), .B(n_395), .Y(n_654) );
AOI21xp33_ASAP7_75t_L g655 ( .A1(n_654), .A2(n_324), .B(n_651), .Y(n_655) );
endmodule