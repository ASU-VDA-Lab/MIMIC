module fake_jpeg_10854_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_3),
.B(n_14),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_24),
.Y(n_49)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

CKINVDCx6p67_ASAP7_75t_R g130 ( 
.A(n_51),
.Y(n_130)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_53),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_5),
.C(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_87),
.Y(n_102)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_55),
.Y(n_135)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_27),
.B(n_2),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_57),
.B(n_58),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_16),
.B(n_15),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_30),
.B(n_2),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_63),
.B(n_73),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_40),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_65),
.Y(n_144)
);

BUFx4f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_72),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_4),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_78),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_17),
.B(n_4),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_79),
.B(n_95),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_82),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_84),
.B(n_88),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_86),
.Y(n_106)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_92),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_17),
.B(n_15),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_93),
.Y(n_134)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_94),
.B1(n_97),
.B2(n_44),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_18),
.B(n_6),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_44),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_51),
.Y(n_112)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_47),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_18),
.B(n_6),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_99),
.B(n_9),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_61),
.A2(n_38),
.B1(n_45),
.B2(n_43),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_100),
.A2(n_119),
.B1(n_67),
.B2(n_64),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_112),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_79),
.A2(n_35),
.B1(n_29),
.B2(n_21),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_113),
.A2(n_140),
.B1(n_105),
.B2(n_126),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_75),
.A2(n_34),
.B1(n_45),
.B2(n_43),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_63),
.B(n_35),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_29),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_59),
.A2(n_33),
.B1(n_36),
.B2(n_34),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_131),
.A2(n_146),
.B1(n_122),
.B2(n_144),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_21),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_138),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_73),
.A2(n_47),
.B1(n_33),
.B2(n_36),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_49),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_65),
.B(n_10),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_10),
.Y(n_169)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_144),
.A2(n_76),
.B1(n_51),
.B2(n_141),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_119),
.B1(n_102),
.B2(n_77),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_154),
.A2(n_155),
.B1(n_158),
.B2(n_170),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_169),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_62),
.B1(n_78),
.B2(n_83),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_130),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_166),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_101),
.B(n_109),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_175),
.C(n_130),
.Y(n_194)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

FAx1_ASAP7_75t_SL g166 ( 
.A(n_116),
.B(n_117),
.CI(n_127),
.CON(n_166),
.SN(n_166)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_111),
.A2(n_66),
.B1(n_44),
.B2(n_97),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_168),
.A2(n_171),
.B1(n_173),
.B2(n_181),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_136),
.A2(n_88),
.B1(n_91),
.B2(n_94),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_141),
.A2(n_0),
.B1(n_115),
.B2(n_129),
.Y(n_171)
);

NAND2xp33_ASAP7_75t_SL g172 ( 
.A(n_106),
.B(n_139),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_176),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_115),
.A2(n_126),
.B1(n_104),
.B2(n_123),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

INVx11_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_106),
.B(n_125),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

OAI32xp33_ASAP7_75t_L g180 ( 
.A1(n_107),
.A2(n_104),
.A3(n_121),
.B1(n_147),
.B2(n_137),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_118),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_132),
.A2(n_114),
.B1(n_142),
.B2(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_110),
.Y(n_183)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_157),
.A2(n_130),
.B(n_105),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_191),
.A2(n_163),
.B(n_183),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_159),
.C(n_153),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_195),
.A2(n_199),
.B1(n_201),
.B2(n_209),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_154),
.A2(n_120),
.B1(n_148),
.B2(n_142),
.Y(n_198)
);

OA22x2_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_212),
.B1(n_185),
.B2(n_184),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_176),
.A2(n_120),
.B1(n_142),
.B2(n_114),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_157),
.A2(n_108),
.B1(n_161),
.B2(n_166),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_166),
.A2(n_180),
.B1(n_175),
.B2(n_156),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_156),
.B(n_169),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_162),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_162),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_167),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_165),
.A2(n_159),
.B1(n_179),
.B2(n_178),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_227),
.Y(n_256)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_217),
.Y(n_249)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_213),
.Y(n_218)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_205),
.Y(n_221)
);

INVx13_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_202),
.A2(n_170),
.B1(n_164),
.B2(n_174),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_223),
.A2(n_234),
.B1(n_235),
.B2(n_206),
.Y(n_247)
);

INVx6_ASAP7_75t_SL g224 ( 
.A(n_205),
.Y(n_224)
);

INVx13_ASAP7_75t_L g255 ( 
.A(n_224),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_190),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_228),
.Y(n_254)
);

AND2x4_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_189),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_210),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_190),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_150),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_229),
.B(n_232),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_165),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_233),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_191),
.C(n_208),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_188),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_186),
.B(n_201),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_186),
.B(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_190),
.B(n_194),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_196),
.Y(n_248)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_224),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_245),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_252),
.C(n_231),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_225),
.A2(n_195),
.B1(n_199),
.B2(n_202),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_241),
.A2(n_219),
.B1(n_223),
.B2(n_230),
.Y(n_263)
);

AND2x6_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_198),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_246),
.A2(n_228),
.B1(n_222),
.B2(n_216),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_247),
.A2(n_219),
.B(n_217),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_231),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_203),
.C(n_196),
.Y(n_252)
);

AND2x6_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_206),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_253),
.B(n_234),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_242),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_259),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_269),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_250),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_265),
.C(n_267),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_263),
.B(n_271),
.Y(n_279)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_264),
.Y(n_276)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_240),
.Y(n_266)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_215),
.C(n_219),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_268),
.A2(n_247),
.B1(n_243),
.B2(n_241),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_232),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_229),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_256),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_203),
.C(n_235),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_256),
.C(n_254),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_272),
.B(n_270),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_260),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_258),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_284),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_273),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_285),
.B(n_269),
.Y(n_289)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_263),
.Y(n_287)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_287),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_286),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_292),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_289),
.B(n_293),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_265),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_282),
.A2(n_249),
.B(n_268),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_294),
.A2(n_243),
.B(n_278),
.Y(n_305)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_286),
.Y(n_295)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_272),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_298),
.C(n_271),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_267),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_281),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_307),
.C(n_293),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_290),
.A2(n_275),
.B(n_287),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_309),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_279),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_304),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_279),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_305),
.A2(n_308),
.B1(n_309),
.B2(n_301),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_283),
.B1(n_284),
.B2(n_278),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_310),
.B(n_312),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_314),
.C(n_316),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_292),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_317),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_298),
.C(n_291),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_289),
.C(n_285),
.Y(n_316)
);

OAI322xp33_ASAP7_75t_L g317 ( 
.A1(n_302),
.A2(n_253),
.A3(n_245),
.B1(n_276),
.B2(n_274),
.C1(n_250),
.C2(n_255),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_312),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_322),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_276),
.C(n_274),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_321),
.B(n_238),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_221),
.Y(n_322)
);

AOI322xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_255),
.A3(n_237),
.B1(n_238),
.B2(n_313),
.C1(n_246),
.C2(n_224),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_325),
.A2(n_192),
.B1(n_214),
.B2(n_193),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_327),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_220),
.Y(n_327)
);

AO21x1_ASAP7_75t_L g328 ( 
.A1(n_323),
.A2(n_218),
.B(n_246),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_246),
.C(n_226),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_329),
.A2(n_324),
.B(n_330),
.Y(n_332)
);

OAI21x1_ASAP7_75t_SL g333 ( 
.A1(n_331),
.A2(n_192),
.B(n_226),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_333),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_319),
.B1(n_226),
.B2(n_193),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_226),
.B1(n_214),
.B2(n_200),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_197),
.Y(n_337)
);


endmodule