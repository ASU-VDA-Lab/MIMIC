module fake_ariane_2896_n_493 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_493);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_493;

wire n_295;
wire n_356;
wire n_190;
wire n_180;
wire n_386;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_373;
wire n_299;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_319;
wire n_416;
wire n_283;
wire n_187;
wire n_367;
wire n_374;
wire n_345;
wire n_318;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_424;
wire n_387;
wire n_406;
wire n_391;
wire n_349;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_462;
wire n_410;
wire n_379;
wire n_445;
wire n_264;
wire n_198;
wire n_232;
wire n_441;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_422;
wire n_269;
wire n_259;
wire n_446;
wire n_405;
wire n_173;
wire n_242;
wire n_309;
wire n_331;
wire n_320;
wire n_401;
wire n_485;
wire n_267;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_398;
wire n_210;
wire n_200;
wire n_253;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_247;
wire n_240;
wire n_369;
wire n_224;
wire n_420;
wire n_439;
wire n_222;
wire n_478;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_330;
wire n_400;
wire n_282;
wire n_328;
wire n_368;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_427;
wire n_303;
wire n_442;
wire n_206;
wire n_352;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_334;
wire n_192;
wire n_488;
wire n_300;
wire n_390;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_260;
wire n_362;
wire n_310;
wire n_236;
wire n_281;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_464;
wire n_297;
wire n_290;
wire n_371;
wire n_199;
wire n_452;
wire n_217;
wire n_178;
wire n_308;
wire n_417;
wire n_201;
wire n_343;
wire n_414;
wire n_287;
wire n_302;
wire n_380;
wire n_284;
wire n_448;
wire n_249;
wire n_355;
wire n_212;
wire n_444;
wire n_278;
wire n_255;
wire n_450;
wire n_257;
wire n_451;
wire n_475;
wire n_409;
wire n_384;
wire n_468;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_407;
wire n_254;
wire n_476;
wire n_460;
wire n_219;
wire n_231;
wire n_366;
wire n_234;
wire n_492;
wire n_280;
wire n_215;
wire n_252;
wire n_454;
wire n_298;
wire n_415;
wire n_216;
wire n_418;
wire n_223;
wire n_403;
wire n_389;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_213;
wire n_304;
wire n_306;
wire n_313;
wire n_430;
wire n_203;
wire n_378;
wire n_436;
wire n_375;
wire n_324;
wire n_337;
wire n_437;
wire n_274;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_292;
wire n_174;
wire n_275;
wire n_204;
wire n_342;
wire n_246;
wire n_428;
wire n_358;
wire n_263;
wire n_434;
wire n_360;
wire n_229;
wire n_394;
wire n_250;
wire n_317;
wire n_243;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_408;
wire n_322;
wire n_251;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_359;

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_102),
.B(n_0),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_144),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_12),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_41),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_28),
.B(n_86),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_7),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_157),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_6),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_25),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_15),
.B(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

INVxp33_ASAP7_75t_SL g184 ( 
.A(n_126),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_88),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_166),
.Y(n_187)
);

INVxp67_ASAP7_75t_SL g188 ( 
.A(n_101),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

BUFx2_ASAP7_75t_SL g190 ( 
.A(n_118),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_89),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_16),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_40),
.B(n_132),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_130),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_64),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_149),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_75),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_111),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_81),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_2),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_121),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_120),
.B(n_99),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_55),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_138),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_83),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_19),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_24),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_3),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_131),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_34),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_2),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_57),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_11),
.B(n_104),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_107),
.B(n_105),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_74),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_8),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_33),
.Y(n_221)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_106),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_66),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_L g224 ( 
.A(n_48),
.B(n_71),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_17),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g226 ( 
.A(n_36),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_59),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_143),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_9),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_82),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_45),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_69),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_127),
.Y(n_233)
);

INVxp67_ASAP7_75t_SL g234 ( 
.A(n_42),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_39),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_49),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_90),
.B(n_134),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_100),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_51),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_78),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_76),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_112),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_60),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_26),
.B(n_161),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_62),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_113),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_94),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_156),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_167),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_29),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_38),
.B(n_20),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_170),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_73),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_87),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_117),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_165),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_27),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_13),
.B(n_5),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_162),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_145),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_85),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_37),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_30),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_140),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_152),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_70),
.Y(n_266)
);

INVxp33_ASAP7_75t_SL g267 ( 
.A(n_160),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_163),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_137),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_10),
.B(n_4),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_92),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_44),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_109),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_97),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_1),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_153),
.B(n_151),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_159),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_95),
.Y(n_278)
);

NOR2xp67_ASAP7_75t_L g279 ( 
.A(n_21),
.B(n_68),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_65),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_80),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_0),
.B(n_164),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_63),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_31),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_91),
.Y(n_285)
);

INVxp67_ASAP7_75t_SL g286 ( 
.A(n_139),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_72),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_3),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_129),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_148),
.B(n_61),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_50),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_43),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_35),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_56),
.Y(n_294)
);

INVxp33_ASAP7_75t_SL g295 ( 
.A(n_22),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_108),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_275),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_210),
.B(n_1),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_191),
.Y(n_299)
);

AND2x6_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_14),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_288),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_179),
.B(n_18),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_178),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_203),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_221),
.Y(n_305)
);

AO22x2_ASAP7_75t_L g306 ( 
.A1(n_175),
.A2(n_23),
.B1(n_32),
.B2(n_46),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_245),
.B(n_47),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_281),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_52),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_212),
.B(n_53),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_194),
.B(n_54),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_177),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_180),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_191),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_183),
.B(n_58),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_191),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_186),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_189),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_195),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_191),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_196),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_181),
.Y(n_322)
);

NAND2x1p5_ASAP7_75t_L g323 ( 
.A(n_263),
.B(n_67),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_197),
.B(n_77),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_198),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_199),
.B(n_79),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_200),
.B(n_84),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_201),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_202),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_206),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_215),
.B(n_93),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_207),
.Y(n_332)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_173),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_225),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_208),
.Y(n_335)
);

BUFx10_ASAP7_75t_L g336 ( 
.A(n_172),
.Y(n_336)
);

NAND3xp33_ASAP7_75t_L g337 ( 
.A(n_243),
.B(n_96),
.C(n_98),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_209),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_211),
.Y(n_339)
);

OR2x2_ASAP7_75t_SL g340 ( 
.A(n_268),
.B(n_103),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_214),
.B(n_110),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_219),
.Y(n_342)
);

NAND3xp33_ASAP7_75t_L g343 ( 
.A(n_199),
.B(n_114),
.C(n_115),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_220),
.B(n_116),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_227),
.B(n_119),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_228),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_230),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_260),
.B(n_122),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_235),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_242),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_247),
.B(n_124),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_248),
.B(n_125),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_252),
.B(n_133),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_257),
.B(n_135),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_232),
.A2(n_158),
.B1(n_147),
.B2(n_150),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_262),
.Y(n_356)
);

INVx2_ASAP7_75t_SL g357 ( 
.A(n_265),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_269),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_271),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_273),
.B(n_136),
.Y(n_360)
);

INVx4_ASAP7_75t_SL g361 ( 
.A(n_274),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_284),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_307),
.B(n_184),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_311),
.B(n_267),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_326),
.B(n_295),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_336),
.B(n_233),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_333),
.B(n_312),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_353),
.B(n_278),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_303),
.B(n_190),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_309),
.B(n_240),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_351),
.B(n_310),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_331),
.B(n_250),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_322),
.B(n_246),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_334),
.B(n_294),
.Y(n_374)
);

NAND2xp33_ASAP7_75t_SL g375 ( 
.A(n_298),
.B(n_293),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_348),
.B(n_216),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_305),
.B(n_229),
.Y(n_377)
);

NAND2xp33_ASAP7_75t_SL g378 ( 
.A(n_302),
.B(n_255),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_308),
.B(n_261),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_304),
.B(n_292),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_359),
.B(n_291),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_359),
.B(n_192),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_321),
.B(n_272),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_335),
.B(n_266),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_317),
.B(n_231),
.Y(n_385)
);

NAND2xp33_ASAP7_75t_SL g386 ( 
.A(n_355),
.B(n_239),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_318),
.B(n_264),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_319),
.B(n_187),
.Y(n_388)
);

XNOR2x2_ASAP7_75t_L g389 ( 
.A(n_306),
.B(n_282),
.Y(n_389)
);

NAND2xp33_ASAP7_75t_SL g390 ( 
.A(n_315),
.B(n_259),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_340),
.B(n_238),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_325),
.B(n_236),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_329),
.B(n_287),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_338),
.B(n_253),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_346),
.B(n_280),
.Y(n_395)
);

NAND2xp33_ASAP7_75t_SL g396 ( 
.A(n_324),
.B(n_254),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_357),
.B(n_204),
.Y(n_397)
);

NAND2xp33_ASAP7_75t_SL g398 ( 
.A(n_327),
.B(n_256),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_347),
.B(n_223),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_350),
.B(n_285),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_358),
.B(n_185),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_362),
.B(n_283),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_323),
.B(n_174),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_391),
.B(n_300),
.Y(n_404)
);

AO21x1_ASAP7_75t_L g405 ( 
.A1(n_386),
.A2(n_341),
.B(n_344),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_393),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_373),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_369),
.B(n_328),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_399),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_374),
.B(n_330),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_395),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g412 ( 
.A(n_380),
.B(n_342),
.Y(n_412)
);

AOI221xp5_ASAP7_75t_L g413 ( 
.A1(n_375),
.A2(n_301),
.B1(n_297),
.B2(n_345),
.C(n_349),
.Y(n_413)
);

OAI21x1_ASAP7_75t_L g414 ( 
.A1(n_370),
.A2(n_354),
.B(n_360),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_401),
.A2(n_300),
.B(n_352),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_371),
.B(n_300),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_380),
.B(n_356),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_367),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_332),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_397),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_364),
.B(n_339),
.Y(n_421)
);

AO21x2_ASAP7_75t_L g422 ( 
.A1(n_403),
.A2(n_337),
.B(n_343),
.Y(n_422)
);

OAI21x1_ASAP7_75t_L g423 ( 
.A1(n_376),
.A2(n_244),
.B(n_237),
.Y(n_423)
);

BUFx10_ASAP7_75t_L g424 ( 
.A(n_389),
.Y(n_424)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_385),
.A2(n_205),
.B(n_313),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_365),
.B(n_361),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_387),
.Y(n_427)
);

OAI221xp5_ASAP7_75t_L g428 ( 
.A1(n_378),
.A2(n_226),
.B1(n_286),
.B2(n_188),
.C(n_234),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_388),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_377),
.B(n_361),
.Y(n_430)
);

OAI21x1_ASAP7_75t_L g431 ( 
.A1(n_392),
.A2(n_222),
.B(n_279),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_394),
.A2(n_224),
.B(n_176),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_390),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_363),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_420),
.B(n_366),
.Y(n_435)
);

OR2x6_ASAP7_75t_L g436 ( 
.A(n_407),
.B(n_379),
.Y(n_436)
);

INVx5_ASAP7_75t_L g437 ( 
.A(n_419),
.Y(n_437)
);

NAND3xp33_ASAP7_75t_SL g438 ( 
.A(n_405),
.B(n_372),
.C(n_398),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_R g439 ( 
.A(n_410),
.B(n_396),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_419),
.B(n_368),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_417),
.B(n_384),
.Y(n_441)
);

NAND2xp33_ASAP7_75t_SL g442 ( 
.A(n_418),
.B(n_277),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_417),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_404),
.B(n_402),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_408),
.B(n_383),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_421),
.Y(n_446)
);

NAND2xp33_ASAP7_75t_R g447 ( 
.A(n_416),
.B(n_213),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_411),
.B(n_412),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_406),
.B(n_400),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_R g450 ( 
.A(n_430),
.B(n_270),
.Y(n_450)
);

NAND2xp33_ASAP7_75t_R g451 ( 
.A(n_430),
.B(n_258),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_448),
.B(n_406),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_434),
.B(n_409),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_424),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_437),
.B(n_424),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_446),
.Y(n_456)
);

NOR2x2_ASAP7_75t_L g457 ( 
.A(n_436),
.B(n_429),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_445),
.Y(n_458)
);

AOI221xp5_ASAP7_75t_L g459 ( 
.A1(n_442),
.A2(n_428),
.B1(n_413),
.B2(n_409),
.C(n_432),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_433),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_436),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_427),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_449),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_441),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_435),
.B(n_426),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_438),
.Y(n_466)
);

A2O1A1Ixp33_ASAP7_75t_L g467 ( 
.A1(n_459),
.A2(n_415),
.B(n_444),
.C(n_414),
.Y(n_467)
);

OR2x6_ASAP7_75t_L g468 ( 
.A(n_454),
.B(n_431),
.Y(n_468)
);

NAND2xp33_ASAP7_75t_R g469 ( 
.A(n_455),
.B(n_423),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_459),
.A2(n_439),
.B1(n_451),
.B2(n_450),
.Y(n_470)
);

NOR2x1_ASAP7_75t_L g471 ( 
.A(n_453),
.B(n_249),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_453),
.B(n_422),
.Y(n_472)
);

AO221x2_ASAP7_75t_L g473 ( 
.A1(n_463),
.A2(n_289),
.B1(n_241),
.B2(n_447),
.C(n_422),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_382),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_461),
.Y(n_475)
);

AOI222xp33_ASAP7_75t_L g476 ( 
.A1(n_470),
.A2(n_456),
.B1(n_464),
.B2(n_460),
.C1(n_471),
.C2(n_474),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_466),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_472),
.B(n_462),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_473),
.B(n_465),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_468),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_468),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_475),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_482),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_477),
.B(n_467),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_481),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_483),
.A2(n_476),
.B1(n_479),
.B2(n_469),
.Y(n_486)
);

NOR4xp75_ASAP7_75t_L g487 ( 
.A(n_484),
.B(n_381),
.C(n_478),
.D(n_476),
.Y(n_487)
);

AOI222xp33_ASAP7_75t_L g488 ( 
.A1(n_485),
.A2(n_480),
.B1(n_182),
.B2(n_193),
.C1(n_217),
.C2(n_218),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_R g489 ( 
.A(n_486),
.B(n_154),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_489),
.Y(n_490)
);

AOI31xp33_ASAP7_75t_L g491 ( 
.A1(n_490),
.A2(n_488),
.A3(n_487),
.B(n_251),
.Y(n_491)
);

AOI222xp33_ASAP7_75t_L g492 ( 
.A1(n_491),
.A2(n_290),
.B1(n_425),
.B2(n_457),
.C1(n_316),
.C2(n_320),
.Y(n_492)
);

OAI221xp5_ASAP7_75t_R g493 ( 
.A1(n_492),
.A2(n_299),
.B1(n_314),
.B2(n_316),
.C(n_320),
.Y(n_493)
);


endmodule