module fake_jpeg_17077_n_274 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_274);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_22),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_19),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_59),
.Y(n_79)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_49),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_17),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_25),
.C(n_17),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_16),
.Y(n_54)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_16),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_57),
.Y(n_82)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NAND2x1_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_25),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_18),
.B1(n_32),
.B2(n_20),
.Y(n_72)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_39),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_63),
.A2(n_18),
.B1(n_17),
.B2(n_19),
.Y(n_66)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_81),
.B(n_88),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_69),
.B(n_51),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_40),
.B1(n_25),
.B2(n_24),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_70),
.A2(n_84),
.B1(n_63),
.B2(n_56),
.Y(n_106)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_18),
.B1(n_19),
.B2(n_28),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_73),
.A2(n_87),
.B1(n_61),
.B2(n_56),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_80),
.Y(n_95)
);

OA22x2_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_24),
.B1(n_32),
.B2(n_20),
.Y(n_77)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_28),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_25),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_48),
.A2(n_18),
.B1(n_28),
.B2(n_21),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_40),
.B1(n_25),
.B2(n_23),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_51),
.A2(n_21),
.B1(n_29),
.B2(n_27),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_44),
.A2(n_21),
.B1(n_29),
.B2(n_26),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_101),
.Y(n_118)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_44),
.B1(n_47),
.B2(n_61),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_100),
.B1(n_102),
.B2(n_106),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_85),
.B(n_70),
.Y(n_123)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_64),
.B1(n_26),
.B2(n_27),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_60),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_68),
.A2(n_50),
.B1(n_23),
.B2(n_45),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_107),
.A2(n_86),
.B1(n_82),
.B2(n_74),
.Y(n_117)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_111),
.Y(n_127)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_73),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_85),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_80),
.Y(n_131)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_77),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_53),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_79),
.B1(n_76),
.B2(n_78),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_95),
.B1(n_90),
.B2(n_102),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_117),
.B(n_126),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_69),
.C(n_79),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_123),
.Y(n_144)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_70),
.C(n_82),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_125),
.A2(n_31),
.B(n_22),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_98),
.Y(n_126)
);

AO22x1_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_70),
.B1(n_84),
.B2(n_50),
.Y(n_128)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_131),
.B(n_137),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_84),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_136),
.Y(n_157)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_92),
.B(n_84),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_98),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_109),
.B1(n_91),
.B2(n_90),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_141),
.A2(n_154),
.B(n_166),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_112),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_150),
.Y(n_176)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_95),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_145),
.B(n_146),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_91),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_93),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_149),
.Y(n_170)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_104),
.B1(n_105),
.B2(n_110),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_151),
.A2(n_164),
.B1(n_122),
.B2(n_134),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_131),
.B(n_113),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_153),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_45),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_99),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_156),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_119),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_158),
.Y(n_181)
);

INVxp33_ASAP7_75t_SL g159 ( 
.A(n_124),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_159),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_53),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_161),
.B(n_8),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_22),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_130),
.Y(n_167)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_163),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_127),
.A2(n_46),
.B1(n_9),
.B2(n_3),
.Y(n_164)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_120),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_146),
.A2(n_136),
.B1(n_118),
.B2(n_121),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_168),
.A2(n_174),
.B1(n_179),
.B2(n_151),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_115),
.C(n_119),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_173),
.C(n_187),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_117),
.Y(n_173)
);

AOI221xp5_ASAP7_75t_L g177 ( 
.A1(n_161),
.A2(n_128),
.B1(n_124),
.B2(n_116),
.C(n_122),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_177),
.B(n_185),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_128),
.B1(n_134),
.B2(n_138),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_152),
.A2(n_9),
.B1(n_15),
.B2(n_3),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_157),
.A2(n_0),
.B(n_2),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_0),
.Y(n_186)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_186),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_46),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_175),
.C(n_182),
.Y(n_192)
);

OAI21x1_ASAP7_75t_L g189 ( 
.A1(n_166),
.A2(n_8),
.B(n_3),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_141),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_154),
.Y(n_191)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_192),
.A2(n_198),
.B1(n_180),
.B2(n_4),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_176),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_201),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_143),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_183),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_150),
.Y(n_197)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_152),
.B1(n_149),
.B2(n_147),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_148),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_162),
.C(n_145),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_179),
.C(n_173),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_184),
.B1(n_186),
.B2(n_174),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_163),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_204),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_140),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_205),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_164),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_208),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_155),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_210),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_155),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_226),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_187),
.C(n_175),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_213),
.B(n_221),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_198),
.A2(n_183),
.B(n_178),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_208),
.B(n_196),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_222),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_219),
.A2(n_224),
.B1(n_193),
.B2(n_201),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_188),
.C(n_165),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_180),
.B1(n_0),
.B2(n_5),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_4),
.C(n_5),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_204),
.B(n_210),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_229),
.B(n_207),
.Y(n_242)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_223),
.A2(n_200),
.B1(n_191),
.B2(n_209),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_234),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_218),
.A2(n_196),
.B(n_195),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_221),
.C(n_211),
.Y(n_239)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_237),
.Y(n_244)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_238),
.B(n_219),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_240),
.C(n_242),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_213),
.C(n_216),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_L g241 ( 
.A1(n_229),
.A2(n_214),
.B(n_215),
.Y(n_241)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_226),
.C(n_225),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_248),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_244),
.B(n_234),
.Y(n_251)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_251),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_231),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_252),
.B(n_250),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_233),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_6),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_241),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_245),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_247),
.A2(n_192),
.B1(n_233),
.B2(n_207),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_256),
.A2(n_236),
.B(n_6),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_260),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_259),
.A2(n_256),
.B(n_10),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_L g261 ( 
.A1(n_254),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_10),
.C2(n_11),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_262),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_263),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_259),
.A2(n_249),
.B(n_255),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_7),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_12),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_269),
.Y(n_271)
);

OAI321xp33_ASAP7_75t_L g272 ( 
.A1(n_271),
.A2(n_270),
.A3(n_266),
.B1(n_268),
.B2(n_264),
.C(n_14),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_272),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_14),
.Y(n_274)
);


endmodule