module real_aes_511_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_735;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_0), .B(n_145), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_1), .A2(n_154), .B(n_159), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_2), .B(n_784), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_3), .B(n_145), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_4), .B(n_161), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_5), .B(n_161), .Y(n_199) );
INVx1_ASAP7_75t_L g152 ( .A(n_6), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_7), .B(n_161), .Y(n_227) );
CKINVDCx16_ASAP7_75t_R g784 ( .A(n_8), .Y(n_784) );
NAND2xp33_ASAP7_75t_L g188 ( .A(n_9), .B(n_163), .Y(n_188) );
AND2x2_ASAP7_75t_L g498 ( .A(n_10), .B(n_182), .Y(n_498) );
AND2x2_ASAP7_75t_L g506 ( .A(n_11), .B(n_139), .Y(n_506) );
INVx2_ASAP7_75t_L g142 ( .A(n_12), .Y(n_142) );
AOI221x1_ASAP7_75t_L g234 ( .A1(n_13), .A2(n_24), .B1(n_145), .B2(n_154), .C(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_14), .B(n_161), .Y(n_458) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_15), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_16), .B(n_145), .Y(n_184) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_17), .A2(n_182), .B(n_183), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_18), .B(n_165), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_19), .B(n_161), .Y(n_175) );
AO21x1_ASAP7_75t_L g194 ( .A1(n_20), .A2(n_145), .B(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_21), .B(n_145), .Y(n_479) );
INVx1_ASAP7_75t_L g118 ( .A(n_22), .Y(n_118) );
NOR2xp33_ASAP7_75t_SL g781 ( .A(n_22), .B(n_119), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_23), .A2(n_90), .B1(n_145), .B2(n_514), .Y(n_513) );
NAND2x1_ASAP7_75t_L g207 ( .A(n_25), .B(n_161), .Y(n_207) );
NAND2x1_ASAP7_75t_L g226 ( .A(n_26), .B(n_163), .Y(n_226) );
OAI22xp5_ASAP7_75t_SL g774 ( .A1(n_27), .A2(n_63), .B1(n_775), .B2(n_776), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_27), .Y(n_775) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_28), .A2(n_87), .B(n_142), .Y(n_141) );
OR2x2_ASAP7_75t_L g167 ( .A(n_28), .B(n_87), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_29), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_30), .B(n_161), .Y(n_187) );
AO21x2_ASAP7_75t_L g453 ( .A1(n_31), .A2(n_139), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_32), .B(n_163), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_33), .A2(n_154), .B(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_34), .B(n_161), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_35), .A2(n_154), .B(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g151 ( .A(n_36), .B(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_L g155 ( .A(n_36), .B(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g522 ( .A(n_36), .Y(n_522) );
OR2x6_ASAP7_75t_L g116 ( .A(n_37), .B(n_117), .Y(n_116) );
NOR3xp33_ASAP7_75t_L g782 ( .A(n_37), .B(n_783), .C(n_785), .Y(n_782) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_38), .B(n_145), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_39), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_40), .B(n_145), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_41), .B(n_161), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_42), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_43), .B(n_163), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_44), .B(n_145), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_45), .A2(n_154), .B(n_502), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_46), .A2(n_154), .B(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_47), .B(n_163), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_48), .A2(n_52), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_48), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_49), .B(n_163), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_50), .B(n_145), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_51), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_52), .Y(n_123) );
INVx1_ASAP7_75t_L g148 ( .A(n_53), .Y(n_148) );
INVx1_ASAP7_75t_L g158 ( .A(n_53), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_54), .B(n_161), .Y(n_504) );
AND2x2_ASAP7_75t_L g470 ( .A(n_55), .B(n_165), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_56), .B(n_163), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_57), .B(n_161), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_58), .B(n_163), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_59), .A2(n_154), .B(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_60), .B(n_145), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_61), .B(n_145), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_62), .A2(n_154), .B(n_463), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_63), .Y(n_776) );
AO21x1_ASAP7_75t_L g196 ( .A1(n_64), .A2(n_154), .B(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g485 ( .A(n_65), .B(n_166), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_66), .B(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_67), .B(n_163), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_68), .B(n_145), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_69), .B(n_163), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_70), .A2(n_95), .B1(n_154), .B2(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g219 ( .A(n_71), .B(n_166), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_72), .B(n_161), .Y(n_482) );
INVx1_ASAP7_75t_L g150 ( .A(n_73), .Y(n_150) );
INVx1_ASAP7_75t_L g156 ( .A(n_73), .Y(n_156) );
AND2x2_ASAP7_75t_L g230 ( .A(n_74), .B(n_139), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_75), .B(n_163), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_76), .A2(n_154), .B(n_474), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_77), .A2(n_154), .B(n_543), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_78), .A2(n_154), .B(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g467 ( .A(n_79), .B(n_166), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_80), .B(n_165), .Y(n_511) );
INVx1_ASAP7_75t_L g119 ( .A(n_81), .Y(n_119) );
AND2x2_ASAP7_75t_L g138 ( .A(n_82), .B(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_83), .B(n_145), .Y(n_177) );
AND2x2_ASAP7_75t_L g546 ( .A(n_84), .B(n_182), .Y(n_546) );
AND2x2_ASAP7_75t_L g195 ( .A(n_85), .B(n_171), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_86), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_88), .B(n_163), .Y(n_176) );
AND2x2_ASAP7_75t_L g211 ( .A(n_89), .B(n_139), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_91), .B(n_161), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_92), .A2(n_154), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_93), .B(n_163), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_94), .A2(n_154), .B(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_96), .B(n_161), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_97), .B(n_161), .Y(n_160) );
BUFx2_ASAP7_75t_L g484 ( .A(n_98), .Y(n_484) );
BUFx2_ASAP7_75t_L g106 ( .A(n_99), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_100), .A2(n_154), .B(n_186), .Y(n_185) );
AOI21xp33_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_780), .B(n_786), .Y(n_101) );
OA21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_121), .B(n_769), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_106), .Y(n_770) );
INVxp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g771 ( .A1(n_108), .A2(n_772), .B(n_777), .Y(n_771) );
NOR2xp33_ASAP7_75t_SL g108 ( .A(n_109), .B(n_120), .Y(n_108) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
BUFx3_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g779 ( .A(n_113), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
OR2x6_ASAP7_75t_SL g129 ( .A(n_114), .B(n_115), .Y(n_129) );
AND2x6_ASAP7_75t_SL g759 ( .A(n_114), .B(n_116), .Y(n_759) );
OR2x2_ASAP7_75t_L g768 ( .A(n_114), .B(n_116), .Y(n_768) );
CKINVDCx16_ASAP7_75t_R g785 ( .A(n_114), .Y(n_785) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_125), .B(n_760), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g760 ( .A1(n_122), .A2(n_761), .B(n_765), .Y(n_760) );
INVxp67_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_130), .B1(n_447), .B2(n_756), .Y(n_126) );
INVx1_ASAP7_75t_SL g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g764 ( .A(n_128), .Y(n_764) );
CKINVDCx11_ASAP7_75t_R g128 ( .A(n_129), .Y(n_128) );
INVx3_ASAP7_75t_L g763 ( .A(n_130), .Y(n_763) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_356), .Y(n_130) );
NOR4xp25_ASAP7_75t_L g131 ( .A(n_132), .B(n_274), .C(n_300), .D(n_340), .Y(n_131) );
OAI211xp5_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_189), .B(n_220), .C(n_260), .Y(n_132) );
INVxp67_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_168), .Y(n_134) );
AND2x2_ASAP7_75t_L g427 ( .A(n_135), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_136), .B(n_168), .Y(n_294) );
BUFx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g221 ( .A(n_137), .B(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_137), .B(n_247), .Y(n_246) );
INVx5_ASAP7_75t_L g280 ( .A(n_137), .Y(n_280) );
NOR2x1_ASAP7_75t_SL g322 ( .A(n_137), .B(n_169), .Y(n_322) );
AND2x2_ASAP7_75t_L g378 ( .A(n_137), .B(n_181), .Y(n_378) );
OR2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_143), .Y(n_137) );
INVx3_ASAP7_75t_L g210 ( .A(n_139), .Y(n_210) );
INVx4_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_140), .A2(n_500), .B(n_506), .Y(n_499) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx4f_ASAP7_75t_L g182 ( .A(n_141), .Y(n_182) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_142), .B(n_167), .Y(n_166) );
AND2x4_ASAP7_75t_L g171 ( .A(n_142), .B(n_167), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_153), .B(n_165), .Y(n_143) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_151), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
AND2x6_ASAP7_75t_L g163 ( .A(n_147), .B(n_156), .Y(n_163) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_L g161 ( .A(n_149), .B(n_158), .Y(n_161) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx5_ASAP7_75t_L g164 ( .A(n_151), .Y(n_164) );
AND2x2_ASAP7_75t_L g157 ( .A(n_152), .B(n_158), .Y(n_157) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_152), .Y(n_517) );
AND2x6_ASAP7_75t_L g154 ( .A(n_155), .B(n_157), .Y(n_154) );
BUFx3_ASAP7_75t_L g518 ( .A(n_155), .Y(n_518) );
INVx2_ASAP7_75t_L g524 ( .A(n_156), .Y(n_524) );
AND2x4_ASAP7_75t_L g520 ( .A(n_157), .B(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g516 ( .A(n_158), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_162), .B(n_164), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_163), .B(n_484), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_164), .A2(n_175), .B(n_176), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_164), .A2(n_187), .B(n_188), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_164), .A2(n_198), .B(n_199), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_164), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_164), .A2(n_216), .B(n_217), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_164), .A2(n_226), .B(n_227), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_164), .A2(n_236), .B(n_237), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_164), .A2(n_458), .B(n_459), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_164), .A2(n_464), .B(n_465), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_164), .A2(n_475), .B(n_476), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_164), .A2(n_482), .B(n_483), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_164), .A2(n_495), .B(n_496), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_164), .A2(n_503), .B(n_504), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_164), .A2(n_544), .B(n_545), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_165), .Y(n_229) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_165), .A2(n_234), .B(n_238), .Y(n_233) );
OA21x2_ASAP7_75t_L g273 ( .A1(n_165), .A2(n_234), .B(n_238), .Y(n_273) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_165), .A2(n_513), .B(n_519), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_165), .A2(n_541), .B(n_542), .Y(n_540) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_180), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_169), .B(n_181), .Y(n_250) );
AND2x2_ASAP7_75t_L g311 ( .A(n_169), .B(n_280), .Y(n_311) );
AO21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_172), .B(n_178), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_170), .B(n_179), .Y(n_178) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_170), .A2(n_172), .B(n_178), .Y(n_264) );
INVx1_ASAP7_75t_SL g170 ( .A(n_171), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_171), .A2(n_184), .B(n_185), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_171), .B(n_201), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_171), .A2(n_455), .B(n_456), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_171), .A2(n_472), .B(n_473), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_177), .Y(n_172) );
AND2x2_ASAP7_75t_L g323 ( .A(n_180), .B(n_247), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_180), .B(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g367 ( .A(n_180), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g400 ( .A(n_180), .B(n_221), .Y(n_400) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g244 ( .A(n_181), .Y(n_244) );
AND2x2_ASAP7_75t_L g277 ( .A(n_181), .B(n_278), .Y(n_277) );
BUFx3_ASAP7_75t_L g312 ( .A(n_181), .Y(n_312) );
OR2x2_ASAP7_75t_L g388 ( .A(n_181), .B(n_247), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_182), .A2(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_SL g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_202), .Y(n_190) );
AOI211x1_ASAP7_75t_SL g317 ( .A1(n_191), .A2(n_309), .B(n_318), .C(n_320), .Y(n_317) );
AND2x2_ASAP7_75t_SL g362 ( .A(n_191), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_191), .B(n_360), .Y(n_407) );
BUFx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g257 ( .A(n_192), .Y(n_257) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g232 ( .A(n_193), .Y(n_232) );
OAI21x1_ASAP7_75t_SL g193 ( .A1(n_194), .A2(n_196), .B(n_200), .Y(n_193) );
INVx1_ASAP7_75t_L g201 ( .A(n_195), .Y(n_201) );
AOI322xp5_ASAP7_75t_L g220 ( .A1(n_202), .A2(n_221), .A3(n_231), .B1(n_239), .B2(n_242), .C1(n_248), .C2(n_251), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_202), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_212), .Y(n_202) );
INVx2_ASAP7_75t_L g255 ( .A(n_203), .Y(n_255) );
INVxp67_ASAP7_75t_L g297 ( .A(n_203), .Y(n_297) );
BUFx3_ASAP7_75t_L g361 ( .A(n_203), .Y(n_361) );
AO21x2_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_210), .B(n_211), .Y(n_203) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_204), .A2(n_210), .B(n_211), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_209), .Y(n_204) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_210), .A2(n_213), .B(n_219), .Y(n_212) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_210), .A2(n_213), .B(n_219), .Y(n_259) );
AO21x1_ASAP7_75t_SL g460 ( .A1(n_210), .A2(n_461), .B(n_467), .Y(n_460) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_210), .A2(n_461), .B(n_467), .Y(n_536) );
INVx2_ASAP7_75t_L g270 ( .A(n_212), .Y(n_270) );
AND2x2_ASAP7_75t_L g319 ( .A(n_212), .B(n_233), .Y(n_319) );
AND2x2_ASAP7_75t_L g363 ( .A(n_212), .B(n_272), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_214), .B(n_218), .Y(n_213) );
AND2x2_ASAP7_75t_L g248 ( .A(n_221), .B(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_221), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_SL g442 ( .A(n_221), .B(n_277), .Y(n_442) );
INVx4_ASAP7_75t_L g247 ( .A(n_222), .Y(n_247) );
AND2x2_ASAP7_75t_L g279 ( .A(n_222), .B(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_222), .Y(n_332) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_229), .B(n_230), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_228), .Y(n_223) );
AOI21x1_ASAP7_75t_L g491 ( .A1(n_229), .A2(n_492), .B(n_498), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g341 ( .A(n_231), .B(n_316), .Y(n_341) );
INVx1_ASAP7_75t_SL g380 ( .A(n_231), .Y(n_380) );
AND2x4_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
AND2x4_ASAP7_75t_L g271 ( .A(n_232), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_232), .B(n_270), .Y(n_339) );
AND2x2_ASAP7_75t_L g391 ( .A(n_232), .B(n_241), .Y(n_391) );
OR2x2_ASAP7_75t_L g415 ( .A(n_232), .B(n_233), .Y(n_415) );
AND2x2_ASAP7_75t_L g239 ( .A(n_233), .B(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g289 ( .A(n_233), .B(n_270), .Y(n_289) );
AND2x2_ASAP7_75t_SL g345 ( .A(n_233), .B(n_257), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_239), .B(n_352), .Y(n_369) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
BUFx2_ASAP7_75t_L g304 ( .A(n_241), .Y(n_304) );
AND2x4_ASAP7_75t_SL g344 ( .A(n_241), .B(n_258), .Y(n_344) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_245), .Y(n_242) );
OR2x2_ASAP7_75t_L g292 ( .A(n_243), .B(n_246), .Y(n_292) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g261 ( .A(n_244), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g409 ( .A(n_244), .B(n_322), .Y(n_409) );
AND2x2_ASAP7_75t_L g425 ( .A(n_244), .B(n_279), .Y(n_425) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AOI311xp33_ASAP7_75t_L g395 ( .A1(n_246), .A2(n_334), .A3(n_396), .B(n_398), .C(n_405), .Y(n_395) );
AND2x4_ASAP7_75t_L g262 ( .A(n_247), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g266 ( .A(n_247), .Y(n_266) );
NAND2x1p5_ASAP7_75t_L g336 ( .A(n_247), .B(n_280), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_247), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g379 ( .A(n_247), .B(n_366), .Y(n_379) );
AND2x2_ASAP7_75t_L g265 ( .A(n_249), .B(n_266), .Y(n_265) );
INVxp67_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
INVxp67_ASAP7_75t_SL g283 ( .A(n_250), .Y(n_283) );
OR2x2_ASAP7_75t_L g372 ( .A(n_250), .B(n_336), .Y(n_372) );
INVx1_ASAP7_75t_L g428 ( .A(n_250), .Y(n_428) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_256), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g337 ( .A(n_254), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g351 ( .A(n_254), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g426 ( .A(n_254), .B(n_299), .Y(n_426) );
BUFx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g269 ( .A(n_255), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g288 ( .A(n_255), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g350 ( .A(n_256), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_256), .A2(n_406), .B1(n_407), .B2(n_408), .Y(n_405) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
AND2x2_ASAP7_75t_L g299 ( .A(n_257), .B(n_270), .Y(n_299) );
AND2x4_ASAP7_75t_L g352 ( .A(n_257), .B(n_259), .Y(n_352) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OAI21xp33_ASAP7_75t_SL g260 ( .A1(n_261), .A2(n_265), .B(n_267), .Y(n_260) );
AOI22xp5_ASAP7_75t_L g346 ( .A1(n_261), .A2(n_347), .B1(n_351), .B2(n_353), .Y(n_346) );
AND2x2_ASAP7_75t_SL g306 ( .A(n_262), .B(n_280), .Y(n_306) );
INVx2_ASAP7_75t_L g368 ( .A(n_262), .Y(n_368) );
AND2x2_ASAP7_75t_L g382 ( .A(n_262), .B(n_378), .Y(n_382) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g278 ( .A(n_264), .Y(n_278) );
INVx1_ASAP7_75t_L g331 ( .A(n_264), .Y(n_331) );
INVx1_ASAP7_75t_L g282 ( .A(n_266), .Y(n_282) );
AND3x2_ASAP7_75t_L g310 ( .A(n_266), .B(n_311), .C(n_312), .Y(n_310) );
INVx1_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
INVx1_ASAP7_75t_L g374 ( .A(n_269), .Y(n_374) );
AND2x2_ASAP7_75t_L g302 ( .A(n_271), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g373 ( .A(n_271), .B(n_374), .Y(n_373) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_271), .A2(n_385), .B1(n_389), .B2(n_392), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_271), .B(n_419), .Y(n_423) );
BUFx2_ASAP7_75t_L g314 ( .A(n_272), .Y(n_314) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g285 ( .A(n_273), .Y(n_285) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_273), .Y(n_404) );
OAI221xp5_ASAP7_75t_SL g274 ( .A1(n_275), .A2(n_284), .B1(n_286), .B2(n_287), .C(n_290), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_276), .B(n_281), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
INVx1_ASAP7_75t_L g366 ( .A(n_278), .Y(n_366) );
INVx2_ASAP7_75t_SL g355 ( .A(n_279), .Y(n_355) );
AND2x2_ASAP7_75t_L g437 ( .A(n_279), .B(n_304), .Y(n_437) );
INVx4_ASAP7_75t_L g328 ( .A(n_280), .Y(n_328) );
INVx1_ASAP7_75t_L g286 ( .A(n_281), .Y(n_286) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x4_ASAP7_75t_L g397 ( .A(n_285), .B(n_352), .Y(n_397) );
INVx1_ASAP7_75t_SL g436 ( .A(n_285), .Y(n_436) );
AND2x2_ASAP7_75t_L g441 ( .A(n_285), .B(n_344), .Y(n_441) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g383 ( .A(n_289), .Y(n_383) );
OAI21xp5_ASAP7_75t_SL g290 ( .A1(n_291), .A2(n_293), .B(n_295), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx1_ASAP7_75t_L g316 ( .A(n_297), .Y(n_316) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g313 ( .A(n_299), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g403 ( .A(n_299), .B(n_404), .Y(n_403) );
OAI211xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_305), .B(n_307), .C(n_324), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g396 ( .A(n_303), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_304), .B(n_319), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_304), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g429 ( .A(n_304), .B(n_352), .Y(n_429) );
OAI221xp5_ASAP7_75t_SL g340 ( .A1(n_305), .A2(n_329), .B1(n_341), .B2(n_342), .C(n_346), .Y(n_340) );
INVx3_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g411 ( .A(n_306), .B(n_312), .Y(n_411) );
OAI32xp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_313), .A3(n_315), .B1(n_317), .B2(n_321), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVxp67_ASAP7_75t_SL g401 ( .A(n_311), .Y(n_401) );
INVx2_ASAP7_75t_L g334 ( .A(n_312), .Y(n_334) );
O2A1O1Ixp33_ASAP7_75t_L g443 ( .A1(n_312), .A2(n_364), .B(n_444), .C(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g349 ( .A(n_314), .Y(n_349) );
OR2x2_ASAP7_75t_L g445 ( .A(n_314), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_318), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g406 ( .A(n_321), .Y(n_406) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g387 ( .A(n_322), .Y(n_387) );
OAI21xp33_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_333), .B(n_337), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
OR2x2_ASAP7_75t_L g364 ( .A(n_327), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_328), .B(n_331), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_330), .A2(n_362), .B1(n_431), .B2(n_434), .C(n_438), .Y(n_430) );
INVx2_ASAP7_75t_L g433 ( .A(n_330), .Y(n_433) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
OR2x2_ASAP7_75t_L g354 ( .A(n_334), .B(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_L g421 ( .A(n_334), .B(n_379), .Y(n_421) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVxp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g419 ( .A(n_344), .Y(n_419) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_352), .B(n_382), .Y(n_439) );
INVx2_ASAP7_75t_L g446 ( .A(n_352), .Y(n_446) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_354), .A2(n_417), .B1(n_420), .B2(n_422), .C(n_424), .Y(n_416) );
AND5x1_ASAP7_75t_L g356 ( .A(n_357), .B(n_395), .C(n_410), .D(n_430), .E(n_440), .Y(n_356) );
NOR2xp33_ASAP7_75t_SL g357 ( .A(n_358), .B(n_375), .Y(n_357) );
OAI221xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_364), .B1(n_367), .B2(n_369), .C(n_370), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g359 ( .A(n_360), .B(n_362), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_373), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI221xp5_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_380), .B1(n_381), .B2(n_383), .C(n_384), .Y(n_375) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_380), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
OR2x2_ASAP7_75t_L g393 ( .A(n_388), .B(n_394), .Y(n_393) );
CKINVDCx16_ASAP7_75t_R g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
AOI21xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .B(n_402), .Y(n_398) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B(n_416), .Y(n_410) );
INVx1_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVxp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_427), .B2(n_429), .Y(n_424) );
O2A1O1Ixp33_ASAP7_75t_L g440 ( .A1(n_426), .A2(n_441), .B(n_442), .C(n_443), .Y(n_440) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx1_ASAP7_75t_L g444 ( .A(n_437), .Y(n_444) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx4_ASAP7_75t_L g762 ( .A(n_447), .Y(n_762) );
OAI22xp5_ASAP7_75t_SL g772 ( .A1(n_447), .A2(n_762), .B1(n_773), .B2(n_774), .Y(n_772) );
AND3x4_ASAP7_75t_L g447 ( .A(n_448), .B(n_634), .C(n_730), .Y(n_447) );
NOR3xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_576), .C(n_603), .Y(n_448) );
OAI211xp5_ASAP7_75t_SL g449 ( .A1(n_450), .A2(n_486), .B(n_525), .C(n_549), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_468), .Y(n_450) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_451), .A2(n_527), .B(n_531), .C(n_537), .Y(n_526) );
OR2x2_ASAP7_75t_L g649 ( .A(n_451), .B(n_586), .Y(n_649) );
INVx2_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g616 ( .A(n_452), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_452), .B(n_587), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_452), .B(n_732), .Y(n_747) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_460), .Y(n_452) );
AND2x2_ASAP7_75t_L g533 ( .A(n_453), .B(n_469), .Y(n_533) );
INVx1_ASAP7_75t_L g553 ( .A(n_453), .Y(n_553) );
OR2x2_ASAP7_75t_L g568 ( .A(n_453), .B(n_477), .Y(n_568) );
INVx2_ASAP7_75t_L g574 ( .A(n_453), .Y(n_574) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_453), .Y(n_629) );
INVx1_ASAP7_75t_L g706 ( .A(n_453), .Y(n_706) );
NOR2x1_ASAP7_75t_SL g555 ( .A(n_460), .B(n_477), .Y(n_555) );
AND2x2_ASAP7_75t_L g585 ( .A(n_460), .B(n_574), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_466), .Y(n_461) );
OR2x2_ASAP7_75t_L g579 ( .A(n_468), .B(n_580), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_468), .B(n_686), .Y(n_685) );
INVx3_ASAP7_75t_L g707 ( .A(n_468), .Y(n_707) );
NAND2x1_ASAP7_75t_L g468 ( .A(n_469), .B(n_477), .Y(n_468) );
OR2x2_ASAP7_75t_SL g567 ( .A(n_469), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g571 ( .A(n_469), .Y(n_571) );
INVx4_ASAP7_75t_L g587 ( .A(n_469), .Y(n_587) );
OR2x2_ASAP7_75t_L g602 ( .A(n_469), .B(n_535), .Y(n_602) );
AND2x2_ASAP7_75t_L g641 ( .A(n_469), .B(n_555), .Y(n_641) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_469), .Y(n_653) );
OR2x6_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
AND2x2_ASAP7_75t_L g534 ( .A(n_477), .B(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g586 ( .A(n_477), .B(n_587), .Y(n_586) );
BUFx2_ASAP7_75t_L g601 ( .A(n_477), .Y(n_601) );
AND2x2_ASAP7_75t_L g617 ( .A(n_477), .B(n_587), .Y(n_617) );
AND2x2_ASAP7_75t_L g630 ( .A(n_477), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g662 ( .A(n_477), .B(n_574), .Y(n_662) );
INVx2_ASAP7_75t_SL g732 ( .A(n_477), .Y(n_732) );
OR2x6_ASAP7_75t_L g477 ( .A(n_478), .B(n_485), .Y(n_477) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NOR2xp67_ASAP7_75t_L g487 ( .A(n_488), .B(n_507), .Y(n_487) );
OAI211xp5_ASAP7_75t_L g603 ( .A1(n_488), .A2(n_604), .B(n_608), .C(n_624), .Y(n_603) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g699 ( .A(n_489), .B(n_538), .Y(n_699) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_499), .Y(n_489) );
INVx2_ASAP7_75t_L g548 ( .A(n_490), .Y(n_548) );
AND2x4_ASAP7_75t_SL g559 ( .A(n_490), .B(n_539), .Y(n_559) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_490), .Y(n_563) );
AND2x2_ASAP7_75t_L g621 ( .A(n_490), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g695 ( .A(n_490), .Y(n_695) );
INVx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_491), .Y(n_597) );
AND2x2_ASAP7_75t_L g640 ( .A(n_491), .B(n_499), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_497), .Y(n_492) );
INVx2_ASAP7_75t_L g530 ( .A(n_499), .Y(n_530) );
AND2x2_ASAP7_75t_L g590 ( .A(n_499), .B(n_539), .Y(n_590) );
INVx2_ASAP7_75t_L g622 ( .A(n_499), .Y(n_622) );
OR2x2_ASAP7_75t_L g645 ( .A(n_499), .B(n_510), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_505), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_507), .B(n_562), .Y(n_669) );
AND2x2_ASAP7_75t_L g703 ( .A(n_507), .B(n_639), .Y(n_703) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OAI31xp33_ASAP7_75t_SL g624 ( .A1(n_508), .A2(n_605), .A3(n_625), .B(n_632), .Y(n_624) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_509), .B(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
BUFx3_ASAP7_75t_L g558 ( .A(n_510), .Y(n_558) );
AND2x2_ASAP7_75t_L g575 ( .A(n_510), .B(n_538), .Y(n_575) );
AND2x4_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
AND2x4_ASAP7_75t_L g565 ( .A(n_511), .B(n_512), .Y(n_565) );
AND2x4_ASAP7_75t_L g514 ( .A(n_515), .B(n_518), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
NOR2x1p5_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g710 ( .A(n_528), .Y(n_710) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NOR2x1_ASAP7_75t_L g592 ( .A(n_530), .B(n_539), .Y(n_592) );
AND2x2_ASAP7_75t_L g633 ( .A(n_530), .B(n_548), .Y(n_633) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
AND2x2_ASAP7_75t_L g613 ( .A(n_534), .B(n_571), .Y(n_613) );
AND2x2_ASAP7_75t_L g572 ( .A(n_535), .B(n_573), .Y(n_572) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_535), .Y(n_581) );
INVx2_ASAP7_75t_L g631 ( .A(n_535), .Y(n_631) );
AND2x2_ASAP7_75t_L g721 ( .A(n_535), .B(n_706), .Y(n_721) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g727 ( .A(n_537), .Y(n_727) );
NAND2x1p5_ASAP7_75t_L g537 ( .A(n_538), .B(n_547), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_538), .B(n_597), .Y(n_666) );
AND2x2_ASAP7_75t_L g714 ( .A(n_538), .B(n_640), .Y(n_714) );
INVx4_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g623 ( .A(n_539), .B(n_595), .Y(n_623) );
AND2x2_ASAP7_75t_L g632 ( .A(n_539), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g644 ( .A(n_539), .Y(n_644) );
BUFx2_ASAP7_75t_L g660 ( .A(n_539), .Y(n_660) );
AND2x4_ASAP7_75t_L g694 ( .A(n_539), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g739 ( .A(n_539), .B(n_640), .Y(n_739) );
OR2x6_ASAP7_75t_L g539 ( .A(n_540), .B(n_546), .Y(n_539) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
AOI222xp33_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_556), .B1(n_560), .B2(n_566), .C1(n_569), .C2(n_575), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_551), .A2(n_615), .B1(n_618), .B2(n_623), .Y(n_614) );
OR2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_554), .Y(n_551) );
AND2x2_ASAP7_75t_L g598 ( .A(n_552), .B(n_599), .Y(n_598) );
AND2x4_ASAP7_75t_SL g612 ( .A(n_552), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_552), .B(n_617), .Y(n_750) );
INVx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g711 ( .A(n_553), .B(n_617), .Y(n_711) );
OR2x2_ASAP7_75t_L g688 ( .A(n_554), .B(n_570), .Y(n_688) );
OR2x2_ASAP7_75t_L g696 ( .A(n_554), .B(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g680 ( .A(n_555), .B(n_573), .Y(n_680) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
OR2x2_ASAP7_75t_L g588 ( .A(n_558), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g738 ( .A(n_558), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g689 ( .A(n_559), .B(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_559), .B(n_718), .Y(n_717) );
INVx2_ASAP7_75t_SL g724 ( .A(n_559), .Y(n_724) );
INVxp67_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
INVx2_ASAP7_75t_L g709 ( .A(n_562), .Y(n_709) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g611 ( .A(n_563), .B(n_590), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_564), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g610 ( .A(n_564), .Y(n_610) );
NOR2x1_ASAP7_75t_L g619 ( .A(n_564), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g713 ( .A(n_564), .B(n_585), .Y(n_713) );
INVx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g647 ( .A(n_565), .B(n_633), .Y(n_647) );
AND2x2_ASAP7_75t_L g690 ( .A(n_565), .B(n_622), .Y(n_690) );
AND2x4_ASAP7_75t_L g605 ( .A(n_566), .B(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g746 ( .A(n_568), .B(n_602), .Y(n_746) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_570), .B(n_585), .Y(n_729) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_571), .B(n_585), .Y(n_651) );
A2O1A1Ixp33_ASAP7_75t_L g712 ( .A1(n_571), .A2(n_612), .B(n_713), .C(n_714), .Y(n_712) );
AND2x2_ASAP7_75t_L g743 ( .A(n_571), .B(n_721), .Y(n_743) );
INVx1_ASAP7_75t_L g654 ( .A(n_572), .Y(n_654) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_575), .B(n_639), .Y(n_638) );
OAI21xp33_ASAP7_75t_SL g576 ( .A1(n_577), .A2(n_588), .B(n_591), .Y(n_576) );
NOR2x1_ASAP7_75t_L g577 ( .A(n_578), .B(n_582), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_579), .A2(n_732), .B1(n_733), .B2(n_735), .Y(n_731) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g607 ( .A(n_581), .Y(n_607) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NOR2xp67_ASAP7_75t_L g628 ( .A(n_587), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g679 ( .A(n_587), .Y(n_679) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OAI21xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B(n_598), .Y(n_591) );
INVx1_ASAP7_75t_L g670 ( .A(n_592), .Y(n_670) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx2_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_612), .B(n_614), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
OR2x2_ASAP7_75t_L g655 ( .A(n_610), .B(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g692 ( .A(n_610), .B(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_610), .B(n_640), .Y(n_728) );
INVx1_ASAP7_75t_L g748 ( .A(n_611), .Y(n_748) );
AOI221xp5_ASAP7_75t_L g715 ( .A1(n_613), .A2(n_716), .B1(n_719), .B2(n_722), .C(n_725), .Y(n_715) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OAI321xp33_ASAP7_75t_L g736 ( .A1(n_618), .A2(n_653), .A3(n_737), .B1(n_740), .B2(n_742), .C(n_744), .Y(n_736) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g677 ( .A(n_622), .Y(n_677) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g671 ( .A(n_627), .Y(n_671) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
INVx1_ASAP7_75t_L g697 ( .A(n_628), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_630), .A2(n_658), .B1(n_662), .B2(n_663), .C(n_668), .Y(n_657) );
INVxp67_ASAP7_75t_L g686 ( .A(n_631), .Y(n_686) );
INVx1_ASAP7_75t_L g656 ( .A(n_633), .Y(n_656) );
NOR2xp67_ASAP7_75t_L g634 ( .A(n_635), .B(n_681), .Y(n_634) );
NAND3xp33_ASAP7_75t_L g635 ( .A(n_636), .B(n_657), .C(n_672), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_641), .B1(n_642), .B2(n_648), .C(n_650), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
BUFx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g755 ( .A(n_640), .Y(n_755) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_643), .B(n_646), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g735 ( .A(n_644), .B(n_690), .Y(n_735) );
INVx2_ASAP7_75t_SL g667 ( .A(n_645), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_646), .A2(n_651), .B1(n_652), .B2(n_655), .Y(n_650) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_654), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_655), .B(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g661 ( .A(n_656), .Y(n_661) );
AOI222xp33_ASAP7_75t_L g700 ( .A1(n_658), .A2(n_701), .B1(n_703), .B2(n_704), .C1(n_708), .C2(n_711), .Y(n_700) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_659), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g734 ( .A(n_659), .B(n_713), .Y(n_734) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_667), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_667), .B(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_667), .B(n_727), .Y(n_726) );
AOI21xp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B(n_671), .Y(n_668) );
NAND2xp33_ASAP7_75t_SL g672 ( .A(n_673), .B(n_678), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
BUFx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_678), .B(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
NAND4xp25_ASAP7_75t_SL g681 ( .A(n_682), .B(n_700), .C(n_712), .D(n_715), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_687), .B(n_689), .C(n_691), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_688), .A2(n_692), .B1(n_696), .B2(n_698), .Y(n_691) );
INVx1_ASAP7_75t_L g718 ( .A(n_690), .Y(n_718) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_707), .Y(n_704) );
BUFx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_707), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVxp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVxp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_724), .A2(n_746), .B1(n_747), .B2(n_748), .Y(n_745) );
AOI21xp33_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_728), .B(n_729), .Y(n_725) );
NOR4xp25_ASAP7_75t_L g730 ( .A(n_731), .B(n_736), .C(n_749), .D(n_751), .Y(n_730) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx4_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx3_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
OAI22x1_ASAP7_75t_L g761 ( .A1(n_758), .A2(n_762), .B1(n_763), .B2(n_764), .Y(n_761) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_759), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
BUFx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_SL g778 ( .A(n_779), .Y(n_778) );
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_780), .Y(n_789) );
AND2x4_ASAP7_75t_SL g780 ( .A(n_781), .B(n_782), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
endmodule