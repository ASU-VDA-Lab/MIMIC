module real_jpeg_12652_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_323;
wire n_176;
wire n_166;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g88 ( 
.A(n_0),
.Y(n_88)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_41),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_3),
.A2(n_30),
.B(n_36),
.C(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_3),
.B(n_45),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_3),
.B(n_31),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_SL g158 ( 
.A1(n_3),
.A2(n_31),
.B(n_143),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_3),
.B(n_65),
.C(n_70),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_3),
.A2(n_41),
.B1(n_50),
.B2(n_54),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_3),
.A2(n_86),
.B1(n_87),
.B2(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_3),
.B(n_114),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_57),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_5),
.A2(n_50),
.B1(n_54),
.B2(n_57),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_5),
.A2(n_57),
.B1(n_69),
.B2(n_70),
.Y(n_173)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_7),
.A2(n_69),
.B1(n_70),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_7),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_7),
.A2(n_50),
.B1(n_54),
.B2(n_90),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_90),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_7),
.A2(n_36),
.B1(n_37),
.B2(n_90),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_8),
.A2(n_69),
.B1(n_70),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_8),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_8),
.A2(n_50),
.B1(n_54),
.B2(n_92),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_92),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_8),
.A2(n_36),
.B1(n_37),
.B2(n_92),
.Y(n_307)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_10),
.A2(n_50),
.B1(n_54),
.B2(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_75),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_10),
.A2(n_69),
.B1(n_70),
.B2(n_75),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_75),
.Y(n_253)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_13),
.A2(n_50),
.B1(n_54),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_13),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_13),
.A2(n_69),
.B1(n_70),
.B2(n_78),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_78),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_78),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_14),
.A2(n_36),
.B1(n_37),
.B2(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_44),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_14),
.A2(n_44),
.B1(n_50),
.B2(n_54),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_14),
.A2(n_44),
.B1(n_69),
.B2(n_70),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_15),
.A2(n_50),
.B1(n_54),
.B2(n_59),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_15),
.A2(n_59),
.B1(n_69),
.B2(n_70),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_15),
.A2(n_36),
.B1(n_37),
.B2(n_59),
.Y(n_224)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_323),
.C(n_327),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_321),
.B(n_325),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_314),
.B(n_320),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_280),
.B(n_311),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_258),
.B(n_279),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_231),
.B(n_257),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_126),
.B(n_207),
.C(n_230),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_105),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_24),
.B(n_105),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_81),
.C(n_96),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_25),
.B(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_46),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_26),
.B(n_60),
.C(n_80),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_40),
.B1(n_42),
.B2(n_45),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_27),
.B(n_276),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_27),
.A2(n_45),
.B(n_253),
.Y(n_327)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_28),
.A2(n_29),
.B1(n_43),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_28),
.A2(n_29),
.B1(n_109),
.B2(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_28),
.A2(n_224),
.B(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_28),
.A2(n_274),
.B(n_275),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_28),
.A2(n_29),
.B1(n_292),
.B2(n_307),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_28),
.A2(n_275),
.B(n_307),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_29),
.A2(n_292),
.B(n_293),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_30),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_31),
.A2(n_32),
.B1(n_52),
.B2(n_53),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_L g95 ( 
.A1(n_31),
.A2(n_34),
.B(n_41),
.Y(n_95)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND3xp33_ASAP7_75t_SL g144 ( 
.A(n_32),
.B(n_52),
.C(n_54),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_41),
.B(n_87),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_41),
.B(n_68),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_45),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_45),
.B(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_60),
.B1(n_61),
.B2(n_80),
.Y(n_46)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_56),
.B2(n_58),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_48),
.A2(n_49),
.B1(n_56),
.B2(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_48),
.A2(n_58),
.B(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_48),
.A2(n_49),
.B1(n_104),
.B2(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_48),
.A2(n_113),
.B(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_48),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_48),
.A2(n_226),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_55),
.Y(n_48)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_49),
.A2(n_248),
.B(n_249),
.Y(n_247)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g54 ( 
.A(n_50),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_54),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_50),
.A2(n_53),
.B(n_142),
.C(n_144),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_50),
.B(n_167),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_73),
.B(n_76),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_62),
.A2(n_136),
.B(n_138),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_62),
.A2(n_68),
.B(n_73),
.Y(n_289)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_63),
.B(n_77),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_63),
.A2(n_79),
.B1(n_137),
.B2(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_63),
.A2(n_79),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_63),
.A2(n_79),
.B1(n_160),
.B2(n_170),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_63),
.A2(n_79),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_63),
.A2(n_217),
.B(n_241),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_68),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_69),
.B(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_87),
.Y(n_86)
);

BUFx4f_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_74),
.B(n_79),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_76),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_81),
.A2(n_82),
.B1(n_96),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_93),
.B2(n_94),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_93),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_88),
.B1(n_89),
.B2(n_91),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_85),
.A2(n_124),
.B(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_85),
.A2(n_88),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_86),
.A2(n_87),
.B1(n_173),
.B2(n_181),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_86),
.A2(n_175),
.B(n_191),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_86),
.A2(n_87),
.B(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_100),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_89),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_88),
.B(n_147),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_91),
.Y(n_122)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.C(n_103),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_102),
.Y(n_134)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_99),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_103),
.B(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_116),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_106),
.B(n_117),
.C(n_125),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_115),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_108),
.B(n_110),
.C(n_115),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_111),
.B(n_249),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_112),
.A2(n_114),
.B(n_250),
.Y(n_317)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_114),
.B(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_114),
.A2(n_250),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_125),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_118),
.B(n_121),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_119),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_120),
.B(n_138),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_205),
.B(n_206),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_148),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_132),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_129),
.B(n_132),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.C(n_139),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_135),
.A2(n_139),
.B1(n_140),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_145),
.B1(n_146),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_147),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_161),
.B(n_204),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_150),
.B(n_153),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.C(n_159),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_154),
.B(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_156),
.A2(n_157),
.B1(n_159),
.B2(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_198),
.B(n_203),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_187),
.B(n_197),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_176),
.B(n_186),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_171),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_171),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_168),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_182),
.B(n_185),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_184),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_189),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_193),
.C(n_196),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_191),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_202),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_229),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_229),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_211),
.C(n_219),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_219),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_218),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_218),
.Y(n_244)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_222),
.C(n_228),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_225),
.B2(n_228),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_225),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_227),
.B(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_233),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_256),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_242),
.B1(n_254),
.B2(n_255),
.Y(n_234)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_235),
.B(n_255),
.C(n_256),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_236),
.A2(n_237),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_239),
.Y(n_270)
);

AOI21xp33_ASAP7_75t_L g295 ( 
.A1(n_237),
.A2(n_270),
.B(n_272),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_247),
.C(n_251),
.Y(n_261)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_248),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_252),
.B(n_293),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_278),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_278),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_277),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_260),
.B(n_263),
.C(n_269),
.Y(n_309)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_269),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_267),
.B(n_268),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_264),
.B(n_267),
.Y(n_268)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_283),
.C(n_295),
.Y(n_282)
);

FAx1_ASAP7_75t_SL g310 ( 
.A(n_268),
.B(n_283),
.CI(n_295),
.CON(n_310),
.SN(n_310)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_308),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g311 ( 
.A1(n_281),
.A2(n_312),
.B(n_313),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_296),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_282),
.B(n_296),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_291),
.B2(n_294),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_289),
.B2(n_290),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_290),
.C(n_291),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_289),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_290),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_289),
.B(n_303),
.C(n_305),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_291),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_291),
.A2(n_294),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_297),
.C(n_300),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_305),
.B2(n_306),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_310),
.Y(n_312)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_310),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_316),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_316),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_323),
.Y(n_326)
);

FAx1_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_318),
.CI(n_319),
.CON(n_316),
.SN(n_316)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_323),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);


endmodule