module real_jpeg_13849_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_273, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_273;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

BUFx10_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_2),
.A2(n_48),
.B1(n_62),
.B2(n_64),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_48),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_2),
.A2(n_31),
.B1(n_33),
.B2(n_48),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_3),
.A2(n_31),
.B1(n_33),
.B2(n_56),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_3),
.A2(n_35),
.B1(n_36),
.B2(n_56),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_3),
.A2(n_56),
.B1(n_62),
.B2(n_64),
.Y(n_154)
);

BUFx16f_ASAP7_75t_L g76 ( 
.A(n_4),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_8),
.A2(n_45),
.B1(n_46),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_8),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_99),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_8),
.A2(n_62),
.B1(n_64),
.B2(n_99),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_8),
.A2(n_31),
.B1(n_33),
.B2(n_99),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_9),
.A2(n_62),
.B1(n_64),
.B2(n_80),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_9),
.A2(n_31),
.B1(n_33),
.B2(n_80),
.Y(n_111)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_11),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_11),
.B(n_62),
.C(n_76),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_11),
.B(n_34),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_11),
.A2(n_65),
.B(n_153),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_11),
.A2(n_32),
.B(n_33),
.C(n_180),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_11),
.A2(n_31),
.B1(n_33),
.B2(n_138),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_11),
.B(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_11),
.B(n_45),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_12),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_61),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_13),
.A2(n_31),
.B1(n_33),
.B2(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_51),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_SL g235 ( 
.A(n_13),
.B(n_31),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_14),
.A2(n_62),
.B1(n_64),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_14),
.A2(n_35),
.B1(n_36),
.B2(n_69),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_15),
.A2(n_31),
.B1(n_33),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_15),
.A2(n_39),
.B1(n_45),
.B2(n_46),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_15),
.A2(n_39),
.B1(n_62),
.B2(n_64),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_16),
.A2(n_31),
.B1(n_33),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_16),
.A2(n_35),
.B1(n_36),
.B2(n_42),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_16),
.A2(n_42),
.B1(n_62),
.B2(n_64),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_126),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_103),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_21),
.B(n_103),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_83),
.C(n_91),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_22),
.A2(n_23),
.B1(n_83),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_57),
.B2(n_82),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_43),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_26),
.B(n_43),
.C(n_82),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_27),
.A2(n_40),
.B1(n_41),
.B2(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_27),
.A2(n_185),
.B(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_27),
.A2(n_40),
.B1(n_199),
.B2(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_27),
.A2(n_186),
.B(n_226),
.Y(n_246)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_28),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_34),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_29)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

AO22x1_ASAP7_75t_SL g34 ( 
.A1(n_30),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_30),
.A2(n_35),
.B(n_138),
.Y(n_180)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

AOI32xp33_ASAP7_75t_L g234 ( 
.A1(n_33),
.A2(n_46),
.A3(n_51),
.B1(n_223),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_34),
.B(n_102),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_35),
.A2(n_36),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_36),
.B(n_142),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_38),
.A2(n_40),
.B(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_40),
.A2(n_101),
.B(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_49),
.B(n_53),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_44),
.A2(n_49),
.B1(n_50),
.B2(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_46),
.A2(n_49),
.B(n_138),
.C(n_222),
.Y(n_221)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_50),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_50),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_50),
.A2(n_98),
.B(n_120),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_54),
.B(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_71),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_58),
.A2(n_71),
.B1(n_72),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_58),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_65),
.B1(n_68),
.B2(n_70),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_66),
.B1(n_67),
.B2(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_64),
.B1(n_76),
.B2(n_77),
.Y(n_78)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_64),
.B(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_64),
.B(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_65),
.A2(n_152),
.B(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_65),
.A2(n_70),
.B1(n_182),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_65),
.A2(n_70),
.B1(n_206),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_67),
.B(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_66),
.A2(n_67),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_66),
.B(n_154),
.Y(n_167)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_67),
.B(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_70),
.A2(n_159),
.B(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_70),
.B(n_138),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_70),
.A2(n_167),
.B(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_79),
.B2(n_81),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_74),
.B1(n_81),
.B2(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_79),
.B1(n_81),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_74),
.B(n_140),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_74),
.A2(n_81),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_78),
.A2(n_89),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_78),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_78),
.B(n_138),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_78),
.A2(n_150),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_81),
.B(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_83),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_87),
.B2(n_90),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_84),
.A2(n_85),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_90),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_87),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_91),
.B(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_97),
.C(n_100),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_92),
.B(n_257),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_93),
.B(n_95),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_94),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_96),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_97),
.B(n_100),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_125),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_113),
.B2(n_114),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_110),
.B(n_112),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_110),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_137),
.B(n_139),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_108),
.A2(n_139),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_123),
.B2(n_124),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_266),
.B(n_271),
.Y(n_127)
);

OAI321xp33_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_240),
.A3(n_259),
.B1(n_264),
.B2(n_265),
.C(n_273),
.Y(n_128)
);

AOI21x1_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_215),
.B(n_239),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_193),
.B(n_214),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_175),
.B(n_192),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_155),
.B(n_174),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_143),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_134),
.B(n_143),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_141),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_136),
.B1(n_141),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_141),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_151),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_148),
.C(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_152),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_163),
.B(n_173),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_161),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_157),
.B(n_161),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_168),
.B(n_172),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_165),
.B(n_166),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_176),
.B(n_177),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_183),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_187),
.C(n_191),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_181),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_187),
.B1(n_190),
.B2(n_191),
.Y(n_183)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_184),
.Y(n_191)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_187),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_189),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_194),
.B(n_195),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_207),
.B2(n_208),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_210),
.C(n_212),
.Y(n_216)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_201),
.C(n_205),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_213),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_209),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_210),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_217),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_230),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_218),
.B(n_231),
.C(n_232),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_224),
.B2(n_229),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_225),
.C(n_227),
.Y(n_251)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_224),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_237),
.Y(n_249)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_252),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_252),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_250),
.C(n_251),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_242),
.A2(n_243),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_249),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_248),
.C(n_249),
.Y(n_258)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_247),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_250),
.B(n_251),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_258),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_256),
.C(n_258),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_260),
.B(n_261),
.Y(n_264)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_270),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_270),
.Y(n_271)
);


endmodule