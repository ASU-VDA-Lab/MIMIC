module fake_jpeg_21143_n_255 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_255);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_42),
.Y(n_49)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_23),
.B(n_31),
.C(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_23),
.B1(n_22),
.B2(n_33),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_50),
.B1(n_17),
.B2(n_18),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_33),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_SL g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_48),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_22),
.B1(n_23),
.B2(n_27),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_22),
.B1(n_28),
.B2(n_30),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_21),
.B1(n_18),
.B2(n_40),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_20),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_20),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_32),
.Y(n_57)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_69),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_61),
.A2(n_68),
.B(n_24),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_52),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_65),
.B(n_67),
.Y(n_90)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_32),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_40),
.B1(n_39),
.B2(n_27),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

INVxp33_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_77),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_29),
.B1(n_31),
.B2(n_17),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_46),
.B(n_29),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_79),
.B(n_82),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_53),
.B1(n_48),
.B2(n_43),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_84),
.B1(n_26),
.B2(n_19),
.Y(n_108)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_57),
.B(n_21),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_55),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_88),
.Y(n_91)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_54),
.A2(n_19),
.B1(n_25),
.B2(n_26),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_50),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_52),
.C(n_50),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_99),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_43),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_51),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_103),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_53),
.B1(n_58),
.B2(n_39),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_104),
.A2(n_108),
.B1(n_111),
.B2(n_74),
.Y(n_136)
);

AOI32xp33_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_19),
.A3(n_24),
.B1(n_58),
.B2(n_26),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_109),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_26),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_68),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_0),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_90),
.B(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_70),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_118),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_84),
.B(n_61),
.Y(n_117)
);

AOI322xp5_ASAP7_75t_L g164 ( 
.A1(n_117),
.A2(n_101),
.A3(n_15),
.B1(n_3),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_71),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_81),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_134),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_122),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_63),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_125),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_95),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_127),
.B(n_138),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_68),
.B1(n_77),
.B2(n_60),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_110),
.B1(n_100),
.B2(n_94),
.Y(n_154)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_66),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_16),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_141),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_136),
.A2(n_110),
.B1(n_86),
.B2(n_74),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_96),
.B(n_68),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_139),
.Y(n_152)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_75),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_93),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_140),
.B(n_115),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_98),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_62),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_101),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_129),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_144),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_116),
.Y(n_146)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_114),
.A3(n_92),
.B1(n_104),
.B2(n_97),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_126),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_130),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_151),
.A2(n_167),
.B(n_120),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_161),
.B1(n_162),
.B2(n_14),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_100),
.Y(n_155)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_94),
.Y(n_160)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_126),
.B1(n_133),
.B2(n_139),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_132),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_SL g172 ( 
.A1(n_163),
.A2(n_164),
.B(n_125),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_165),
.B(n_119),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_166),
.A2(n_141),
.B1(n_138),
.B2(n_124),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_0),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_121),
.B(n_127),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_171),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_179),
.B1(n_182),
.B2(n_184),
.Y(n_201)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_119),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_176),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_180),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_158),
.A2(n_133),
.B(n_127),
.Y(n_178)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_SL g179 ( 
.A1(n_145),
.A2(n_142),
.B(n_128),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_144),
.B(n_131),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_181),
.A2(n_186),
.B1(n_161),
.B2(n_154),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_158),
.A2(n_124),
.B1(n_3),
.B2(n_5),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_1),
.C(n_6),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_185),
.C(n_188),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_1),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_162),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_157),
.C(n_166),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_157),
.C(n_149),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_198),
.Y(n_209)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_187),
.Y(n_197)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_149),
.C(n_145),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_200),
.Y(n_210)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_206),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_153),
.C(n_150),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_183),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_185),
.A2(n_143),
.B1(n_151),
.B2(n_156),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_198),
.B(n_156),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_208),
.B(n_215),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_201),
.A2(n_195),
.B1(n_204),
.B2(n_193),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_211),
.A2(n_186),
.B1(n_169),
.B2(n_194),
.Y(n_225)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

OA21x2_ASAP7_75t_SL g215 ( 
.A1(n_190),
.A2(n_192),
.B(n_193),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_188),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_150),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_217),
.B(n_190),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_220),
.B(n_216),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_212),
.A2(n_203),
.B1(n_184),
.B2(n_205),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_221),
.A2(n_228),
.B(n_212),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_194),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_225),
.C(n_229),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_159),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_230),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_211),
.A2(n_159),
.B(n_153),
.Y(n_227)
);

NOR3xp33_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_210),
.C(n_213),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_173),
.C(n_168),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_207),
.Y(n_230)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_233),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_223),
.B(n_210),
.Y(n_234)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

OAI321xp33_ASAP7_75t_L g240 ( 
.A1(n_235),
.A2(n_238),
.A3(n_148),
.B1(n_167),
.B2(n_225),
.C(n_229),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_L g236 ( 
.A1(n_228),
.A2(n_213),
.B(n_219),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_236),
.A2(n_227),
.B1(n_221),
.B2(n_148),
.Y(n_239)
);

AOI31xp33_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_218),
.A3(n_214),
.B(n_168),
.Y(n_238)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_239),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_240),
.A2(n_242),
.B1(n_231),
.B2(n_12),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_235),
.A2(n_222),
.B(n_8),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_241),
.Y(n_245)
);

BUFx24_ASAP7_75t_SL g247 ( 
.A(n_243),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_248),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_245),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_250),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_252)
);

NOR4xp25_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_244),
.C(n_241),
.D(n_237),
.Y(n_251)
);

AO21x2_ASAP7_75t_L g253 ( 
.A1(n_251),
.A2(n_11),
.B(n_13),
.Y(n_253)
);

O2A1O1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_252),
.A2(n_253),
.B(n_249),
.C(n_13),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_254),
.B(n_14),
.Y(n_255)
);


endmodule