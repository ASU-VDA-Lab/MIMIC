module fake_jpeg_24703_n_242 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_33),
.B(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_27),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_31),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_25),
.B1(n_20),
.B2(n_19),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_46),
.A2(n_62),
.B1(n_22),
.B2(n_16),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_25),
.B1(n_20),
.B2(n_19),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_22),
.B1(n_16),
.B2(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_55),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_21),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_57),
.Y(n_67)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_63),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_21),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_20),
.B1(n_25),
.B2(n_22),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_22),
.B1(n_37),
.B2(n_21),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_60),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_25),
.B1(n_20),
.B2(n_19),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_33),
.B(n_26),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_21),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_32),
.B(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_66),
.A2(n_72),
.B1(n_75),
.B2(n_83),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_68),
.A2(n_71),
.B1(n_15),
.B2(n_28),
.Y(n_101)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_82),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_31),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_61),
.B1(n_44),
.B2(n_49),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_34),
.B1(n_36),
.B2(n_24),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_55),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_15),
.B(n_28),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_15),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_39),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_65),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_36),
.B1(n_34),
.B2(n_42),
.Y(n_83)
);

MAJx2_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_53),
.C(n_57),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_88),
.B(n_92),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_91),
.Y(n_112)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_14),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_76),
.Y(n_91)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_97),
.Y(n_123)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_45),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_100),
.Y(n_114)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_102),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_68),
.B1(n_85),
.B2(n_83),
.Y(n_120)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_103),
.Y(n_129)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_104),
.Y(n_124)
);

INVxp33_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_43),
.B1(n_50),
.B2(n_51),
.Y(n_118)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_108),
.Y(n_128)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_81),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_109),
.A2(n_130),
.B(n_56),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_99),
.A2(n_72),
.B1(n_61),
.B2(n_85),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_121),
.B1(n_48),
.B2(n_63),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_79),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_126),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_50),
.B1(n_51),
.B2(n_42),
.Y(n_142)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_119),
.B(n_122),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_26),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_102),
.A2(n_66),
.B1(n_43),
.B2(n_48),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_125),
.B(n_127),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_76),
.Y(n_126)
);

NAND2xp33_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_81),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_107),
.Y(n_131)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_134),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_112),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_133),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_115),
.B(n_88),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_86),
.C(n_99),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_143),
.C(n_114),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_90),
.A3(n_101),
.B1(n_70),
.B2(n_74),
.C1(n_80),
.C2(n_93),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_141),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_74),
.Y(n_138)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_124),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_142),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_140),
.A2(n_144),
.B1(n_120),
.B2(n_109),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_106),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_41),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_110),
.B1(n_127),
.B2(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_146),
.Y(n_158)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_149),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_124),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_150),
.Y(n_164)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_152),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_51),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_154),
.B(n_171),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_155),
.A2(n_160),
.B1(n_143),
.B2(n_137),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_147),
.A2(n_110),
.B(n_109),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_170),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_128),
.B1(n_114),
.B2(n_119),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_162),
.A2(n_151),
.B1(n_132),
.B2(n_137),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_169),
.C(n_41),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_126),
.Y(n_169)
);

INVx6_ASAP7_75t_SL g170 ( 
.A(n_139),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

BUFx12_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_133),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_175),
.B(n_186),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_173),
.A2(n_140),
.B1(n_149),
.B2(n_134),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_176),
.A2(n_178),
.B1(n_163),
.B2(n_161),
.Y(n_204)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_150),
.B1(n_145),
.B2(n_138),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_162),
.B(n_128),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_187),
.C(n_188),
.Y(n_197)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_183),
.Y(n_200)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_129),
.B1(n_106),
.B2(n_24),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_190),
.B1(n_168),
.B2(n_154),
.Y(n_192)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_1),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_189),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_170),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_41),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_50),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_29),
.B1(n_17),
.B2(n_31),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_172),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_194),
.C(n_199),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_192),
.A2(n_195),
.B1(n_204),
.B2(n_185),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_159),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_169),
.C(n_160),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_167),
.C(n_163),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_175),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_156),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_176),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_179),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_209),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_206),
.B(n_203),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_208),
.B(n_214),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_185),
.B1(n_29),
.B2(n_26),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_210),
.A2(n_198),
.B1(n_196),
.B2(n_30),
.Y(n_218)
);

O2A1O1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_29),
.B(n_42),
.C(n_27),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_211),
.A2(n_212),
.B(n_30),
.Y(n_221)
);

O2A1O1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_198),
.A2(n_42),
.B(n_27),
.C(n_38),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_41),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_215),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_201),
.Y(n_214)
);

BUFx24_ASAP7_75t_SL g215 ( 
.A(n_200),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_218),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_207),
.B(n_14),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_219),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_SL g220 ( 
.A1(n_211),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_221),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_222),
.A2(n_212),
.B(n_205),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_226),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_2),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_220),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_225),
.B(n_223),
.Y(n_230)
);

AOI322xp5_ASAP7_75t_L g235 ( 
.A1(n_230),
.A2(n_232),
.A3(n_233),
.B1(n_234),
.B2(n_229),
.C1(n_228),
.C2(n_7),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_38),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_224),
.B(n_27),
.Y(n_234)
);

AOI322xp5_ASAP7_75t_L g238 ( 
.A1(n_235),
.A2(n_237),
.A3(n_5),
.B1(n_6),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_231),
.A2(n_38),
.B(n_6),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_5),
.Y(n_239)
);

AOI322xp5_ASAP7_75t_L g237 ( 
.A1(n_230),
.A2(n_38),
.A3(n_27),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_5),
.Y(n_237)
);

AOI321xp33_ASAP7_75t_L g240 ( 
.A1(n_238),
.A2(n_239),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_240),
.A2(n_16),
.B(n_12),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_11),
.Y(n_242)
);


endmodule