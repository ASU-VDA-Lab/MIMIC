module fake_jpeg_17888_n_57 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_57);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_57;

wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx8_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_12),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_32),
.Y(n_35)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_39),
.B1(n_14),
.B2(n_24),
.Y(n_40)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_26),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_13),
.B1(n_23),
.B2(n_5),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_46),
.B1(n_47),
.B2(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_45),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_1),
.B1(n_3),
.B2(n_6),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_44),
.B1(n_16),
.B2(n_18),
.Y(n_52)
);

AOI21x1_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_44),
.B(n_41),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_53),
.A2(n_48),
.B1(n_42),
.B2(n_27),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_54),
.A2(n_48),
.B(n_27),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_56),
.A2(n_52),
.B1(n_15),
.B2(n_19),
.Y(n_57)
);


endmodule