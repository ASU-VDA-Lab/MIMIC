module fake_jpeg_4532_n_21 (n_0, n_3, n_2, n_1, n_21);

input n_0;
input n_3;
input n_2;
input n_1;

output n_21;

wire n_13;
wire n_10;
wire n_6;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_4;
wire n_16;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

BUFx5_ASAP7_75t_L g4 ( 
.A(n_2),
.Y(n_4)
);

INVx1_ASAP7_75t_L g5 ( 
.A(n_3),
.Y(n_5)
);

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_2),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_5),
.B(n_1),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_8),
.B(n_9),
.Y(n_12)
);

A2O1A1Ixp33_ASAP7_75t_L g9 ( 
.A1(n_6),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_9)
);

INVx13_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

AOI22xp5_ASAP7_75t_L g11 ( 
.A1(n_10),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_11)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_12),
.B(n_4),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_14),
.B(n_8),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_13),
.A2(n_11),
.B1(n_12),
.B2(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_16),
.B(n_14),
.Y(n_18)
);

AOI321xp33_ASAP7_75t_L g19 ( 
.A1(n_18),
.A2(n_15),
.A3(n_11),
.B1(n_1),
.B2(n_7),
.C(n_0),
.Y(n_19)
);

AOI322xp5_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_0),
.A3(n_7),
.B1(n_17),
.B2(n_14),
.C1(n_16),
.C2(n_12),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_20),
.B(n_17),
.CI(n_0),
.CON(n_21),
.SN(n_21)
);


endmodule