module fake_jpeg_1764_n_151 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_151);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_151;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx6_ASAP7_75t_SL g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_11),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_32),
.B(n_26),
.Y(n_78)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_17),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_37),
.Y(n_67)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_12),
.B(n_3),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_46),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_6),
.C(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_23),
.Y(n_55)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_14),
.A2(n_10),
.B1(n_13),
.B2(n_26),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_52),
.B(n_28),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_SL g45 ( 
.A(n_17),
.B(n_19),
.C(n_20),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_21),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_19),
.B(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_12),
.B(n_29),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_50),
.Y(n_75)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_13),
.A2(n_26),
.B1(n_22),
.B2(n_23),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_57),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_60),
.B(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_25),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_65),
.B(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_16),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_16),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_69),
.B(n_70),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_72),
.Y(n_91)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_84),
.B(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

OR2x4_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_52),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_30),
.C(n_44),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_93),
.C(n_94),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_16),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_88),
.B(n_90),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_16),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_66),
.B1(n_102),
.B2(n_83),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_62),
.A2(n_73),
.B1(n_54),
.B2(n_56),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_92),
.A2(n_66),
.B1(n_81),
.B2(n_84),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_77),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_58),
.B(n_56),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_99),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_79),
.B(n_74),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_74),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_101),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_66),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_104),
.B(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_63),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_86),
.B1(n_94),
.B2(n_98),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_85),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_98),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_106),
.B1(n_113),
.B2(n_121),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_115),
.B(n_87),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_111),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_87),
.C(n_105),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_126),
.C(n_107),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_114),
.B1(n_103),
.B2(n_118),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_125),
.A2(n_110),
.B1(n_116),
.B2(n_112),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_108),
.C(n_107),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_133),
.C(n_135),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_132),
.Y(n_137)
);

BUFx12_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_106),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_128),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_126),
.B(n_120),
.Y(n_139)
);

BUFx24_ASAP7_75t_SL g138 ( 
.A(n_130),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_138),
.B(n_130),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_129),
.C(n_136),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_142),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_127),
.B(n_134),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_144),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_127),
.C(n_134),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_146),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_148),
.A2(n_145),
.B(n_149),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_147),
.Y(n_151)
);


endmodule