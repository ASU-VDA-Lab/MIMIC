module fake_aes_8789_n_625 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_625);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_625;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_476;
wire n_227;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g73 ( .A(n_35), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_40), .Y(n_74) );
BUFx3_ASAP7_75t_L g75 ( .A(n_9), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_42), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_39), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_12), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_21), .Y(n_79) );
BUFx3_ASAP7_75t_L g80 ( .A(n_48), .Y(n_80) );
BUFx6f_ASAP7_75t_L g81 ( .A(n_10), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_36), .Y(n_82) );
CKINVDCx16_ASAP7_75t_R g83 ( .A(n_44), .Y(n_83) );
CKINVDCx16_ASAP7_75t_R g84 ( .A(n_19), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_58), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_24), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_43), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_53), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_21), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_61), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_28), .Y(n_91) );
CKINVDCx16_ASAP7_75t_R g92 ( .A(n_2), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_26), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_59), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_71), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_7), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_37), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_0), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_56), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_49), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_5), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_63), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_32), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_47), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_1), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_22), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_10), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_30), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_8), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_13), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_51), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_15), .Y(n_113) );
INVxp33_ASAP7_75t_SL g114 ( .A(n_6), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_46), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_45), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_15), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_19), .Y(n_118) );
INVxp33_ASAP7_75t_SL g119 ( .A(n_57), .Y(n_119) );
INVxp33_ASAP7_75t_SL g120 ( .A(n_20), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_25), .Y(n_121) );
OA21x2_ASAP7_75t_L g122 ( .A1(n_73), .A2(n_31), .B(n_70), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_73), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_84), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_108), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_92), .B(n_0), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_78), .B(n_1), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_116), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_83), .Y(n_129) );
INVxp67_ASAP7_75t_L g130 ( .A(n_75), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_118), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_74), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_81), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_99), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_78), .Y(n_135) );
CKINVDCx11_ASAP7_75t_R g136 ( .A(n_102), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_89), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_104), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_89), .B(n_3), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_74), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_76), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_76), .Y(n_142) );
NOR2xp33_ASAP7_75t_R g143 ( .A(n_104), .B(n_33), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_85), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_119), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_116), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_81), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_116), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_119), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_101), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_116), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_85), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_101), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_113), .B(n_3), .Y(n_154) );
NOR2xp33_ASAP7_75t_R g155 ( .A(n_113), .B(n_34), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_116), .Y(n_156) );
NOR2xp33_ASAP7_75t_R g157 ( .A(n_80), .B(n_38), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_86), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_86), .Y(n_159) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_88), .A2(n_29), .B(n_69), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_114), .Y(n_161) );
INVx4_ASAP7_75t_L g162 ( .A(n_80), .Y(n_162) );
CKINVDCx16_ASAP7_75t_R g163 ( .A(n_75), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_114), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_98), .B(n_4), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_130), .B(n_98), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_165), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_128), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_128), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_165), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_165), .Y(n_171) );
BUFx2_ASAP7_75t_L g172 ( .A(n_150), .Y(n_172) );
NOR2x1p5_ASAP7_75t_L g173 ( .A(n_153), .B(n_129), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_165), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_128), .Y(n_175) );
INVx4_ASAP7_75t_L g176 ( .A(n_162), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_163), .B(n_120), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_163), .B(n_120), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_161), .A2(n_164), .B1(n_149), .B2(n_145), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_162), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_123), .B(n_117), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_123), .B(n_117), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_162), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_128), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_128), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_162), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_128), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_132), .B(n_96), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_138), .B(n_77), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_133), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_122), .Y(n_191) );
NAND3x1_ASAP7_75t_L g192 ( .A(n_126), .B(n_79), .C(n_105), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_133), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_151), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_122), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_132), .B(n_93), .Y(n_196) );
AND2x6_ASAP7_75t_L g197 ( .A(n_140), .B(n_121), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_151), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_133), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_133), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_147), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_147), .Y(n_202) );
NAND3xp33_ASAP7_75t_L g203 ( .A(n_140), .B(n_121), .C(n_115), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_151), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_142), .B(n_106), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_142), .B(n_94), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_147), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_144), .B(n_107), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_122), .Y(n_209) );
BUFx3_ASAP7_75t_L g210 ( .A(n_122), .Y(n_210) );
INVx4_ASAP7_75t_L g211 ( .A(n_160), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_160), .Y(n_212) );
AND2x6_ASAP7_75t_L g213 ( .A(n_144), .B(n_115), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_159), .B(n_110), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_147), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_151), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_134), .B(n_112), .Y(n_217) );
OAI22xp33_ASAP7_75t_L g218 ( .A1(n_135), .A2(n_111), .B1(n_109), .B2(n_81), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_151), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_159), .B(n_103), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_151), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_156), .Y(n_222) );
AO22x2_ASAP7_75t_L g223 ( .A1(n_141), .A2(n_90), .B1(n_97), .B2(n_88), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_141), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_152), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_152), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_156), .Y(n_227) );
NAND3x1_ASAP7_75t_L g228 ( .A(n_127), .B(n_97), .C(n_91), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_158), .B(n_100), .Y(n_229) );
BUFx3_ASAP7_75t_L g230 ( .A(n_160), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_156), .Y(n_231) );
BUFx2_ASAP7_75t_L g232 ( .A(n_172), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_188), .B(n_158), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_224), .Y(n_234) );
NOR3xp33_ASAP7_75t_SL g235 ( .A(n_218), .B(n_125), .C(n_154), .Y(n_235) );
NOR3xp33_ASAP7_75t_SL g236 ( .A(n_177), .B(n_139), .C(n_87), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_182), .B(n_95), .Y(n_237) );
NOR2xp33_ASAP7_75t_R g238 ( .A(n_172), .B(n_136), .Y(n_238) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_223), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_188), .B(n_143), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_224), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_225), .Y(n_242) );
NOR3xp33_ASAP7_75t_SL g243 ( .A(n_178), .B(n_82), .C(n_90), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_192), .A2(n_228), .B1(n_217), .B2(n_167), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_225), .Y(n_245) );
NOR3xp33_ASAP7_75t_SL g246 ( .A(n_189), .B(n_91), .C(n_124), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_226), .Y(n_247) );
BUFx3_ASAP7_75t_L g248 ( .A(n_197), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_182), .B(n_157), .Y(n_249) );
NAND2x1p5_ASAP7_75t_L g250 ( .A(n_182), .B(n_81), .Y(n_250) );
INVx4_ASAP7_75t_L g251 ( .A(n_176), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_223), .A2(n_81), .B1(n_155), .B2(n_137), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_226), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_188), .B(n_160), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_223), .Y(n_255) );
BUFx12f_ASAP7_75t_L g256 ( .A(n_173), .Y(n_256) );
OR2x2_ASAP7_75t_L g257 ( .A(n_166), .B(n_131), .Y(n_257) );
NOR2xp33_ASAP7_75t_R g258 ( .A(n_167), .B(n_4), .Y(n_258) );
BUFx12f_ASAP7_75t_L g259 ( .A(n_173), .Y(n_259) );
OR2x2_ASAP7_75t_SL g260 ( .A(n_179), .B(n_5), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_180), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_180), .Y(n_262) );
OR2x6_ASAP7_75t_L g263 ( .A(n_223), .B(n_148), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_223), .Y(n_264) );
INVx4_ASAP7_75t_L g265 ( .A(n_176), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_205), .B(n_6), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_182), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_197), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_170), .Y(n_269) );
INVx3_ASAP7_75t_SL g270 ( .A(n_197), .Y(n_270) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_195), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_166), .B(n_7), .Y(n_272) );
AOI22xp33_ASAP7_75t_SL g273 ( .A1(n_181), .A2(n_156), .B1(n_9), .B2(n_11), .Y(n_273) );
BUFx2_ASAP7_75t_L g274 ( .A(n_197), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_188), .B(n_148), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_179), .Y(n_276) );
NOR3xp33_ASAP7_75t_SL g277 ( .A(n_206), .B(n_8), .C(n_11), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_180), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_170), .B(n_156), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_180), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g281 ( .A1(n_171), .A2(n_148), .B(n_146), .C(n_156), .Y(n_281) );
INVx5_ASAP7_75t_L g282 ( .A(n_197), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_171), .B(n_146), .Y(n_283) );
INVx3_ASAP7_75t_L g284 ( .A(n_197), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_181), .B(n_146), .Y(n_285) );
NOR2xp33_ASAP7_75t_SL g286 ( .A(n_197), .B(n_12), .Y(n_286) );
CKINVDCx8_ASAP7_75t_R g287 ( .A(n_197), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_174), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_205), .B(n_13), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_208), .B(n_14), .Y(n_290) );
NOR2x1p5_ASAP7_75t_L g291 ( .A(n_208), .B(n_214), .Y(n_291) );
INVx5_ASAP7_75t_L g292 ( .A(n_213), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_213), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_213), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_174), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_214), .Y(n_296) );
OR2x6_ASAP7_75t_L g297 ( .A(n_192), .B(n_14), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_L g298 ( .A1(n_220), .A2(n_16), .B(n_17), .C(n_18), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_196), .B(n_16), .Y(n_299) );
BUFx3_ASAP7_75t_L g300 ( .A(n_213), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_229), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g302 ( .A1(n_239), .A2(n_228), .B1(n_203), .B2(n_209), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_241), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_301), .B(n_229), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_232), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_241), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_270), .A2(n_263), .B1(n_264), .B2(n_255), .Y(n_307) );
NOR2xp67_ASAP7_75t_SL g308 ( .A(n_287), .B(n_209), .Y(n_308) );
INVx4_ASAP7_75t_L g309 ( .A(n_270), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_261), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_238), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_291), .B(n_209), .Y(n_312) );
CKINVDCx16_ASAP7_75t_R g313 ( .A(n_238), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_296), .B(n_210), .Y(n_314) );
OAI21x1_ASAP7_75t_L g315 ( .A1(n_254), .A2(n_203), .B(n_183), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_261), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_251), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_251), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_251), .Y(n_319) );
INVx8_ASAP7_75t_L g320 ( .A(n_263), .Y(n_320) );
NOR2xp33_ASAP7_75t_R g321 ( .A(n_276), .B(n_213), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_266), .B(n_210), .Y(n_322) );
OAI221xp5_ASAP7_75t_L g323 ( .A1(n_244), .A2(n_191), .B1(n_211), .B2(n_195), .C(n_210), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_257), .B(n_176), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_266), .A2(n_213), .B1(n_191), .B2(n_211), .Y(n_325) );
INVx1_ASAP7_75t_SL g326 ( .A(n_258), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_263), .Y(n_327) );
BUFx4f_ASAP7_75t_L g328 ( .A(n_263), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_248), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_247), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_267), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_279), .A2(n_212), .B(n_230), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_258), .Y(n_333) );
INVxp67_ASAP7_75t_L g334 ( .A(n_266), .Y(n_334) );
AOI21x1_ASAP7_75t_L g335 ( .A1(n_279), .A2(n_175), .B(n_169), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_265), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_262), .A2(n_212), .B(n_230), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_272), .Y(n_338) );
NOR2x1_ASAP7_75t_L g339 ( .A(n_297), .B(n_211), .Y(n_339) );
INVx2_ASAP7_75t_SL g340 ( .A(n_250), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_267), .B(n_213), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_267), .B(n_213), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_276), .B(n_186), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_233), .B(n_186), .Y(n_344) );
A2O1A1Ixp33_ASAP7_75t_L g345 ( .A1(n_269), .A2(n_212), .B(n_230), .C(n_195), .Y(n_345) );
OAI22xp33_ASAP7_75t_L g346 ( .A1(n_297), .A2(n_191), .B1(n_211), .B2(n_186), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_248), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_293), .B(n_191), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_293), .B(n_300), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_271), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_250), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_300), .B(n_186), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_252), .A2(n_176), .B1(n_183), .B2(n_200), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_262), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_278), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_304), .B(n_289), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_350), .Y(n_357) );
INVx4_ASAP7_75t_L g358 ( .A(n_320), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_304), .B(n_290), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_350), .Y(n_360) );
AND2x4_ASAP7_75t_L g361 ( .A(n_312), .B(n_265), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_303), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_303), .Y(n_363) );
CKINVDCx16_ASAP7_75t_R g364 ( .A(n_313), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_305), .B(n_256), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_312), .A2(n_297), .B1(n_256), .B2(n_259), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_343), .B(n_259), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_334), .B(n_260), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_312), .A2(n_237), .B1(n_295), .B2(n_288), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_306), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_314), .A2(n_237), .B1(n_249), .B2(n_240), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_328), .A2(n_247), .B1(n_253), .B2(n_294), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_306), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_330), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_350), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_314), .A2(n_249), .B1(n_299), .B2(n_273), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_322), .A2(n_245), .B1(n_242), .B2(n_234), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_351), .Y(n_378) );
INVx1_ASAP7_75t_SL g379 ( .A(n_351), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_330), .Y(n_380) );
AOI21x1_ASAP7_75t_L g381 ( .A1(n_335), .A2(n_285), .B(n_275), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_338), .B(n_235), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_350), .Y(n_383) );
INVx4_ASAP7_75t_SL g384 ( .A(n_327), .Y(n_384) );
OA21x2_ASAP7_75t_L g385 ( .A1(n_345), .A2(n_281), .B(n_298), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_328), .A2(n_286), .B1(n_236), .B2(n_243), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_310), .Y(n_387) );
OAI21x1_ASAP7_75t_L g388 ( .A1(n_335), .A2(n_253), .B(n_284), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_356), .B(n_322), .Y(n_389) );
OAI221xp5_ASAP7_75t_L g390 ( .A1(n_368), .A2(n_246), .B1(n_324), .B2(n_298), .C(n_326), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_368), .A2(n_333), .B1(n_320), .B2(n_339), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_362), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_382), .A2(n_320), .B1(n_311), .B2(n_321), .Y(n_393) );
OAI22xp33_ASAP7_75t_L g394 ( .A1(n_386), .A2(n_320), .B1(n_311), .B2(n_327), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_358), .Y(n_395) );
OAI222xp33_ASAP7_75t_L g396 ( .A1(n_386), .A2(n_346), .B1(n_323), .B2(n_302), .C1(n_307), .C2(n_340), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_367), .A2(n_331), .B1(n_317), .B2(n_336), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_359), .A2(n_325), .B1(n_340), .B2(n_271), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_376), .A2(n_319), .B1(n_317), .B2(n_318), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g400 ( .A1(n_366), .A2(n_277), .B1(n_342), .B2(n_341), .C(n_344), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_362), .A2(n_271), .B1(n_350), .B2(n_309), .Y(n_401) );
OAI22xp33_ASAP7_75t_L g402 ( .A1(n_358), .A2(n_309), .B1(n_319), .B2(n_336), .Y(n_402) );
AOI22xp33_ASAP7_75t_SL g403 ( .A1(n_358), .A2(n_379), .B1(n_378), .B2(n_364), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_363), .A2(n_271), .B1(n_309), .B2(n_294), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_387), .Y(n_405) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_358), .A2(n_364), .B1(n_370), .B2(n_373), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_387), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_363), .Y(n_408) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_371), .A2(n_353), .B1(n_283), .B2(n_281), .C(n_317), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_370), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_373), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_374), .B(n_310), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g413 ( .A1(n_365), .A2(n_283), .B1(n_319), .B2(n_318), .C(n_336), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_374), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_380), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_380), .A2(n_318), .B1(n_316), .B2(n_354), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_405), .B(n_385), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_414), .B(n_385), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_414), .Y(n_419) );
OAI211xp5_ASAP7_75t_L g420 ( .A1(n_390), .A2(n_369), .B(n_377), .C(n_385), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_414), .B(n_385), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_405), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_405), .B(n_384), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_390), .A2(n_361), .B1(n_372), .B2(n_348), .Y(n_424) );
INVx2_ASAP7_75t_SL g425 ( .A(n_395), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_406), .A2(n_361), .B1(n_355), .B2(n_354), .C(n_183), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_416), .A2(n_360), .B(n_357), .Y(n_427) );
INVx1_ASAP7_75t_SL g428 ( .A(n_403), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_415), .B(n_361), .Y(n_429) );
AO21x2_ASAP7_75t_L g430 ( .A1(n_416), .A2(n_388), .B(n_381), .Y(n_430) );
NAND3xp33_ASAP7_75t_L g431 ( .A(n_399), .B(n_357), .C(n_383), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_415), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_407), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_415), .Y(n_434) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_407), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_394), .A2(n_361), .B1(n_348), .B2(n_355), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_407), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_392), .Y(n_438) );
OA211x2_ASAP7_75t_L g439 ( .A1(n_391), .A2(n_384), .B(n_18), .C(n_20), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_389), .A2(n_384), .B1(n_308), .B2(n_348), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_411), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_412), .B(n_384), .Y(n_442) );
A2O1A1Ixp33_ASAP7_75t_L g443 ( .A1(n_395), .A2(n_308), .B(n_337), .C(n_352), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_412), .B(n_384), .Y(n_444) );
NAND3xp33_ASAP7_75t_L g445 ( .A(n_409), .B(n_383), .C(n_357), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_408), .Y(n_446) );
AO21x2_ASAP7_75t_L g447 ( .A1(n_398), .A2(n_388), .B(n_381), .Y(n_447) );
AOI211xp5_ASAP7_75t_SL g448 ( .A1(n_396), .A2(n_332), .B(n_375), .C(n_383), .Y(n_448) );
OAI33xp33_ASAP7_75t_L g449 ( .A1(n_408), .A2(n_190), .A3(n_193), .B1(n_199), .B2(n_200), .B3(n_201), .Y(n_449) );
OAI221xp5_ASAP7_75t_L g450 ( .A1(n_400), .A2(n_265), .B1(n_375), .B2(n_280), .C(n_278), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_395), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_438), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_418), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_422), .B(n_410), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_418), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_446), .Y(n_456) );
INVx3_ASAP7_75t_L g457 ( .A(n_435), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_421), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_428), .B(n_389), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_446), .Y(n_460) );
AOI221xp5_ASAP7_75t_L g461 ( .A1(n_441), .A2(n_397), .B1(n_409), .B2(n_413), .C(n_393), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_437), .B(n_395), .Y(n_462) );
AOI221xp5_ASAP7_75t_SL g463 ( .A1(n_424), .A2(n_398), .B1(n_402), .B2(n_404), .C(n_401), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_425), .B(n_401), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_419), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_437), .B(n_375), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_437), .B(n_360), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_419), .B(n_360), .Y(n_468) );
OAI31xp33_ASAP7_75t_L g469 ( .A1(n_420), .A2(n_404), .A3(n_352), .B(n_274), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_432), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_421), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g472 ( .A(n_442), .Y(n_472) );
AOI322xp5_ASAP7_75t_L g473 ( .A1(n_432), .A2(n_17), .A3(n_22), .B1(n_352), .B2(n_349), .C1(n_185), .C2(n_198), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_434), .B(n_360), .Y(n_474) );
BUFx2_ASAP7_75t_L g475 ( .A(n_433), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_436), .A2(n_360), .B1(n_347), .B2(n_329), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_434), .Y(n_477) );
INVx4_ASAP7_75t_L g478 ( .A(n_451), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_417), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_429), .B(n_360), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_429), .B(n_349), .Y(n_481) );
OAI31xp33_ASAP7_75t_L g482 ( .A1(n_442), .A2(n_349), .A3(n_347), .B(n_329), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_417), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_435), .Y(n_484) );
OAI221xp5_ASAP7_75t_SL g485 ( .A1(n_440), .A2(n_175), .B1(n_168), .B2(n_169), .C(n_184), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_435), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_435), .Y(n_487) );
OAI33xp33_ASAP7_75t_L g488 ( .A1(n_445), .A2(n_201), .A3(n_202), .B1(n_207), .B2(n_215), .B3(n_221), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_444), .B(n_315), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_423), .B(n_451), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_430), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_430), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_430), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_451), .B(n_23), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_472), .B(n_425), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_472), .B(n_452), .Y(n_496) );
NOR2x1_ASAP7_75t_L g497 ( .A(n_478), .B(n_431), .Y(n_497) );
NAND2xp33_ASAP7_75t_R g498 ( .A(n_475), .B(n_427), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_475), .B(n_448), .Y(n_499) );
INVxp67_ASAP7_75t_L g500 ( .A(n_459), .Y(n_500) );
NOR2xp33_ASAP7_75t_R g501 ( .A(n_478), .B(n_439), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_465), .Y(n_502) );
NOR3xp33_ASAP7_75t_SL g503 ( .A(n_461), .B(n_449), .C(n_450), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_470), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_470), .B(n_447), .Y(n_505) );
NAND2xp67_ASAP7_75t_L g506 ( .A(n_490), .B(n_439), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_477), .B(n_447), .Y(n_507) );
INVx2_ASAP7_75t_SL g508 ( .A(n_478), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_490), .B(n_454), .Y(n_509) );
NAND2xp33_ASAP7_75t_R g510 ( .A(n_457), .B(n_447), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_454), .B(n_426), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_477), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_456), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_479), .B(n_443), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_456), .Y(n_515) );
OR2x6_ASAP7_75t_L g516 ( .A(n_462), .B(n_194), .Y(n_516) );
AND2x2_ASAP7_75t_SL g517 ( .A(n_494), .B(n_268), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_481), .A2(n_280), .B1(n_284), .B2(n_268), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_462), .B(n_27), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_460), .B(n_41), .Y(n_520) );
INVxp67_ASAP7_75t_L g521 ( .A(n_494), .Y(n_521) );
NOR3xp33_ASAP7_75t_SL g522 ( .A(n_469), .B(n_488), .C(n_482), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g523 ( .A(n_480), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_483), .Y(n_524) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_491), .A2(n_169), .B(n_222), .Y(n_525) );
INVx1_ASAP7_75t_SL g526 ( .A(n_466), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_453), .B(n_50), .Y(n_527) );
INVxp67_ASAP7_75t_SL g528 ( .A(n_491), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_SL g529 ( .A1(n_492), .A2(n_185), .B(n_175), .C(n_168), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_455), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_455), .B(n_458), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_458), .B(n_52), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_500), .A2(n_469), .B1(n_489), .B2(n_464), .Y(n_533) );
OAI21xp33_ASAP7_75t_SL g534 ( .A1(n_508), .A2(n_473), .B(n_482), .Y(n_534) );
AOI211xp5_ASAP7_75t_L g535 ( .A1(n_499), .A2(n_463), .B(n_485), .C(n_476), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_496), .B(n_471), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_L g537 ( .A1(n_522), .A2(n_493), .B(n_492), .C(n_476), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_513), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_515), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_524), .B(n_493), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_523), .B(n_474), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_509), .B(n_466), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_526), .Y(n_543) );
INVxp67_ASAP7_75t_SL g544 ( .A(n_528), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_503), .A2(n_457), .B1(n_484), .B2(n_487), .Y(n_545) );
OAI21xp33_ASAP7_75t_L g546 ( .A1(n_506), .A2(n_487), .B(n_468), .Y(n_546) );
AOI211xp5_ASAP7_75t_L g547 ( .A1(n_501), .A2(n_486), .B(n_467), .C(n_198), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_502), .Y(n_548) );
OAI22xp33_ASAP7_75t_L g549 ( .A1(n_521), .A2(n_292), .B1(n_282), .B2(n_284), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_531), .B(n_54), .Y(n_550) );
O2A1O1Ixp33_ASAP7_75t_L g551 ( .A1(n_520), .A2(n_185), .B(n_221), .C(n_227), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_502), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_504), .Y(n_553) );
OAI32xp33_ASAP7_75t_L g554 ( .A1(n_498), .A2(n_495), .A3(n_510), .B1(n_514), .B2(n_532), .Y(n_554) );
OAI32xp33_ASAP7_75t_L g555 ( .A1(n_498), .A2(n_268), .A3(n_222), .B1(n_187), .B2(n_221), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_529), .A2(n_292), .B(n_282), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_504), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_517), .A2(n_292), .B1(n_282), .B2(n_183), .Y(n_558) );
AOI222xp33_ASAP7_75t_L g559 ( .A1(n_511), .A2(n_168), .B1(n_227), .B2(n_222), .C1(n_216), .C2(n_204), .Y(n_559) );
OAI222xp33_ASAP7_75t_L g560 ( .A1(n_516), .A2(n_55), .B1(n_60), .B2(n_62), .C1(n_64), .C2(n_65), .Y(n_560) );
OAI22xp33_ASAP7_75t_SL g561 ( .A1(n_516), .A2(n_66), .B1(n_67), .B2(n_68), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_531), .B(n_72), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_512), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_512), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_548), .Y(n_565) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_544), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_538), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_539), .Y(n_568) );
XOR2x2_ASAP7_75t_L g569 ( .A(n_547), .B(n_517), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_534), .B(n_497), .Y(n_570) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_543), .Y(n_571) );
INVx1_ASAP7_75t_SL g572 ( .A(n_541), .Y(n_572) );
NAND3xp33_ASAP7_75t_L g573 ( .A(n_535), .B(n_507), .C(n_505), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_542), .B(n_530), .Y(n_574) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_536), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_540), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_536), .B(n_519), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_552), .B(n_527), .Y(n_578) );
NAND2x1_ASAP7_75t_L g579 ( .A(n_553), .B(n_525), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_557), .B(n_525), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_563), .B(n_518), .Y(n_581) );
NOR3xp33_ASAP7_75t_SL g582 ( .A(n_554), .B(n_194), .C(n_219), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_533), .A2(n_204), .B1(n_216), .B2(n_194), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_564), .Y(n_584) );
NAND2x1_ASAP7_75t_L g585 ( .A(n_545), .B(n_194), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_565), .Y(n_586) );
AND4x1_ASAP7_75t_L g587 ( .A(n_582), .B(n_533), .C(n_537), .D(n_546), .Y(n_587) );
OAI21xp5_ASAP7_75t_L g588 ( .A1(n_570), .A2(n_560), .B(n_561), .Y(n_588) );
AOI222xp33_ASAP7_75t_L g589 ( .A1(n_570), .A2(n_560), .B1(n_562), .B2(n_550), .C1(n_555), .C2(n_558), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_565), .Y(n_590) );
INVxp67_ASAP7_75t_L g591 ( .A(n_571), .Y(n_591) );
OAI21xp33_ASAP7_75t_SL g592 ( .A1(n_566), .A2(n_559), .B(n_556), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_574), .B(n_549), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_573), .B(n_551), .Y(n_594) );
OAI22xp33_ASAP7_75t_SL g595 ( .A1(n_575), .A2(n_219), .B1(n_231), .B2(n_585), .Y(n_595) );
XNOR2x1_ASAP7_75t_L g596 ( .A(n_572), .B(n_219), .Y(n_596) );
AOI21xp33_ASAP7_75t_L g597 ( .A1(n_585), .A2(n_219), .B(n_231), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_576), .B(n_231), .Y(n_598) );
OAI22xp33_ASAP7_75t_SL g599 ( .A1(n_577), .A2(n_567), .B1(n_568), .B2(n_579), .Y(n_599) );
AOI21xp33_ASAP7_75t_L g600 ( .A1(n_592), .A2(n_583), .B(n_580), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_591), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_591), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_593), .Y(n_603) );
OAI21xp5_ASAP7_75t_L g604 ( .A1(n_588), .A2(n_569), .B(n_579), .Y(n_604) );
NOR2xp33_ASAP7_75t_R g605 ( .A(n_594), .B(n_569), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_589), .A2(n_581), .B1(n_578), .B2(n_584), .Y(n_606) );
INVx1_ASAP7_75t_SL g607 ( .A(n_596), .Y(n_607) );
AOI211xp5_ASAP7_75t_L g608 ( .A1(n_599), .A2(n_595), .B(n_597), .C(n_598), .Y(n_608) );
OAI22xp33_ASAP7_75t_L g609 ( .A1(n_586), .A2(n_590), .B1(n_587), .B2(n_598), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_L g610 ( .A1(n_590), .A2(n_570), .B(n_592), .C(n_588), .Y(n_610) );
NOR2x1_ASAP7_75t_L g611 ( .A(n_588), .B(n_570), .Y(n_611) );
NOR3xp33_ASAP7_75t_SL g612 ( .A(n_588), .B(n_592), .C(n_570), .Y(n_612) );
OR4x2_ASAP7_75t_L g613 ( .A(n_605), .B(n_611), .C(n_604), .D(n_612), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_606), .B(n_603), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_601), .Y(n_615) );
OAI211xp5_ASAP7_75t_SL g616 ( .A1(n_610), .A2(n_606), .B(n_609), .C(n_607), .Y(n_616) );
INVx1_ASAP7_75t_SL g617 ( .A(n_602), .Y(n_617) );
OAI211xp5_ASAP7_75t_L g618 ( .A1(n_616), .A2(n_605), .B(n_600), .C(n_608), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_617), .Y(n_619) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_619), .Y(n_620) );
XOR2x1_ASAP7_75t_L g621 ( .A(n_618), .B(n_613), .Y(n_621) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_620), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_621), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_622), .Y(n_624) );
OA22x2_ASAP7_75t_L g625 ( .A1(n_624), .A2(n_623), .B1(n_614), .B2(n_615), .Y(n_625) );
endmodule