module real_aes_9341_n_297 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_286, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_287, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_293, n_124, n_22, n_173, n_191, n_209, n_296, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_288, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_295, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_294, n_227, n_67, n_92, n_33, n_206, n_258, n_291, n_148, n_88, n_1758, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_292, n_116, n_94, n_229, n_289, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_290, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_297);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_286;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_287;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_293;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_296;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_288;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_295;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_294;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_291;
input n_148;
input n_88;
input n_1758;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_292;
input n_116;
input n_94;
input n_229;
input n_289;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_290;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_297;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1744;
wire n_1044;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1382;
wire n_875;
wire n_951;
wire n_1225;
wire n_1199;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_1745;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_1712;
wire n_667;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1741;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_602;
wire n_402;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_492;
wire n_407;
wire n_419;
wire n_1699;
wire n_730;
wire n_1023;
wire n_1748;
wire n_1403;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1172;
wire n_459;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_1185;
wire n_661;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1175;
wire n_1170;
wire n_778;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_317;
wire n_1595;
wire n_321;
wire n_1735;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1360;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_1430;
wire n_907;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_1352;
wire n_394;
wire n_1280;
wire n_1323;
wire n_729;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
INVxp33_ASAP7_75t_L g1014 ( .A(n_0), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_0), .A2(n_36), .B1(n_892), .B2(n_1042), .Y(n_1041) );
OAI222xp33_ASAP7_75t_L g1408 ( .A1(n_1), .A2(n_43), .B1(n_176), .B2(n_1409), .C1(n_1411), .C2(n_1412), .Y(n_1408) );
AOI221xp5_ASAP7_75t_L g1434 ( .A1(n_1), .A2(n_176), .B1(n_1435), .B2(n_1436), .C(n_1437), .Y(n_1434) );
INVx1_ASAP7_75t_L g1516 ( .A(n_2), .Y(n_1516) );
INVx1_ASAP7_75t_L g1167 ( .A(n_3), .Y(n_1167) );
AOI22xp33_ASAP7_75t_L g1703 ( .A1(n_4), .A2(n_15), .B1(n_475), .B2(n_1704), .Y(n_1703) );
OAI22xp5_ASAP7_75t_L g1732 ( .A1(n_4), .A2(n_15), .B1(n_566), .B2(n_1136), .Y(n_1732) );
OAI221xp5_ASAP7_75t_L g682 ( .A1(n_5), .A2(n_285), .B1(n_442), .B2(n_683), .C(n_684), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g739 ( .A1(n_5), .A2(n_290), .B1(n_740), .B2(n_741), .C(n_743), .Y(n_739) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_6), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_6), .B(n_226), .Y(n_331) );
AND2x2_ASAP7_75t_L g440 ( .A(n_6), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g490 ( .A(n_6), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g1309 ( .A1(n_7), .A2(n_14), .B1(n_810), .B2(n_1207), .Y(n_1309) );
INVx1_ASAP7_75t_L g1333 ( .A(n_7), .Y(n_1333) );
OA22x2_ASAP7_75t_L g1336 ( .A1(n_8), .A2(n_1337), .B1(n_1388), .B2(n_1389), .Y(n_1336) );
INVxp67_ASAP7_75t_SL g1389 ( .A(n_8), .Y(n_1389) );
INVxp67_ASAP7_75t_L g1021 ( .A(n_9), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_9), .A2(n_89), .B1(n_888), .B2(n_892), .Y(n_1047) );
INVxp33_ASAP7_75t_SL g420 ( .A(n_10), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_10), .A2(n_243), .B1(n_473), .B2(n_477), .Y(n_481) );
INVx1_ASAP7_75t_L g775 ( .A(n_11), .Y(n_775) );
AOI21xp5_ASAP7_75t_L g383 ( .A1(n_12), .A2(n_384), .B(n_388), .Y(n_383) );
INVx1_ASAP7_75t_L g457 ( .A(n_12), .Y(n_457) );
OAI332xp33_ASAP7_75t_L g1348 ( .A1(n_13), .A2(n_486), .A3(n_520), .B1(n_1349), .B2(n_1352), .B3(n_1355), .C1(n_1358), .C2(n_1361), .Y(n_1348) );
INVx1_ASAP7_75t_L g1386 ( .A(n_13), .Y(n_1386) );
AOI221xp5_ASAP7_75t_L g1328 ( .A1(n_14), .A2(n_129), .B1(n_1329), .B2(n_1331), .C(n_1332), .Y(n_1328) );
INVx1_ASAP7_75t_L g1575 ( .A(n_16), .Y(n_1575) );
INVx1_ASAP7_75t_L g968 ( .A(n_17), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_18), .A2(n_121), .B1(n_901), .B2(n_902), .Y(n_900) );
INVxp67_ASAP7_75t_SL g934 ( .A(n_18), .Y(n_934) );
INVxp33_ASAP7_75t_L g1253 ( .A(n_19), .Y(n_1253) );
AOI221xp5_ASAP7_75t_L g1280 ( .A1(n_19), .A2(n_162), .B1(n_401), .B2(n_576), .C(n_984), .Y(n_1280) );
INVx1_ASAP7_75t_L g906 ( .A(n_20), .Y(n_906) );
INVx1_ASAP7_75t_L g770 ( .A(n_21), .Y(n_770) );
INVx1_ASAP7_75t_L g1470 ( .A(n_22), .Y(n_1470) );
INVx1_ASAP7_75t_L g580 ( .A(n_23), .Y(n_580) );
AO221x2_ASAP7_75t_L g1480 ( .A1(n_24), .A2(n_63), .B1(n_1452), .B2(n_1460), .C(n_1481), .Y(n_1480) );
INVx2_ASAP7_75t_L g340 ( .A(n_25), .Y(n_340) );
OR2x2_ASAP7_75t_L g357 ( .A(n_25), .B(n_338), .Y(n_357) );
INVx1_ASAP7_75t_L g1283 ( .A(n_26), .Y(n_1283) );
INVx1_ASAP7_75t_L g1482 ( .A(n_27), .Y(n_1482) );
AOI221xp5_ASAP7_75t_L g1205 ( .A1(n_28), .A2(n_53), .B1(n_1206), .B2(n_1207), .C(n_1208), .Y(n_1205) );
INVx1_ASAP7_75t_L g1238 ( .A(n_28), .Y(n_1238) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_29), .Y(n_614) );
INVx1_ASAP7_75t_L g904 ( .A(n_30), .Y(n_904) );
AOI22xp33_ASAP7_75t_SL g890 ( .A1(n_31), .A2(n_159), .B1(n_891), .B2(n_892), .Y(n_890) );
INVxp33_ASAP7_75t_SL g917 ( .A(n_31), .Y(n_917) );
OR2x2_ASAP7_75t_L g330 ( .A(n_32), .B(n_331), .Y(n_330) );
BUFx2_ASAP7_75t_L g334 ( .A(n_32), .Y(n_334) );
BUFx2_ASAP7_75t_L g429 ( .A(n_32), .Y(n_429) );
INVx1_ASAP7_75t_L g439 ( .A(n_32), .Y(n_439) );
OAI221xp5_ASAP7_75t_L g1148 ( .A1(n_33), .A2(n_193), .B1(n_697), .B2(n_919), .C(n_921), .Y(n_1148) );
OAI22xp33_ASAP7_75t_SL g1178 ( .A1(n_33), .A2(n_193), .B1(n_1179), .B2(n_1180), .Y(n_1178) );
CKINVDCx5p33_ASAP7_75t_R g1351 ( .A(n_34), .Y(n_1351) );
INVx1_ASAP7_75t_L g1573 ( .A(n_35), .Y(n_1573) );
INVxp33_ASAP7_75t_L g1010 ( .A(n_36), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_37), .A2(n_179), .B1(n_658), .B2(n_1111), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g1131 ( .A1(n_37), .A2(n_179), .B1(n_611), .B2(n_804), .Y(n_1131) );
AOI221xp5_ASAP7_75t_L g1112 ( .A1(n_38), .A2(n_133), .B1(n_435), .B2(n_521), .C(n_1113), .Y(n_1112) );
INVx1_ASAP7_75t_L g1127 ( .A(n_38), .Y(n_1127) );
CKINVDCx5p33_ASAP7_75t_R g1356 ( .A(n_39), .Y(n_1356) );
INVxp67_ASAP7_75t_L g709 ( .A(n_40), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g748 ( .A1(n_40), .A2(n_197), .B1(n_749), .B2(n_750), .C(n_754), .Y(n_748) );
INVxp33_ASAP7_75t_L g1146 ( .A(n_41), .Y(n_1146) );
AOI221xp5_ASAP7_75t_L g1172 ( .A1(n_41), .A2(n_46), .B1(n_409), .B2(n_984), .C(n_1173), .Y(n_1172) );
AOI221xp5_ASAP7_75t_L g1308 ( .A1(n_42), .A2(n_129), .B1(n_374), .B2(n_740), .C(n_899), .Y(n_1308) );
INVx1_ASAP7_75t_L g1334 ( .A(n_42), .Y(n_1334) );
INVx1_ASAP7_75t_L g1438 ( .A(n_43), .Y(n_1438) );
INVxp67_ASAP7_75t_L g704 ( .A(n_44), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_44), .A2(n_199), .B1(n_408), .B2(n_756), .Y(n_755) );
CKINVDCx16_ASAP7_75t_R g1290 ( .A(n_45), .Y(n_1290) );
INVxp33_ASAP7_75t_L g1144 ( .A(n_46), .Y(n_1144) );
AOI22xp33_ASAP7_75t_SL g1705 ( .A1(n_47), .A2(n_88), .B1(n_1105), .B2(n_1113), .Y(n_1705) );
INVx1_ASAP7_75t_L g1731 ( .A(n_47), .Y(n_1731) );
INVx1_ASAP7_75t_L g1569 ( .A(n_48), .Y(n_1569) );
INVx1_ASAP7_75t_L g1265 ( .A(n_49), .Y(n_1265) );
INVxp33_ASAP7_75t_SL g1147 ( .A(n_50), .Y(n_1147) );
AOI22xp33_ASAP7_75t_L g1175 ( .A1(n_50), .A2(n_280), .B1(n_1176), .B2(n_1177), .Y(n_1175) );
INVx1_ASAP7_75t_L g1165 ( .A(n_51), .Y(n_1165) );
AOI22xp33_ASAP7_75t_SL g1701 ( .A1(n_52), .A2(n_236), .B1(n_1105), .B2(n_1113), .Y(n_1701) );
AOI22xp33_ASAP7_75t_L g1722 ( .A1(n_52), .A2(n_217), .B1(n_981), .B2(n_1189), .Y(n_1722) );
INVx1_ASAP7_75t_L g1241 ( .A(n_53), .Y(n_1241) );
INVx1_ASAP7_75t_L g1222 ( .A(n_54), .Y(n_1222) );
INVx1_ASAP7_75t_L g686 ( .A(n_55), .Y(n_686) );
INVx1_ASAP7_75t_L g907 ( .A(n_56), .Y(n_907) );
AOI221xp5_ASAP7_75t_SL g1303 ( .A1(n_57), .A2(n_77), .B1(n_409), .B2(n_889), .C(n_1304), .Y(n_1303) );
INVx1_ASAP7_75t_L g1319 ( .A(n_57), .Y(n_1319) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_58), .A2(n_218), .B1(n_584), .B2(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g659 ( .A(n_58), .Y(n_659) );
AOI22xp33_ASAP7_75t_SL g803 ( .A1(n_59), .A2(n_265), .B1(n_804), .B2(n_806), .Y(n_803) );
INVxp67_ASAP7_75t_SL g866 ( .A(n_59), .Y(n_866) );
INVx1_ASAP7_75t_L g1300 ( .A(n_60), .Y(n_1300) );
INVx1_ASAP7_75t_L g1121 ( .A(n_61), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_61), .A2(n_167), .B1(n_804), .B2(n_1135), .Y(n_1134) );
OAI221xp5_ASAP7_75t_L g953 ( .A1(n_62), .A2(n_143), .B1(n_690), .B2(n_696), .C(n_700), .Y(n_953) );
OAI33xp33_ASAP7_75t_L g986 ( .A1(n_62), .A2(n_143), .A3(n_415), .B1(n_735), .B2(n_987), .B3(n_1758), .Y(n_986) );
XNOR2x2_ASAP7_75t_L g1694 ( .A(n_63), .B(n_1695), .Y(n_1694) );
AOI22xp33_ASAP7_75t_L g1740 ( .A1(n_63), .A2(n_1741), .B1(n_1744), .B2(n_1749), .Y(n_1740) );
INVx1_ASAP7_75t_L g1299 ( .A(n_64), .Y(n_1299) );
CKINVDCx5p33_ASAP7_75t_R g1357 ( .A(n_65), .Y(n_1357) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_66), .Y(n_824) );
AOI22xp33_ASAP7_75t_SL g811 ( .A1(n_67), .A2(n_137), .B1(n_806), .B2(n_812), .Y(n_811) );
OAI221xp5_ASAP7_75t_L g853 ( .A1(n_67), .A2(n_854), .B1(n_856), .B2(n_863), .C(n_873), .Y(n_853) );
OAI222xp33_ASAP7_75t_L g1413 ( .A1(n_68), .A2(n_154), .B1(n_234), .B2(n_1180), .C1(n_1311), .C2(n_1414), .Y(n_1413) );
INVx1_ASAP7_75t_L g1419 ( .A(n_68), .Y(n_1419) );
INVx1_ASAP7_75t_L g1493 ( .A(n_69), .Y(n_1493) );
CKINVDCx16_ASAP7_75t_R g1498 ( .A(n_70), .Y(n_1498) );
AOI22xp33_ASAP7_75t_SL g1702 ( .A1(n_71), .A2(n_217), .B1(n_1101), .B2(n_1111), .Y(n_1702) );
AOI21xp33_ASAP7_75t_L g1723 ( .A1(n_71), .A2(n_563), .B(n_805), .Y(n_1723) );
OAI22xp5_ASAP7_75t_L g1339 ( .A1(n_72), .A2(n_223), .B1(n_1340), .B2(n_1342), .Y(n_1339) );
CKINVDCx5p33_ASAP7_75t_R g1385 ( .A(n_72), .Y(n_1385) );
INVxp33_ASAP7_75t_SL g509 ( .A(n_73), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g564 ( .A1(n_73), .A2(n_281), .B1(n_552), .B2(n_565), .C(n_568), .Y(n_564) );
INVx1_ASAP7_75t_L g716 ( .A(n_74), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g1399 ( .A1(n_75), .A2(n_104), .B1(n_815), .B2(n_1218), .Y(n_1399) );
INVx1_ASAP7_75t_L g1424 ( .A(n_75), .Y(n_1424) );
AOI22xp33_ASAP7_75t_L g1402 ( .A1(n_76), .A2(n_157), .B1(n_892), .B2(n_1403), .Y(n_1402) );
INVx1_ASAP7_75t_L g1431 ( .A(n_76), .Y(n_1431) );
INVx1_ASAP7_75t_L g1318 ( .A(n_77), .Y(n_1318) );
INVxp67_ASAP7_75t_L g1019 ( .A(n_78), .Y(n_1019) );
AOI221xp5_ASAP7_75t_L g1046 ( .A1(n_78), .A2(n_200), .B1(n_374), .B2(n_401), .C(n_899), .Y(n_1046) );
INVxp33_ASAP7_75t_L g780 ( .A(n_79), .Y(n_780) );
AOI221xp5_ASAP7_75t_L g842 ( .A1(n_79), .A2(n_264), .B1(n_843), .B2(n_845), .C(n_846), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_80), .A2(n_198), .B1(n_815), .B2(n_816), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g874 ( .A1(n_80), .A2(n_198), .B1(n_875), .B2(n_877), .Y(n_874) );
INVx1_ASAP7_75t_L g1517 ( .A(n_81), .Y(n_1517) );
CKINVDCx5p33_ASAP7_75t_R g1118 ( .A(n_82), .Y(n_1118) );
INVxp67_ASAP7_75t_SL g962 ( .A(n_83), .Y(n_962) );
AOI221xp5_ASAP7_75t_L g991 ( .A1(n_83), .A2(n_147), .B1(n_992), .B2(n_993), .C(n_994), .Y(n_991) );
OAI221xp5_ASAP7_75t_L g1294 ( .A1(n_84), .A2(n_244), .B1(n_1295), .B2(n_1296), .C(n_1297), .Y(n_1294) );
INVx1_ASAP7_75t_L g1326 ( .A(n_84), .Y(n_1326) );
INVxp67_ASAP7_75t_SL g398 ( .A(n_85), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_85), .A2(n_208), .B1(n_471), .B2(n_479), .Y(n_482) );
INVx1_ASAP7_75t_L g722 ( .A(n_86), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g1343 ( .A1(n_87), .A2(n_163), .B1(n_329), .B2(n_1344), .Y(n_1343) );
CKINVDCx5p33_ASAP7_75t_R g1383 ( .A(n_87), .Y(n_1383) );
NOR2xp33_ASAP7_75t_L g1717 ( .A(n_88), .B(n_419), .Y(n_1717) );
INVxp67_ASAP7_75t_L g1023 ( .A(n_89), .Y(n_1023) );
OAI221xp5_ASAP7_75t_L g689 ( .A1(n_90), .A2(n_189), .B1(n_690), .B2(n_695), .C(n_700), .Y(n_689) );
OAI221xp5_ASAP7_75t_SL g732 ( .A1(n_90), .A2(n_189), .B1(n_733), .B2(n_734), .C(n_736), .Y(n_732) );
INVx1_ASAP7_75t_L g1714 ( .A(n_91), .Y(n_1714) );
AOI22xp33_ASAP7_75t_L g1726 ( .A1(n_91), .A2(n_145), .B1(n_805), .B2(n_981), .Y(n_1726) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_92), .A2(n_118), .B1(n_369), .B2(n_374), .C(n_375), .Y(n_368) );
INVxp33_ASAP7_75t_L g450 ( .A(n_92), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_93), .A2(n_263), .B1(n_553), .B2(n_601), .C(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g642 ( .A(n_93), .Y(n_642) );
XNOR2xp5_ASAP7_75t_L g1058 ( .A(n_94), .B(n_1059), .Y(n_1058) );
INVxp33_ASAP7_75t_L g1154 ( .A(n_95), .Y(n_1154) );
AOI22xp33_ASAP7_75t_L g1186 ( .A1(n_95), .A2(n_250), .B1(n_369), .B2(n_1187), .Y(n_1186) );
AOI22xp5_ASAP7_75t_L g1473 ( .A1(n_96), .A2(n_158), .B1(n_1474), .B2(n_1477), .Y(n_1473) );
CKINVDCx16_ASAP7_75t_R g1501 ( .A(n_97), .Y(n_1501) );
INVx1_ASAP7_75t_L g338 ( .A(n_98), .Y(n_338) );
INVx1_ASAP7_75t_L g391 ( .A(n_98), .Y(n_391) );
INVx1_ASAP7_75t_L g941 ( .A(n_99), .Y(n_941) );
CKINVDCx5p33_ASAP7_75t_R g1077 ( .A(n_100), .Y(n_1077) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_101), .A2(n_251), .B1(n_359), .B2(n_364), .Y(n_358) );
INVxp67_ASAP7_75t_SL g501 ( .A(n_101), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_102), .A2(n_229), .B1(n_369), .B2(n_408), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_102), .A2(n_229), .B1(n_471), .B2(n_473), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g1202 ( .A1(n_103), .A2(n_293), .B1(n_895), .B2(n_1203), .Y(n_1202) );
INVx1_ASAP7_75t_L g1226 ( .A(n_103), .Y(n_1226) );
INVx1_ASAP7_75t_L g1421 ( .A(n_104), .Y(n_1421) );
INVx1_ASAP7_75t_L g956 ( .A(n_105), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_105), .A2(n_187), .B1(n_997), .B2(n_998), .Y(n_996) );
OAI221xp5_ASAP7_75t_L g1015 ( .A1(n_106), .A2(n_132), .B1(n_919), .B2(n_920), .C(n_1016), .Y(n_1015) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_106), .A2(n_132), .B1(n_895), .B2(n_1044), .Y(n_1043) );
INVxp67_ASAP7_75t_SL g1259 ( .A(n_107), .Y(n_1259) );
AOI221xp5_ASAP7_75t_L g1277 ( .A1(n_107), .A2(n_230), .B1(n_630), .B2(n_740), .C(n_899), .Y(n_1277) );
INVx1_ASAP7_75t_L g1298 ( .A(n_108), .Y(n_1298) );
AOI221xp5_ASAP7_75t_L g1320 ( .A1(n_108), .A2(n_244), .B1(n_1321), .B2(n_1323), .C(n_1325), .Y(n_1320) );
INVx1_ASAP7_75t_L g1708 ( .A(n_109), .Y(n_1708) );
AOI21xp5_ASAP7_75t_L g1727 ( .A1(n_109), .A2(n_555), .B(n_617), .Y(n_1727) );
INVxp33_ASAP7_75t_SL g1250 ( .A(n_110), .Y(n_1250) );
AOI22xp33_ASAP7_75t_L g1281 ( .A1(n_110), .A2(n_128), .B1(n_374), .B2(n_586), .Y(n_1281) );
INVxp33_ASAP7_75t_L g948 ( .A(n_111), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_111), .A2(n_273), .B1(n_980), .B2(n_981), .Y(n_979) );
CKINVDCx5p33_ASAP7_75t_R g728 ( .A(n_112), .Y(n_728) );
INVx1_ASAP7_75t_L g1081 ( .A(n_113), .Y(n_1081) );
OAI221xp5_ASAP7_75t_L g1106 ( .A1(n_113), .A2(n_190), .B1(n_852), .B2(n_1107), .C(n_1109), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_114), .A2(n_242), .B1(n_756), .B2(n_809), .Y(n_808) );
INVxp67_ASAP7_75t_SL g860 ( .A(n_114), .Y(n_860) );
INVx1_ASAP7_75t_L g965 ( .A(n_115), .Y(n_965) );
INVx1_ASAP7_75t_L g1467 ( .A(n_116), .Y(n_1467) );
INVx1_ASAP7_75t_L g1072 ( .A(n_117), .Y(n_1072) );
AOI221xp5_ASAP7_75t_L g1100 ( .A1(n_117), .A2(n_174), .B1(n_444), .B2(n_1101), .C(n_1102), .Y(n_1100) );
OAI221xp5_ASAP7_75t_L g431 ( .A1(n_118), .A2(n_155), .B1(n_432), .B2(n_442), .C(n_449), .Y(n_431) );
INVx1_ASAP7_75t_L g1312 ( .A(n_119), .Y(n_1312) );
AO221x2_ASAP7_75t_L g1514 ( .A1(n_120), .A2(n_206), .B1(n_1460), .B2(n_1500), .C(n_1515), .Y(n_1514) );
INVxp33_ASAP7_75t_L g924 ( .A(n_121), .Y(n_924) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_122), .Y(n_604) );
INVx1_ASAP7_75t_L g893 ( .A(n_123), .Y(n_893) );
OAI22xp33_ASAP7_75t_SL g628 ( .A1(n_124), .A2(n_231), .B1(n_557), .B2(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g666 ( .A(n_124), .Y(n_666) );
INVx1_ASAP7_75t_L g1162 ( .A(n_125), .Y(n_1162) );
INVx1_ASAP7_75t_L g1262 ( .A(n_126), .Y(n_1262) );
AOI22xp33_ASAP7_75t_L g1278 ( .A1(n_126), .A2(n_188), .B1(n_892), .B2(n_1187), .Y(n_1278) );
INVx1_ASAP7_75t_L g303 ( .A(n_127), .Y(n_303) );
INVxp33_ASAP7_75t_SL g1254 ( .A(n_128), .Y(n_1254) );
INVx1_ASAP7_75t_L g532 ( .A(n_130), .Y(n_532) );
AOI221xp5_ASAP7_75t_L g551 ( .A1(n_130), .A2(n_228), .B1(n_552), .B2(n_553), .C(n_556), .Y(n_551) );
XNOR2x1_ASAP7_75t_L g1005 ( .A(n_131), .B(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g1130 ( .A(n_133), .Y(n_1130) );
AOI221xp5_ASAP7_75t_L g608 ( .A1(n_134), .A2(n_172), .B1(n_609), .B2(n_611), .C(n_613), .Y(n_608) );
INVx1_ASAP7_75t_L g671 ( .A(n_134), .Y(n_671) );
INVx1_ASAP7_75t_L g1027 ( .A(n_135), .Y(n_1027) );
INVx1_ASAP7_75t_L g1215 ( .A(n_136), .Y(n_1215) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_136), .A2(n_181), .B1(n_471), .B2(n_843), .Y(n_1236) );
OAI211xp5_ASAP7_75t_SL g834 ( .A1(n_137), .A2(n_835), .B(n_839), .C(n_848), .Y(n_834) );
INVx1_ASAP7_75t_L g970 ( .A(n_138), .Y(n_970) );
CKINVDCx5p33_ASAP7_75t_R g1117 ( .A(n_139), .Y(n_1117) );
CKINVDCx5p33_ASAP7_75t_R g615 ( .A(n_140), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g1479 ( .A1(n_141), .A2(n_196), .B1(n_1452), .B2(n_1460), .Y(n_1479) );
INVx1_ASAP7_75t_L g581 ( .A(n_142), .Y(n_581) );
AOI221xp5_ASAP7_75t_L g1400 ( .A1(n_144), .A2(n_204), .B1(n_401), .B2(n_563), .C(n_1401), .Y(n_1400) );
AOI221xp5_ASAP7_75t_L g1428 ( .A1(n_144), .A2(n_157), .B1(n_1321), .B2(n_1429), .C(n_1430), .Y(n_1428) );
INVx1_ASAP7_75t_L g1711 ( .A(n_145), .Y(n_1711) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_146), .A2(n_268), .B1(n_741), .B2(n_1218), .Y(n_1217) );
AOI22xp33_ASAP7_75t_L g1232 ( .A1(n_146), .A2(n_160), .B1(n_478), .B2(n_937), .Y(n_1232) );
INVxp33_ASAP7_75t_L g957 ( .A(n_147), .Y(n_957) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_148), .A2(n_177), .B1(n_374), .B2(n_400), .C(n_404), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_148), .A2(n_177), .B1(n_477), .B2(n_479), .Y(n_476) );
INVx1_ASAP7_75t_L g1243 ( .A(n_149), .Y(n_1243) );
OAI221xp5_ASAP7_75t_L g1347 ( .A1(n_150), .A2(n_248), .B1(n_690), .B2(n_696), .C(n_921), .Y(n_1347) );
OAI222xp33_ASAP7_75t_L g1373 ( .A1(n_150), .A2(n_163), .B1(n_248), .B2(n_733), .C1(n_734), .C2(n_1311), .Y(n_1373) );
OAI22xp5_ASAP7_75t_L g894 ( .A1(n_151), .A2(n_207), .B1(n_364), .B2(n_895), .Y(n_894) );
OAI221xp5_ASAP7_75t_L g918 ( .A1(n_151), .A2(n_207), .B1(n_919), .B2(n_920), .C(n_921), .Y(n_918) );
INVx1_ASAP7_75t_L g1483 ( .A(n_152), .Y(n_1483) );
AOI221xp5_ASAP7_75t_L g1398 ( .A1(n_153), .A2(n_169), .B1(n_409), .B2(n_889), .C(n_1304), .Y(n_1398) );
INVx1_ASAP7_75t_L g1422 ( .A(n_153), .Y(n_1422) );
INVx1_ASAP7_75t_L g1425 ( .A(n_154), .Y(n_1425) );
INVx1_ASAP7_75t_L g382 ( .A(n_155), .Y(n_382) );
INVx1_ASAP7_75t_L g790 ( .A(n_156), .Y(n_790) );
INVxp33_ASAP7_75t_L g912 ( .A(n_159), .Y(n_912) );
AOI221xp5_ASAP7_75t_L g1216 ( .A1(n_160), .A2(n_166), .B1(n_563), .B2(n_623), .C(n_1176), .Y(n_1216) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_161), .A2(n_238), .B1(n_435), .B2(n_548), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_161), .A2(n_258), .B1(n_584), .B2(n_585), .Y(n_583) );
INVxp33_ASAP7_75t_L g1251 ( .A(n_162), .Y(n_1251) );
INVx1_ASAP7_75t_L g1035 ( .A(n_164), .Y(n_1035) );
CKINVDCx5p33_ASAP7_75t_R g1698 ( .A(n_165), .Y(n_1698) );
AOI22xp33_ASAP7_75t_SL g1229 ( .A1(n_166), .A2(n_268), .B1(n_1230), .B2(n_1231), .Y(n_1229) );
INVx1_ASAP7_75t_L g1120 ( .A(n_167), .Y(n_1120) );
INVx1_ASAP7_75t_L g1221 ( .A(n_168), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g1233 ( .A1(n_168), .A2(n_202), .B1(n_478), .B2(n_1234), .Y(n_1233) );
INVx1_ASAP7_75t_L g1427 ( .A(n_169), .Y(n_1427) );
CKINVDCx5p33_ASAP7_75t_R g1407 ( .A(n_170), .Y(n_1407) );
AOI22xp5_ASAP7_75t_L g1508 ( .A1(n_171), .A2(n_191), .B1(n_1474), .B2(n_1477), .Y(n_1508) );
INVx1_ASAP7_75t_L g673 ( .A(n_172), .Y(n_673) );
INVx1_ASAP7_75t_L g908 ( .A(n_173), .Y(n_908) );
INVx1_ASAP7_75t_L g1092 ( .A(n_174), .Y(n_1092) );
OAI221xp5_ASAP7_75t_L g1255 ( .A1(n_175), .A2(n_294), .B1(n_697), .B2(n_919), .C(n_1016), .Y(n_1255) );
OAI22xp33_ASAP7_75t_L g1282 ( .A1(n_175), .A2(n_294), .B1(n_1179), .B2(n_1180), .Y(n_1282) );
INVx1_ASAP7_75t_L g518 ( .A(n_178), .Y(n_518) );
CKINVDCx16_ASAP7_75t_R g324 ( .A(n_180), .Y(n_324) );
INVx1_ASAP7_75t_L g1220 ( .A(n_181), .Y(n_1220) );
CKINVDCx5p33_ASAP7_75t_R g1699 ( .A(n_182), .Y(n_1699) );
XNOR2xp5_ASAP7_75t_L g1137 ( .A(n_183), .B(n_1138), .Y(n_1137) );
AOI22xp5_ASAP7_75t_L g1509 ( .A1(n_183), .A2(n_235), .B1(n_1500), .B2(n_1510), .Y(n_1509) );
CKINVDCx5p33_ASAP7_75t_R g622 ( .A(n_184), .Y(n_622) );
INVx1_ASAP7_75t_L g1245 ( .A(n_185), .Y(n_1245) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_186), .Y(n_305) );
AND3x2_ASAP7_75t_L g1453 ( .A(n_186), .B(n_303), .C(n_1454), .Y(n_1453) );
NAND2xp5_ASAP7_75t_L g1464 ( .A(n_186), .B(n_303), .Y(n_1464) );
INVx1_ASAP7_75t_L g961 ( .A(n_187), .Y(n_961) );
INVxp67_ASAP7_75t_SL g1258 ( .A(n_188), .Y(n_1258) );
INVx1_ASAP7_75t_L g1086 ( .A(n_190), .Y(n_1086) );
INVx1_ASAP7_75t_L g966 ( .A(n_192), .Y(n_966) );
INVx2_ASAP7_75t_L g316 ( .A(n_194), .Y(n_316) );
INVx1_ASAP7_75t_L g1301 ( .A(n_195), .Y(n_1301) );
XNOR2x2_ASAP7_75t_L g505 ( .A(n_196), .B(n_506), .Y(n_505) );
INVxp67_ASAP7_75t_SL g713 ( .A(n_197), .Y(n_713) );
INVxp33_ASAP7_75t_SL g706 ( .A(n_199), .Y(n_706) );
INVxp33_ASAP7_75t_L g1025 ( .A(n_200), .Y(n_1025) );
INVxp67_ASAP7_75t_L g1157 ( .A(n_201), .Y(n_1157) );
AOI221xp5_ASAP7_75t_L g1184 ( .A1(n_201), .A2(n_270), .B1(n_740), .B2(n_899), .C(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1201 ( .A(n_202), .Y(n_1201) );
CKINVDCx5p33_ASAP7_75t_R g1359 ( .A(n_203), .Y(n_1359) );
INVx1_ASAP7_75t_L g1433 ( .A(n_204), .Y(n_1433) );
AOI22xp5_ASAP7_75t_L g1504 ( .A1(n_205), .A2(n_213), .B1(n_1452), .B2(n_1460), .Y(n_1504) );
INVx1_ASAP7_75t_L g679 ( .A(n_206), .Y(n_679) );
INVxp33_ASAP7_75t_SL g417 ( .A(n_208), .Y(n_417) );
INVx1_ASAP7_75t_L g1030 ( .A(n_209), .Y(n_1030) );
AOI221xp5_ASAP7_75t_L g897 ( .A1(n_210), .A2(n_284), .B1(n_353), .B2(n_898), .C(n_899), .Y(n_897) );
INVxp67_ASAP7_75t_SL g930 ( .A(n_210), .Y(n_930) );
INVx1_ASAP7_75t_L g1454 ( .A(n_211), .Y(n_1454) );
INVx1_ASAP7_75t_L g528 ( .A(n_212), .Y(n_528) );
CKINVDCx16_ASAP7_75t_R g1458 ( .A(n_214), .Y(n_1458) );
INVx1_ASAP7_75t_L g511 ( .A(n_215), .Y(n_511) );
INVx1_ASAP7_75t_L g1571 ( .A(n_216), .Y(n_1571) );
INVx1_ASAP7_75t_L g661 ( .A(n_218), .Y(n_661) );
CKINVDCx5p33_ASAP7_75t_R g1350 ( .A(n_219), .Y(n_1350) );
INVx1_ASAP7_75t_L g1715 ( .A(n_220), .Y(n_1715) );
OAI211xp5_ASAP7_75t_L g1729 ( .A1(n_220), .A2(n_1311), .B(n_1730), .C(n_1733), .Y(n_1729) );
INVx1_ASAP7_75t_L g1268 ( .A(n_221), .Y(n_1268) );
CKINVDCx5p33_ASAP7_75t_R g974 ( .A(n_222), .Y(n_974) );
CKINVDCx5p33_ASAP7_75t_R g1381 ( .A(n_223), .Y(n_1381) );
CKINVDCx5p33_ASAP7_75t_R g1360 ( .A(n_224), .Y(n_1360) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_225), .Y(n_637) );
INVx1_ASAP7_75t_L g318 ( .A(n_226), .Y(n_318) );
INVx2_ASAP7_75t_L g441 ( .A(n_226), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g635 ( .A(n_227), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_228), .A2(n_232), .B1(n_534), .B2(n_537), .Y(n_533) );
INVxp67_ASAP7_75t_SL g1261 ( .A(n_230), .Y(n_1261) );
INVx1_ASAP7_75t_L g656 ( .A(n_231), .Y(n_656) );
INVx1_ASAP7_75t_L g559 ( .A(n_232), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g1503 ( .A1(n_233), .A2(n_257), .B1(n_1474), .B2(n_1477), .Y(n_1503) );
INVx1_ASAP7_75t_L g1418 ( .A(n_234), .Y(n_1418) );
INVx1_ASAP7_75t_L g1720 ( .A(n_236), .Y(n_1720) );
INVxp33_ASAP7_75t_L g1013 ( .A(n_237), .Y(n_1013) );
AOI221xp5_ASAP7_75t_L g1040 ( .A1(n_237), .A2(n_240), .B1(n_409), .B2(n_887), .C(n_889), .Y(n_1040) );
OAI22xp33_ASAP7_75t_L g587 ( .A1(n_238), .A2(n_272), .B1(n_588), .B2(n_589), .Y(n_587) );
INVx1_ASAP7_75t_L g949 ( .A(n_239), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g985 ( .A(n_239), .B(n_384), .Y(n_985) );
INVxp33_ASAP7_75t_L g1011 ( .A(n_240), .Y(n_1011) );
INVx1_ASAP7_75t_L g719 ( .A(n_241), .Y(n_719) );
INVxp67_ASAP7_75t_SL g872 ( .A(n_242), .Y(n_872) );
INVxp67_ASAP7_75t_SL g349 ( .A(n_243), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g1306 ( .A1(n_245), .A2(n_260), .B1(n_891), .B2(n_902), .Y(n_1306) );
OAI221xp5_ASAP7_75t_L g1316 ( .A1(n_245), .A2(n_260), .B1(n_707), .B2(n_840), .C(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g796 ( .A(n_246), .Y(n_796) );
INVx1_ASAP7_75t_L g1266 ( .A(n_247), .Y(n_1266) );
INVx1_ASAP7_75t_L g943 ( .A(n_249), .Y(n_943) );
INVxp67_ASAP7_75t_L g1160 ( .A(n_250), .Y(n_1160) );
INVxp67_ASAP7_75t_SL g496 ( .A(n_251), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g1354 ( .A(n_252), .Y(n_1354) );
INVx1_ASAP7_75t_L g1494 ( .A(n_253), .Y(n_1494) );
INVx1_ASAP7_75t_L g1032 ( .A(n_254), .Y(n_1032) );
AOI221xp5_ASAP7_75t_L g886 ( .A1(n_255), .A2(n_296), .B1(n_887), .B2(n_888), .C(n_889), .Y(n_886) );
INVxp33_ASAP7_75t_L g916 ( .A(n_255), .Y(n_916) );
INVx1_ASAP7_75t_L g1457 ( .A(n_256), .Y(n_1457) );
NAND2xp5_ASAP7_75t_L g1469 ( .A(n_256), .B(n_1466), .Y(n_1469) );
INVxp67_ASAP7_75t_SL g546 ( .A(n_258), .Y(n_546) );
XOR2x2_ASAP7_75t_L g765 ( .A(n_259), .B(n_766), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g1745 ( .A1(n_261), .A2(n_1746), .B1(n_1747), .B2(n_1748), .Y(n_1745) );
CKINVDCx5p33_ASAP7_75t_R g1746 ( .A(n_261), .Y(n_1746) );
INVxp33_ASAP7_75t_L g951 ( .A(n_262), .Y(n_951) );
AOI21xp33_ASAP7_75t_L g983 ( .A1(n_262), .A2(n_576), .B(n_984), .Y(n_983) );
INVx1_ASAP7_75t_L g654 ( .A(n_263), .Y(n_654) );
INVxp33_ASAP7_75t_L g784 ( .A(n_264), .Y(n_784) );
INVxp67_ASAP7_75t_SL g857 ( .A(n_265), .Y(n_857) );
CKINVDCx5p33_ASAP7_75t_R g1037 ( .A(n_266), .Y(n_1037) );
INVx1_ASAP7_75t_L g1191 ( .A(n_267), .Y(n_1191) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_269), .Y(n_346) );
INVxp33_ASAP7_75t_L g1155 ( .A(n_270), .Y(n_1155) );
AOI21xp5_ASAP7_75t_L g1210 ( .A1(n_271), .A2(n_389), .B(n_1211), .Y(n_1210) );
INVx1_ASAP7_75t_L g1240 ( .A(n_271), .Y(n_1240) );
INVxp67_ASAP7_75t_SL g544 ( .A(n_272), .Y(n_544) );
INVxp33_ASAP7_75t_L g952 ( .A(n_273), .Y(n_952) );
INVx1_ASAP7_75t_L g1089 ( .A(n_274), .Y(n_1089) );
AOI21xp5_ASAP7_75t_L g1104 ( .A1(n_274), .A2(n_846), .B(n_1105), .Y(n_1104) );
INVx2_ASAP7_75t_L g315 ( .A(n_275), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g1068 ( .A(n_276), .Y(n_1068) );
INVx1_ASAP7_75t_L g1168 ( .A(n_277), .Y(n_1168) );
XNOR2x1_ASAP7_75t_L g1394 ( .A(n_278), .B(n_1395), .Y(n_1394) );
XNOR2x2_ASAP7_75t_L g597 ( .A(n_279), .B(n_598), .Y(n_597) );
INVxp33_ASAP7_75t_L g1142 ( .A(n_280), .Y(n_1142) );
INVxp33_ASAP7_75t_SL g513 ( .A(n_281), .Y(n_513) );
INVx1_ASAP7_75t_L g717 ( .A(n_282), .Y(n_717) );
INVx1_ASAP7_75t_L g515 ( .A(n_283), .Y(n_515) );
INVxp33_ASAP7_75t_SL g927 ( .A(n_284), .Y(n_927) );
INVx1_ASAP7_75t_L g738 ( .A(n_285), .Y(n_738) );
INVx1_ASAP7_75t_L g1269 ( .A(n_286), .Y(n_1269) );
BUFx3_ASAP7_75t_L g343 ( .A(n_287), .Y(n_343) );
INVx1_ASAP7_75t_L g373 ( .A(n_287), .Y(n_373) );
BUFx3_ASAP7_75t_L g345 ( .A(n_288), .Y(n_345) );
INVx1_ASAP7_75t_L g355 ( .A(n_288), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g605 ( .A(n_289), .Y(n_605) );
INVxp33_ASAP7_75t_SL g685 ( .A(n_290), .Y(n_685) );
CKINVDCx5p33_ASAP7_75t_R g1353 ( .A(n_291), .Y(n_1353) );
CKINVDCx5p33_ASAP7_75t_R g1209 ( .A(n_292), .Y(n_1209) );
INVx1_ASAP7_75t_L g1225 ( .A(n_293), .Y(n_1225) );
CKINVDCx5p33_ASAP7_75t_R g1712 ( .A(n_295), .Y(n_1712) );
INVxp33_ASAP7_75t_L g914 ( .A(n_296), .Y(n_914) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_319), .B(n_1442), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_301), .B(n_306), .Y(n_300) );
AND2x4_ASAP7_75t_L g1739 ( .A(n_301), .B(n_307), .Y(n_1739) );
NOR2xp33_ASAP7_75t_SL g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_SL g1743 ( .A(n_302), .Y(n_1743) );
NAND2xp5_ASAP7_75t_L g1756 ( .A(n_302), .B(n_304), .Y(n_1756) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g1742 ( .A(n_304), .B(n_1743), .Y(n_1742) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_308), .B(n_312), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g469 ( .A(n_310), .B(n_318), .Y(n_469) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g521 ( .A(n_311), .B(n_522), .Y(n_521) );
OR2x6_ASAP7_75t_L g312 ( .A(n_313), .B(n_317), .Y(n_312) );
OR2x2_ASAP7_75t_L g329 ( .A(n_313), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g644 ( .A(n_313), .Y(n_644) );
INVx2_ASAP7_75t_SL g859 ( .A(n_313), .Y(n_859) );
BUFx6f_ASAP7_75t_L g926 ( .A(n_313), .Y(n_926) );
INVx2_ASAP7_75t_SL g960 ( .A(n_313), .Y(n_960) );
BUFx2_ASAP7_75t_L g1432 ( .A(n_313), .Y(n_1432) );
OAI22xp33_ASAP7_75t_L g1437 ( .A1(n_313), .A2(n_664), .B1(n_1407), .B2(n_1438), .Y(n_1437) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
AND2x2_ASAP7_75t_L g437 ( .A(n_315), .B(n_316), .Y(n_437) );
INVx2_ASAP7_75t_L g446 ( .A(n_315), .Y(n_446) );
AND2x4_ASAP7_75t_L g455 ( .A(n_315), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g462 ( .A(n_315), .Y(n_462) );
INVx1_ASAP7_75t_L g500 ( .A(n_315), .Y(n_500) );
INVx1_ASAP7_75t_L g448 ( .A(n_316), .Y(n_448) );
INVx2_ASAP7_75t_L g456 ( .A(n_316), .Y(n_456) );
INVx1_ASAP7_75t_L g494 ( .A(n_316), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_316), .B(n_446), .Y(n_527) );
INVx1_ASAP7_75t_L g649 ( .A(n_316), .Y(n_649) );
INVx2_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
OAI22xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_1053), .B1(n_1054), .B2(n_1441), .Y(n_319) );
INVx3_ASAP7_75t_L g1441 ( .A(n_320), .Y(n_1441) );
AO22x2_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_762), .B1(n_1051), .B2(n_1052), .Y(n_320) );
INVx1_ASAP7_75t_L g1052 ( .A(n_321), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_677), .B1(n_678), .B2(n_761), .Y(n_321) );
INVx2_ASAP7_75t_L g761 ( .A(n_322), .Y(n_761) );
AO22x2_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_503), .B1(n_504), .B2(n_676), .Y(n_322) );
INVx2_ASAP7_75t_SL g676 ( .A(n_323), .Y(n_676) );
XNOR2x1_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_430), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_346), .B(n_347), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g1270 ( .A1(n_327), .A2(n_425), .B1(n_1271), .B2(n_1283), .Y(n_1270) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx5_ASAP7_75t_L g727 ( .A(n_328), .Y(n_727) );
INVx1_ASAP7_75t_L g973 ( .A(n_328), .Y(n_973) );
INVx2_ASAP7_75t_L g1192 ( .A(n_328), .Y(n_1192) );
AND2x4_ASAP7_75t_L g328 ( .A(n_329), .B(n_332), .Y(n_328) );
INVx2_ASAP7_75t_L g516 ( .A(n_329), .Y(n_516) );
INVx3_ASAP7_75t_L g495 ( .A(n_330), .Y(n_495) );
INVx1_ASAP7_75t_L g831 ( .A(n_331), .Y(n_831) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x6_ASAP7_75t_L g825 ( .A(n_333), .B(n_826), .Y(n_825) );
AND2x4_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
AND2x4_ASAP7_75t_L g818 ( .A(n_334), .B(n_390), .Y(n_818) );
INVx2_ASAP7_75t_L g1311 ( .A(n_335), .Y(n_1311) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_341), .Y(n_335) );
AND2x4_ASAP7_75t_L g360 ( .A(n_336), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g365 ( .A(n_336), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g415 ( .A(n_336), .Y(n_415) );
BUFx2_ASAP7_75t_L g578 ( .A(n_336), .Y(n_578) );
AND2x4_ASAP7_75t_L g634 ( .A(n_336), .B(n_361), .Y(n_634) );
AND2x4_ASAP7_75t_L g636 ( .A(n_336), .B(n_366), .Y(n_636) );
NAND2x1p5_ASAP7_75t_L g795 ( .A(n_336), .B(n_487), .Y(n_795) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_336), .B(n_366), .Y(n_1204) );
AND2x4_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g390 ( .A(n_339), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g406 ( .A(n_340), .B(n_391), .Y(n_406) );
INVx1_ASAP7_75t_L g1066 ( .A(n_340), .Y(n_1066) );
HB1xp67_ASAP7_75t_L g1071 ( .A(n_340), .Y(n_1071) );
INVx1_ASAP7_75t_L g1075 ( .A(n_340), .Y(n_1075) );
INVx6_ASAP7_75t_L g411 ( .A(n_341), .Y(n_411) );
BUFx2_ASAP7_75t_L g576 ( .A(n_341), .Y(n_576) );
INVx2_ASAP7_75t_L g783 ( .A(n_341), .Y(n_783) );
AND2x4_ASAP7_75t_L g1069 ( .A(n_341), .B(n_1070), .Y(n_1069) );
AND2x4_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
INVx1_ASAP7_75t_L g367 ( .A(n_342), .Y(n_367) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g354 ( .A(n_343), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g397 ( .A(n_343), .B(n_345), .Y(n_397) );
INVx1_ASAP7_75t_L g363 ( .A(n_344), .Y(n_363) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g372 ( .A(n_345), .B(n_373), .Y(n_372) );
AOI31xp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_392), .A3(n_416), .B(n_424), .Y(n_347) );
AOI211xp5_ASAP7_75t_SL g348 ( .A1(n_349), .A2(n_350), .B(n_358), .C(n_368), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g976 ( .A1(n_350), .A2(n_965), .B(n_977), .Y(n_976) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_352), .Y(n_731) );
AOI221xp5_ASAP7_75t_L g885 ( .A1(n_352), .A2(n_886), .B1(n_890), .B2(n_893), .C(n_894), .Y(n_885) );
AOI221xp5_ASAP7_75t_L g1039 ( .A1(n_352), .A2(n_1027), .B1(n_1040), .B2(n_1041), .C(n_1043), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_352), .A2(n_418), .B1(n_1162), .B2(n_1167), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_352), .A2(n_418), .B1(n_1220), .B2(n_1221), .Y(n_1219) );
AND2x4_ASAP7_75t_L g352 ( .A(n_353), .B(n_356), .Y(n_352) );
INVx2_ASAP7_75t_SL g737 ( .A(n_353), .Y(n_737) );
BUFx3_ASAP7_75t_L g891 ( .A(n_353), .Y(n_891) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx2_ASAP7_75t_L g374 ( .A(n_354), .Y(n_374) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_354), .Y(n_561) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_354), .Y(n_567) );
INVx2_ASAP7_75t_SL g610 ( .A(n_354), .Y(n_610) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_354), .Y(n_630) );
BUFx3_ASAP7_75t_L g805 ( .A(n_354), .Y(n_805) );
BUFx2_ASAP7_75t_L g980 ( .A(n_354), .Y(n_980) );
AND2x6_ASAP7_75t_L g1093 ( .A(n_354), .B(n_1065), .Y(n_1093) );
HB1xp67_ASAP7_75t_L g1185 ( .A(n_354), .Y(n_1185) );
HB1xp67_ASAP7_75t_L g1401 ( .A(n_354), .Y(n_1401) );
INVx1_ASAP7_75t_L g381 ( .A(n_355), .Y(n_381) );
AND2x4_ASAP7_75t_L g395 ( .A(n_356), .B(n_396), .Y(n_395) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_356), .A2(n_583), .B(n_587), .Y(n_582) );
OAI21xp33_ASAP7_75t_L g625 ( .A1(n_356), .A2(n_626), .B(n_628), .Y(n_625) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_356), .B(n_630), .Y(n_1275) );
AOI222xp33_ASAP7_75t_L g1293 ( .A1(n_356), .A2(n_360), .B1(n_365), .B2(n_1294), .C1(n_1300), .C2(n_1301), .Y(n_1293) );
AOI221xp5_ASAP7_75t_L g1406 ( .A1(n_356), .A2(n_418), .B1(n_1407), .B2(n_1408), .C(n_1413), .Y(n_1406) );
A2O1A1Ixp33_ASAP7_75t_L g1730 ( .A1(n_356), .A2(n_887), .B(n_1731), .C(n_1732), .Y(n_1730) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g419 ( .A(n_357), .B(n_379), .Y(n_419) );
OR2x2_ASAP7_75t_L g422 ( .A(n_357), .B(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g774 ( .A(n_357), .B(n_439), .Y(n_774) );
A2O1A1Ixp33_ASAP7_75t_SL g1364 ( .A1(n_357), .A2(n_1365), .B(n_1368), .C(n_1372), .Y(n_1364) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_360), .A2(n_365), .B1(n_580), .B2(n_581), .Y(n_579) );
INVx2_ASAP7_75t_SL g733 ( .A(n_360), .Y(n_733) );
INVx2_ASAP7_75t_SL g895 ( .A(n_360), .Y(n_895) );
INVxp67_ASAP7_75t_L g987 ( .A(n_361), .Y(n_987) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g793 ( .A(n_362), .Y(n_793) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g1085 ( .A(n_363), .Y(n_1085) );
INVx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g735 ( .A(n_366), .Y(n_735) );
BUFx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x6_ASAP7_75t_L g1087 ( .A(n_367), .B(n_1066), .Y(n_1087) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI221xp5_ASAP7_75t_L g736 ( .A1(n_370), .A2(n_686), .B1(n_737), .B2(n_738), .C(n_739), .Y(n_736) );
INVx1_ASAP7_75t_L g1218 ( .A(n_370), .Y(n_1218) );
OAI22xp5_ASAP7_75t_L g1380 ( .A1(n_370), .A2(n_1381), .B1(n_1382), .B2(n_1383), .Y(n_1380) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_371), .Y(n_552) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_371), .Y(n_601) );
INVx1_ASAP7_75t_L g757 ( .A(n_371), .Y(n_757) );
INVx1_ASAP7_75t_L g999 ( .A(n_371), .Y(n_999) );
AND2x6_ASAP7_75t_L g1073 ( .A(n_371), .B(n_1074), .Y(n_1073) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g423 ( .A(n_372), .Y(n_423) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_372), .Y(n_612) );
INVx1_ASAP7_75t_L g778 ( .A(n_372), .Y(n_778) );
INVx1_ASAP7_75t_L g903 ( .A(n_372), .Y(n_903) );
INVx1_ASAP7_75t_L g380 ( .A(n_373), .Y(n_380) );
OAI21xp5_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_382), .B(n_383), .Y(n_375) );
OAI221xp5_ASAP7_75t_L g1133 ( .A1(n_376), .A2(n_1117), .B1(n_1118), .B2(n_1128), .C(n_1134), .Y(n_1133) );
OAI22xp5_ASAP7_75t_L g1375 ( .A1(n_376), .A2(n_1351), .B1(n_1353), .B2(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g584 ( .A(n_378), .Y(n_584) );
INVx2_ASAP7_75t_L g1126 ( .A(n_378), .Y(n_1126) );
INVx2_ASAP7_75t_L g1295 ( .A(n_378), .Y(n_1295) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g572 ( .A(n_379), .Y(n_572) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
AND2x2_ASAP7_75t_L g387 ( .A(n_380), .B(n_381), .Y(n_387) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI221xp5_ASAP7_75t_L g1377 ( .A1(n_385), .A2(n_405), .B1(n_1350), .B2(n_1354), .C(n_1378), .Y(n_1377) );
OAI221xp5_ASAP7_75t_L g1384 ( .A1(n_385), .A2(n_1126), .B1(n_1385), .B2(n_1386), .C(n_1387), .Y(n_1384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx2_ASAP7_75t_L g558 ( .A(n_387), .Y(n_558) );
BUFx4f_ASAP7_75t_L g570 ( .A(n_387), .Y(n_570) );
INVx2_ASAP7_75t_L g787 ( .A(n_387), .Y(n_787) );
INVx1_ASAP7_75t_L g1410 ( .A(n_387), .Y(n_1410) );
BUFx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_390), .Y(n_573) );
INVx2_ASAP7_75t_SL g617 ( .A(n_390), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g889 ( .A(n_390), .Y(n_889) );
INVx1_ASAP7_75t_L g984 ( .A(n_390), .Y(n_984) );
INVx1_ASAP7_75t_L g1095 ( .A(n_391), .Y(n_1095) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_398), .B1(n_399), .B2(n_407), .C(n_412), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx6f_ASAP7_75t_L g747 ( .A(n_395), .Y(n_747) );
AOI221xp5_ASAP7_75t_L g896 ( .A1(n_395), .A2(n_413), .B1(n_897), .B2(n_900), .C(n_904), .Y(n_896) );
INVx1_ASAP7_75t_L g990 ( .A(n_395), .Y(n_990) );
INVx1_ASAP7_75t_L g1183 ( .A(n_395), .Y(n_1183) );
INVx2_ASAP7_75t_SL g1214 ( .A(n_395), .Y(n_1214) );
BUFx3_ASAP7_75t_L g740 ( .A(n_396), .Y(n_740) );
BUFx6f_ASAP7_75t_L g807 ( .A(n_396), .Y(n_807) );
BUFx4f_ASAP7_75t_L g887 ( .A(n_396), .Y(n_887) );
INVx1_ASAP7_75t_L g1174 ( .A(n_396), .Y(n_1174) );
INVx2_ASAP7_75t_SL g1305 ( .A(n_396), .Y(n_1305) );
AND2x4_ASAP7_75t_L g1405 ( .A(n_396), .B(n_578), .Y(n_1405) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_397), .Y(n_403) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
A2O1A1Ixp33_ASAP7_75t_L g575 ( .A1(n_401), .A2(n_515), .B(n_576), .C(n_577), .Y(n_575) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x4_ASAP7_75t_L g413 ( .A(n_402), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g624 ( .A(n_402), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g1297 ( .A1(n_402), .A2(n_630), .B1(n_1298), .B2(n_1299), .Y(n_1297) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g753 ( .A(n_403), .Y(n_753) );
AND2x4_ASAP7_75t_L g1063 ( .A(n_403), .B(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx3_ASAP7_75t_L g899 ( .A(n_405), .Y(n_899) );
BUFx3_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_SL g563 ( .A(n_406), .Y(n_563) );
INVx1_ASAP7_75t_L g607 ( .A(n_406), .Y(n_607) );
INVx2_ASAP7_75t_L g802 ( .A(n_406), .Y(n_802) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g742 ( .A(n_410), .Y(n_742) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g555 ( .A(n_411), .Y(n_555) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_411), .Y(n_621) );
INVx1_ASAP7_75t_L g810 ( .A(n_411), .Y(n_810) );
INVx2_ASAP7_75t_L g1091 ( .A(n_411), .Y(n_1091) );
INVx2_ASAP7_75t_SL g1189 ( .A(n_411), .Y(n_1189) );
INVx2_ASAP7_75t_L g1211 ( .A(n_411), .Y(n_1211) );
HB1xp67_ASAP7_75t_L g1404 ( .A(n_411), .Y(n_1404) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g759 ( .A(n_413), .Y(n_759) );
AOI221xp5_ASAP7_75t_L g988 ( .A1(n_413), .A2(n_970), .B1(n_989), .B2(n_991), .C(n_996), .Y(n_988) );
AOI221xp5_ASAP7_75t_L g1045 ( .A1(n_413), .A2(n_747), .B1(n_1035), .B2(n_1046), .C(n_1047), .Y(n_1045) );
AOI221xp5_ASAP7_75t_L g1181 ( .A1(n_413), .A2(n_1168), .B1(n_1182), .B2(n_1184), .C(n_1186), .Y(n_1181) );
AOI221xp5_ASAP7_75t_L g1212 ( .A1(n_413), .A2(n_1213), .B1(n_1215), .B2(n_1216), .C(n_1217), .Y(n_1212) );
AOI221xp5_ASAP7_75t_L g1276 ( .A1(n_413), .A2(n_1213), .B1(n_1269), .B2(n_1277), .C(n_1278), .Y(n_1276) );
AOI21xp33_ASAP7_75t_L g1302 ( .A1(n_413), .A2(n_1303), .B(n_1306), .Y(n_1302) );
INVx1_ASAP7_75t_L g1372 ( .A(n_413), .Y(n_1372) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g734 ( .A(n_415), .B(n_735), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B1(n_420), .B2(n_421), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_418), .A2(n_421), .B1(n_717), .B2(n_719), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_418), .A2(n_421), .B1(n_906), .B2(n_907), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_418), .A2(n_421), .B1(n_966), .B2(n_968), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_418), .A2(n_421), .B1(n_1030), .B2(n_1032), .Y(n_1048) );
AOI22xp5_ASAP7_75t_L g1272 ( .A1(n_418), .A2(n_1265), .B1(n_1268), .B2(n_1273), .Y(n_1272) );
INVx6_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g1171 ( .A1(n_421), .A2(n_1165), .B1(n_1172), .B2(n_1175), .C(n_1178), .Y(n_1171) );
AOI211xp5_ASAP7_75t_L g1200 ( .A1(n_421), .A2(n_1201), .B(n_1202), .C(n_1205), .Y(n_1200) );
AOI221xp5_ASAP7_75t_L g1279 ( .A1(n_421), .A2(n_1266), .B1(n_1280), .B2(n_1281), .C(n_1282), .Y(n_1279) );
INVx4_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g586 ( .A(n_423), .Y(n_586) );
INVx2_ASAP7_75t_L g982 ( .A(n_423), .Y(n_982) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g1169 ( .A1(n_425), .A2(n_1170), .B1(n_1191), .B2(n_1192), .Y(n_1169) );
INVx5_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AOI31xp33_ASAP7_75t_L g729 ( .A1(n_426), .A2(n_730), .A3(n_744), .B(n_760), .Y(n_729) );
OAI31xp33_ASAP7_75t_L g833 ( .A1(n_426), .A2(n_834), .A3(n_853), .B(n_874), .Y(n_833) );
AOI31xp33_ASAP7_75t_L g1038 ( .A1(n_426), .A2(n_1039), .A3(n_1045), .B(n_1048), .Y(n_1038) );
AOI221x1_ASAP7_75t_SL g1059 ( .A1(n_426), .A2(n_1060), .B1(n_1094), .B2(n_1096), .C(n_1122), .Y(n_1059) );
BUFx8_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g883 ( .A(n_427), .Y(n_883) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx2_ASAP7_75t_L g638 ( .A(n_428), .Y(n_638) );
AND2x4_ASAP7_75t_L g1094 ( .A(n_428), .B(n_1095), .Y(n_1094) );
BUFx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g468 ( .A(n_429), .Y(n_468) );
OR2x6_ASAP7_75t_L g520 ( .A(n_429), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_431), .B(n_463), .Y(n_430) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_433), .A2(n_615), .B(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_433), .A2(n_685), .B1(n_686), .B2(n_687), .Y(n_684) );
BUFx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_434), .A2(n_518), .B(n_519), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_434), .A2(n_674), .B1(n_916), .B2(n_917), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_434), .A2(n_514), .B1(n_951), .B2(n_952), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_434), .A2(n_443), .B1(n_1013), .B2(n_1014), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_434), .A2(n_443), .B1(n_1146), .B2(n_1147), .Y(n_1145) );
AOI22xp33_ASAP7_75t_L g1239 ( .A1(n_434), .A2(n_1240), .B1(n_1241), .B2(n_1242), .Y(n_1239) );
AOI22xp33_ASAP7_75t_L g1252 ( .A1(n_434), .A2(n_1242), .B1(n_1253), .B2(n_1254), .Y(n_1252) );
NAND2xp5_ASAP7_75t_L g1707 ( .A(n_434), .B(n_1708), .Y(n_1707) );
AND2x4_ASAP7_75t_L g434 ( .A(n_435), .B(n_438), .Y(n_434) );
INVx2_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g472 ( .A(n_436), .Y(n_472) );
INVx2_ASAP7_75t_SL g832 ( .A(n_436), .Y(n_832) );
INVx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_437), .Y(n_536) );
AND2x2_ASAP7_75t_L g443 ( .A(n_438), .B(n_444), .Y(n_443) );
AND2x4_ASAP7_75t_L g452 ( .A(n_438), .B(n_453), .Y(n_452) );
AND2x6_ASAP7_75t_L g459 ( .A(n_438), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g514 ( .A(n_438), .B(n_444), .Y(n_514) );
AND2x2_ASAP7_75t_L g674 ( .A(n_438), .B(n_444), .Y(n_674) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_438), .B(n_444), .Y(n_1242) );
AOI22xp33_ASAP7_75t_L g1315 ( .A1(n_438), .A2(n_668), .B1(n_1316), .B2(n_1320), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_438), .B(n_444), .Y(n_1341) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_438), .B(n_1029), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_438), .B(n_832), .Y(n_1362) );
AND2x4_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
INVx1_ASAP7_75t_L g487 ( .A(n_439), .Y(n_487) );
INVx2_ASAP7_75t_L g838 ( .A(n_440), .Y(n_838) );
AND2x4_ASAP7_75t_L g855 ( .A(n_440), .B(n_536), .Y(n_855) );
AND2x2_ASAP7_75t_L g876 ( .A(n_440), .B(n_445), .Y(n_876) );
INVx1_ASAP7_75t_L g489 ( .A(n_441), .Y(n_489) );
INVx1_ASAP7_75t_L g522 ( .A(n_441), .Y(n_522) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g478 ( .A(n_445), .Y(n_478) );
BUFx6f_ASAP7_75t_L g1111 ( .A(n_445), .Y(n_1111) );
INVx1_ASAP7_75t_L g1322 ( .A(n_445), .Y(n_1322) );
INVx1_ASAP7_75t_L g1330 ( .A(n_445), .Y(n_1330) );
BUFx6f_ASAP7_75t_L g1704 ( .A(n_445), .Y(n_1704) );
AND2x4_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g699 ( .A(n_446), .Y(n_699) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .B1(n_457), .B2(n_458), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g1423 ( .A1(n_451), .A2(n_516), .B1(n_1424), .B2(n_1425), .Y(n_1423) );
BUFx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx2_ASAP7_75t_L g510 ( .A(n_452), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_452), .A2(n_459), .B1(n_614), .B2(n_671), .Y(n_670) );
BUFx2_ASAP7_75t_L g688 ( .A(n_452), .Y(n_688) );
BUFx2_ASAP7_75t_L g913 ( .A(n_452), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_452), .A2(n_459), .B1(n_1010), .B2(n_1011), .Y(n_1009) );
BUFx2_ASAP7_75t_L g1143 ( .A(n_452), .Y(n_1143) );
BUFx3_ASAP7_75t_L g937 ( .A(n_453), .Y(n_937) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_454), .Y(n_531) );
INVx3_ASAP7_75t_L g1029 ( .A(n_454), .Y(n_1029) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_455), .Y(n_475) );
INVx1_ASAP7_75t_L g871 ( .A(n_455), .Y(n_871) );
AND2x4_ASAP7_75t_L g461 ( .A(n_456), .B(n_462), .Y(n_461) );
INVxp67_ASAP7_75t_SL g683 ( .A(n_458), .Y(n_683) );
BUFx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_459), .A2(n_509), .B1(n_510), .B2(n_511), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_459), .A2(n_912), .B1(n_913), .B2(n_914), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_459), .A2(n_688), .B1(n_948), .B2(n_949), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g1141 ( .A1(n_459), .A2(n_1142), .B1(n_1143), .B2(n_1144), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_459), .A2(n_913), .B1(n_1209), .B2(n_1238), .Y(n_1237) );
AOI22xp33_ASAP7_75t_L g1249 ( .A1(n_459), .A2(n_913), .B1(n_1250), .B2(n_1251), .Y(n_1249) );
INVx1_ASAP7_75t_SL g1342 ( .A(n_459), .Y(n_1342) );
AOI22xp5_ASAP7_75t_L g1420 ( .A1(n_459), .A2(n_1242), .B1(n_1421), .B2(n_1422), .Y(n_1420) );
AOI22xp33_ASAP7_75t_L g1710 ( .A1(n_459), .A2(n_1341), .B1(n_1711), .B2(n_1712), .Y(n_1710) );
NAND2x1p5_ASAP7_75t_L g700 ( .A(n_460), .B(n_495), .Y(n_700) );
BUFx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx2_ASAP7_75t_L g480 ( .A(n_461), .Y(n_480) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_461), .Y(n_539) );
BUFx3_ASAP7_75t_L g549 ( .A(n_461), .Y(n_549) );
BUFx6f_ASAP7_75t_L g844 ( .A(n_461), .Y(n_844) );
INVx1_ASAP7_75t_L g1114 ( .A(n_461), .Y(n_1114) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_464), .B(n_491), .Y(n_463) );
AOI33xp33_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_470), .A3(n_476), .B1(n_481), .B2(n_482), .B3(n_483), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
BUFx2_ASAP7_75t_L g591 ( .A(n_468), .Y(n_591) );
OR2x6_ASAP7_75t_L g801 ( .A(n_468), .B(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g827 ( .A(n_468), .Y(n_827) );
AOI31xp33_ASAP7_75t_L g975 ( .A1(n_468), .A2(n_976), .A3(n_988), .B(n_1000), .Y(n_975) );
AND2x4_ASAP7_75t_L g1228 ( .A(n_468), .B(n_469), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1706 ( .A(n_468), .B(n_847), .Y(n_1706) );
INVx1_ASAP7_75t_L g862 ( .A(n_469), .Y(n_862) );
BUFx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_474), .A2(n_1019), .B1(n_1020), .B2(n_1021), .Y(n_1018) );
OAI22xp5_ASAP7_75t_L g1260 ( .A1(n_474), .A2(n_1158), .B1(n_1261), .B2(n_1262), .Y(n_1260) );
OAI22xp5_ASAP7_75t_L g1263 ( .A1(n_474), .A2(n_1264), .B1(n_1265), .B2(n_1266), .Y(n_1263) );
OAI22xp5_ASAP7_75t_L g1349 ( .A1(n_474), .A2(n_712), .B1(n_1350), .B2(n_1351), .Y(n_1349) );
INVx4_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_SL g545 ( .A(n_475), .Y(n_545) );
INVx2_ASAP7_75t_SL g707 ( .A(n_475), .Y(n_707) );
INVx2_ASAP7_75t_SL g841 ( .A(n_475), .Y(n_841) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x4_ASAP7_75t_L g502 ( .A(n_480), .B(n_495), .Y(n_502) );
INVx1_ASAP7_75t_L g723 ( .A(n_483), .Y(n_723) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_484), .A2(n_520), .B1(n_523), .B2(n_540), .Y(n_519) );
OAI33xp33_ASAP7_75t_L g922 ( .A1(n_484), .A2(n_520), .A3(n_923), .B1(n_929), .B2(n_935), .B3(n_938), .Y(n_922) );
OAI33xp33_ASAP7_75t_L g1017 ( .A1(n_484), .A2(n_520), .A3(n_1018), .B1(n_1022), .B2(n_1026), .B3(n_1031), .Y(n_1017) );
OAI33xp33_ASAP7_75t_L g1149 ( .A1(n_484), .A2(n_1150), .A3(n_1151), .B1(n_1156), .B2(n_1161), .B3(n_1166), .Y(n_1149) );
OAI33xp33_ASAP7_75t_L g1256 ( .A1(n_484), .A2(n_1150), .A3(n_1257), .B1(n_1260), .B2(n_1263), .B3(n_1267), .Y(n_1256) );
CKINVDCx8_ASAP7_75t_R g484 ( .A(n_485), .Y(n_484) );
INVx5_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx6_ASAP7_75t_L g668 ( .A(n_486), .Y(n_668) );
OR2x6_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx2_ASAP7_75t_L g847 ( .A(n_488), .Y(n_847) );
NAND2x1p5_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
AOI221xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_496), .B1(n_497), .B2(n_501), .C(n_502), .Y(n_491) );
INVx1_ASAP7_75t_L g596 ( .A(n_492), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g1224 ( .A1(n_492), .A2(n_497), .B1(n_502), .B2(n_1225), .C(n_1226), .Y(n_1224) );
AOI221xp5_ASAP7_75t_L g1335 ( .A1(n_492), .A2(n_497), .B1(n_502), .B2(n_1300), .C(n_1301), .Y(n_1335) );
AOI221xp5_ASAP7_75t_L g1417 ( .A1(n_492), .A2(n_497), .B1(n_502), .B2(n_1418), .C(n_1419), .Y(n_1417) );
AOI221xp5_ASAP7_75t_L g1697 ( .A1(n_492), .A2(n_497), .B1(n_502), .B2(n_1698), .C(n_1699), .Y(n_1697) );
AND2x4_ASAP7_75t_L g492 ( .A(n_493), .B(n_495), .Y(n_492) );
AND2x2_ASAP7_75t_L g850 ( .A(n_493), .B(n_829), .Y(n_850) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g694 ( .A(n_494), .Y(n_694) );
AND2x4_ASAP7_75t_L g497 ( .A(n_495), .B(n_498), .Y(n_497) );
NAND2x1_ASAP7_75t_SL g692 ( .A(n_495), .B(n_693), .Y(n_692) );
NAND2x1p5_ASAP7_75t_L g697 ( .A(n_495), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g594 ( .A(n_497), .Y(n_594) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g648 ( .A(n_500), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_500), .B(n_649), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g592 ( .A1(n_502), .A2(n_580), .B1(n_581), .B2(n_593), .C(n_595), .Y(n_592) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_502), .A2(n_593), .B1(n_595), .B2(n_635), .C(n_637), .Y(n_675) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
XOR2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_597), .Y(n_504) );
NAND4xp25_ASAP7_75t_L g506 ( .A(n_507), .B(n_517), .C(n_550), .D(n_592), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_512), .Y(n_507) );
OAI221xp5_ASAP7_75t_L g568 ( .A1(n_511), .A2(n_518), .B1(n_569), .B2(n_571), .C(n_573), .Y(n_568) );
AOI22xp33_ASAP7_75t_SL g512 ( .A1(n_513), .A2(n_514), .B1(n_515), .B2(n_516), .Y(n_512) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_516), .A2(n_622), .B1(n_673), .B2(n_674), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g1327 ( .A1(n_516), .A2(n_1228), .B1(n_1312), .B2(n_1328), .Y(n_1327) );
AOI22xp33_ASAP7_75t_L g1713 ( .A1(n_516), .A2(n_1345), .B1(n_1714), .B2(n_1715), .Y(n_1713) );
OAI33xp33_ASAP7_75t_L g640 ( .A1(n_520), .A2(n_641), .A3(n_650), .B1(n_655), .B2(n_660), .B3(n_667), .Y(n_640) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_520), .Y(n_702) );
HB1xp67_ASAP7_75t_L g1150 ( .A(n_520), .Y(n_1150) );
OAI221xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_528), .B1(n_529), .B2(n_532), .C(n_533), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g1355 ( .A1(n_524), .A2(n_1028), .B1(n_1356), .B2(n_1357), .Y(n_1355) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g543 ( .A(n_527), .Y(n_543) );
INVx1_ASAP7_75t_L g653 ( .A(n_527), .Y(n_653) );
OAI221xp5_ASAP7_75t_L g556 ( .A1(n_528), .A2(n_557), .B1(n_559), .B2(n_560), .C(n_562), .Y(n_556) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_531), .A2(n_605), .B1(n_651), .B2(n_654), .Y(n_650) );
INVx3_ASAP7_75t_L g658 ( .A(n_531), .Y(n_658) );
INVx2_ASAP7_75t_L g1101 ( .A(n_531), .Y(n_1101) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_SL g845 ( .A(n_535), .Y(n_845) );
INVx2_ASAP7_75t_L g1105 ( .A(n_535), .Y(n_1105) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx6f_ASAP7_75t_L g1230 ( .A(n_536), .Y(n_1230) );
AOI22xp5_ASAP7_75t_L g1317 ( .A1(n_537), .A2(n_1230), .B1(n_1318), .B2(n_1319), .Y(n_1317) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g1231 ( .A(n_538), .Y(n_1231) );
INVx2_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
OAI221xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_544), .B1(n_545), .B2(n_546), .C(n_547), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_541), .A2(n_656), .B1(n_657), .B2(n_659), .Y(n_655) );
BUFx2_ASAP7_75t_L g964 ( .A(n_541), .Y(n_964) );
INVx2_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g712 ( .A(n_542), .Y(n_712) );
INVx2_ASAP7_75t_L g840 ( .A(n_542), .Y(n_840) );
BUFx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g933 ( .A(n_543), .Y(n_933) );
OAI22xp5_ASAP7_75t_SL g929 ( .A1(n_545), .A2(n_930), .B1(n_931), .B2(n_934), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_545), .A2(n_964), .B1(n_965), .B2(n_966), .Y(n_963) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x4_ASAP7_75t_L g836 ( .A(n_549), .B(n_837), .Y(n_836) );
OAI31xp33_ASAP7_75t_SL g550 ( .A1(n_551), .A2(n_564), .A3(n_574), .B(n_590), .Y(n_550) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
HB1xp67_ASAP7_75t_L g997 ( .A(n_555), .Y(n_997) );
OAI21xp5_ASAP7_75t_SL g1208 ( .A1(n_557), .A2(n_1209), .B(n_1210), .Y(n_1208) );
INVx2_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g603 ( .A(n_558), .Y(n_603) );
OAI221xp5_ASAP7_75t_L g602 ( .A1(n_560), .A2(n_603), .B1(n_604), .B2(n_605), .C(n_606), .Y(n_602) );
INVx1_ASAP7_75t_L g1176 ( .A(n_560), .Y(n_1176) );
INVx2_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
BUFx3_ASAP7_75t_L g1379 ( .A(n_561), .Y(n_1379) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
BUFx2_ASAP7_75t_L g754 ( .A(n_563), .Y(n_754) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g588 ( .A(n_567), .Y(n_588) );
BUFx2_ASAP7_75t_L g749 ( .A(n_567), .Y(n_749) );
BUFx3_ASAP7_75t_L g815 ( .A(n_567), .Y(n_815) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_SL g589 ( .A(n_570), .Y(n_589) );
INVx1_ASAP7_75t_L g1721 ( .A(n_570), .Y(n_1721) );
OAI221xp5_ASAP7_75t_L g613 ( .A1(n_571), .A2(n_589), .B1(n_614), .B2(n_615), .C(n_616), .Y(n_613) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND3xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_579), .C(n_582), .Y(n_574) );
A2O1A1Ixp33_ASAP7_75t_SL g619 ( .A1(n_577), .A2(n_620), .B(n_622), .C(n_623), .Y(n_619) );
BUFx3_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g1206 ( .A(n_588), .Y(n_1206) );
OAI31xp33_ASAP7_75t_L g1363 ( .A1(n_590), .A2(n_1364), .A3(n_1373), .B(n_1374), .Y(n_1363) );
CKINVDCx8_ASAP7_75t_R g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND4xp25_ASAP7_75t_L g598 ( .A(n_599), .B(n_639), .C(n_669), .D(n_675), .Y(n_598) );
OAI31xp33_ASAP7_75t_SL g599 ( .A1(n_600), .A2(n_608), .A3(n_618), .B(n_638), .Y(n_599) );
INVx2_ASAP7_75t_SL g1412 ( .A(n_601), .Y(n_1412) );
OAI22xp33_ASAP7_75t_L g641 ( .A1(n_604), .A2(n_642), .B1(n_643), .B2(n_645), .Y(n_641) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g772 ( .A(n_610), .Y(n_772) );
BUFx3_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g627 ( .A(n_612), .Y(n_627) );
INVx1_ASAP7_75t_L g817 ( .A(n_612), .Y(n_817) );
BUFx6f_ASAP7_75t_L g892 ( .A(n_612), .Y(n_892) );
INVx1_ASAP7_75t_L g743 ( .A(n_616), .Y(n_743) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND3xp33_ASAP7_75t_SL g618 ( .A(n_619), .B(n_625), .C(n_631), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g813 ( .A(n_621), .Y(n_813) );
INVx4_ASAP7_75t_L g888 ( .A(n_621), .Y(n_888) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g898 ( .A(n_624), .Y(n_898) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_635), .B1(n_636), .B2(n_637), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx4_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g1179 ( .A(n_634), .Y(n_1179) );
INVx1_ASAP7_75t_SL g1414 ( .A(n_634), .Y(n_1414) );
AOI22xp33_ASAP7_75t_L g1733 ( .A1(n_634), .A2(n_636), .B1(n_1698), .B2(n_1699), .Y(n_1733) );
INVx2_ASAP7_75t_SL g1044 ( .A(n_636), .Y(n_1044) );
INVx2_ASAP7_75t_L g1180 ( .A(n_636), .Y(n_1180) );
AOI22xp5_ASAP7_75t_L g1198 ( .A1(n_638), .A2(n_727), .B1(n_1199), .B2(n_1222), .Y(n_1198) );
INVx2_ASAP7_75t_L g1415 ( .A(n_638), .Y(n_1415) );
OAI31xp33_ASAP7_75t_L g1716 ( .A1(n_638), .A2(n_1717), .A3(n_1718), .B(n_1729), .Y(n_1716) );
OAI22xp33_ASAP7_75t_L g660 ( .A1(n_643), .A2(n_661), .B1(n_662), .B2(n_666), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g1352 ( .A1(n_643), .A2(n_721), .B1(n_1353), .B2(n_1354), .Y(n_1352) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g705 ( .A(n_644), .Y(n_705) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g1103 ( .A(n_646), .Y(n_1103) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g873 ( .A(n_647), .B(n_830), .Y(n_873) );
HB1xp67_ASAP7_75t_L g969 ( .A(n_647), .Y(n_969) );
OR2x6_ASAP7_75t_L g1099 ( .A(n_647), .B(n_830), .Y(n_1099) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g928 ( .A(n_648), .Y(n_928) );
BUFx2_ASAP7_75t_L g940 ( .A(n_648), .Y(n_940) );
INVx3_ASAP7_75t_L g1034 ( .A(n_648), .Y(n_1034) );
BUFx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
HB1xp67_ASAP7_75t_L g865 ( .A(n_653), .Y(n_865) );
INVx2_ASAP7_75t_L g1159 ( .A(n_653), .Y(n_1159) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g714 ( .A(n_663), .Y(n_714) );
INVx1_ASAP7_75t_L g1024 ( .A(n_663), .Y(n_1024) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
BUFx3_ASAP7_75t_L g721 ( .A(n_664), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g1430 ( .A1(n_664), .A2(n_1431), .B1(n_1432), .B2(n_1433), .Y(n_1430) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g971 ( .A(n_668), .Y(n_971) );
AOI33xp33_ASAP7_75t_L g1227 ( .A1(n_668), .A2(n_1228), .A3(n_1229), .B1(n_1232), .B2(n_1233), .B3(n_1236), .Y(n_1227) );
AOI222xp33_ASAP7_75t_L g1426 ( .A1(n_668), .A2(n_1228), .B1(n_1362), .B2(n_1427), .C1(n_1428), .C2(n_1434), .Y(n_1426) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .Y(n_669) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
XNOR2x1_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_724), .Y(n_680) );
NOR3xp33_ASAP7_75t_SL g681 ( .A(n_682), .B(n_689), .C(n_701), .Y(n_681) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_SL g919 ( .A(n_691), .Y(n_919) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND2x1p5_ASAP7_75t_L g1107 ( .A(n_693), .B(n_1108), .Y(n_1107) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
BUFx4f_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
BUFx4f_ASAP7_75t_L g920 ( .A(n_697), .Y(n_920) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OR2x6_ASAP7_75t_L g852 ( .A(n_699), .B(n_830), .Y(n_852) );
BUFx3_ASAP7_75t_L g921 ( .A(n_700), .Y(n_921) );
BUFx2_ASAP7_75t_L g1016 ( .A(n_700), .Y(n_1016) );
OAI33xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .A3(n_708), .B1(n_715), .B2(n_718), .B3(n_723), .Y(n_701) );
OAI33xp33_ASAP7_75t_L g954 ( .A1(n_702), .A2(n_955), .A3(n_958), .B1(n_963), .B2(n_967), .B3(n_971), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_705), .B1(n_706), .B2(n_707), .Y(n_703) );
OAI22xp33_ASAP7_75t_L g718 ( .A1(n_705), .A2(n_719), .B1(n_720), .B2(n_722), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_707), .A2(n_710), .B1(n_716), .B2(n_717), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g1156 ( .A1(n_707), .A2(n_1157), .B1(n_1158), .B2(n_1160), .Y(n_1156) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_710), .B1(n_713), .B2(n_714), .Y(n_708) );
OAI22xp33_ASAP7_75t_SL g958 ( .A1(n_710), .A2(n_959), .B1(n_961), .B2(n_962), .Y(n_958) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g1161 ( .A1(n_712), .A2(n_1162), .B1(n_1163), .B2(n_1165), .Y(n_1161) );
OAI22xp33_ASAP7_75t_L g955 ( .A1(n_714), .A2(n_841), .B1(n_956), .B2(n_957), .Y(n_955) );
OAI22xp33_ASAP7_75t_L g1267 ( .A1(n_714), .A2(n_1152), .B1(n_1268), .B2(n_1269), .Y(n_1267) );
OAI22xp5_ASAP7_75t_SL g1358 ( .A1(n_714), .A2(n_926), .B1(n_1359), .B2(n_1360), .Y(n_1358) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_716), .A2(n_731), .B(n_732), .Y(n_730) );
OAI221xp5_ASAP7_75t_L g856 ( .A1(n_720), .A2(n_857), .B1(n_858), .B2(n_860), .C(n_861), .Y(n_856) );
BUFx3_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g744 ( .A1(n_722), .A2(n_745), .B1(n_748), .B2(n_755), .C(n_758), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_728), .B(n_729), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_727), .A2(n_883), .B1(n_884), .B2(n_908), .Y(n_882) );
AOI21xp33_ASAP7_75t_SL g1036 ( .A1(n_727), .A2(n_1037), .B(n_1038), .Y(n_1036) );
OR2x6_ASAP7_75t_L g798 ( .A(n_735), .B(n_795), .Y(n_798) );
INVx1_ASAP7_75t_L g992 ( .A(n_737), .Y(n_992) );
INVx1_ASAP7_75t_L g1042 ( .A(n_737), .Y(n_1042) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx3_ASAP7_75t_L g1080 ( .A(n_753), .Y(n_1080) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g1051 ( .A(n_762), .Y(n_1051) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_764), .B1(n_1003), .B2(n_1049), .Y(n_762) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
XNOR2x1_ASAP7_75t_L g764 ( .A(n_765), .B(n_879), .Y(n_764) );
NAND3xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_823), .C(n_833), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_788), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_779), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_771), .B1(n_775), .B2(n_776), .Y(n_769) );
OAI221xp5_ASAP7_75t_L g839 ( .A1(n_770), .A2(n_775), .B1(n_840), .B2(n_841), .C(n_842), .Y(n_839) );
AND2x2_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
AND2x2_ASAP7_75t_L g781 ( .A(n_773), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OR2x6_ASAP7_75t_L g777 ( .A(n_774), .B(n_778), .Y(n_777) );
OR2x6_ASAP7_75t_L g786 ( .A(n_774), .B(n_787), .Y(n_786) );
CKINVDCx6p67_ASAP7_75t_R g776 ( .A(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g1367 ( .A(n_778), .Y(n_1367) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_781), .B1(n_784), .B2(n_785), .Y(n_779) );
INVx2_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g901 ( .A(n_783), .Y(n_901) );
CKINVDCx6p67_ASAP7_75t_R g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g1129 ( .A(n_787), .Y(n_1129) );
BUFx3_ASAP7_75t_L g1725 ( .A(n_787), .Y(n_1725) );
NAND3xp33_ASAP7_75t_SL g788 ( .A(n_789), .B(n_799), .C(n_819), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_791), .B1(n_796), .B2(n_797), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_790), .A2(n_796), .B1(n_849), .B2(n_851), .Y(n_848) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
NAND2x1p5_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .Y(n_792) );
INVx2_ASAP7_75t_SL g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g822 ( .A(n_795), .Y(n_822) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
AOI33xp33_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_803), .A3(n_808), .B1(n_811), .B2(n_814), .B3(n_818), .Y(n_799) );
CKINVDCx5p33_ASAP7_75t_R g800 ( .A(n_801), .Y(n_800) );
INVx2_ASAP7_75t_L g1124 ( .A(n_801), .Y(n_1124) );
INVx1_ASAP7_75t_L g995 ( .A(n_802), .Y(n_995) );
BUFx3_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx2_ASAP7_75t_SL g1370 ( .A(n_805), .Y(n_1370) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_807), .B(n_822), .Y(n_821) );
BUFx2_ASAP7_75t_SL g1371 ( .A(n_807), .Y(n_1371) );
BUFx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
HB1xp67_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx4_ASAP7_75t_L g1132 ( .A(n_818), .Y(n_1132) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
NOR2xp67_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
INVx2_ASAP7_75t_L g1313 ( .A(n_827), .Y(n_1313) );
INVx1_ASAP7_75t_L g1116 ( .A(n_828), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_829), .B(n_832), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g1108 ( .A(n_830), .Y(n_1108) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx8_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
AOI222xp33_ASAP7_75t_L g1115 ( .A1(n_836), .A2(n_855), .B1(n_1068), .B2(n_1116), .C1(n_1117), .C2(n_1118), .Y(n_1115) );
AND2x4_ASAP7_75t_L g878 ( .A(n_837), .B(n_870), .Y(n_878) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVxp67_ASAP7_75t_L g1331 ( .A(n_841), .Y(n_1331) );
BUFx6f_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx2_ASAP7_75t_SL g846 ( .A(n_847), .Y(n_846) );
HB1xp67_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
CKINVDCx11_ASAP7_75t_R g851 ( .A(n_852), .Y(n_851) );
CKINVDCx6p67_ASAP7_75t_R g854 ( .A(n_855), .Y(n_854) );
OAI22xp33_ASAP7_75t_L g1022 ( .A1(n_858), .A2(n_1023), .B1(n_1024), .B2(n_1025), .Y(n_1022) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx2_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_866), .B1(n_867), .B2(n_872), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx3_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_876), .A2(n_878), .B1(n_1120), .B2(n_1121), .Y(n_1119) );
INVx3_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
AO22x2_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_942), .B1(n_1001), .B2(n_1002), .Y(n_879) );
INVx1_ASAP7_75t_L g1002 ( .A(n_880), .Y(n_1002) );
XOR2x2_ASAP7_75t_L g880 ( .A(n_881), .B(n_941), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_882), .B(n_909), .Y(n_881) );
NAND3xp33_ASAP7_75t_L g884 ( .A(n_885), .B(n_896), .C(n_905), .Y(n_884) );
BUFx2_ASAP7_75t_L g993 ( .A(n_887), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g1365 ( .A1(n_888), .A2(n_1357), .B1(n_1359), .B2(n_1366), .Y(n_1365) );
INVxp67_ASAP7_75t_L g1382 ( .A(n_891), .Y(n_1382) );
INVx1_ASAP7_75t_L g1376 ( .A(n_892), .Y(n_1376) );
OAI22xp5_ASAP7_75t_L g935 ( .A1(n_893), .A2(n_907), .B1(n_931), .B2(n_936), .Y(n_935) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx1_ASAP7_75t_L g1177 ( .A(n_903), .Y(n_1177) );
INVx1_ASAP7_75t_L g1207 ( .A(n_903), .Y(n_1207) );
OAI22xp33_ASAP7_75t_L g938 ( .A1(n_904), .A2(n_906), .B1(n_925), .B2(n_939), .Y(n_938) );
NOR3xp33_ASAP7_75t_L g909 ( .A(n_910), .B(n_918), .C(n_922), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_911), .B(n_915), .Y(n_910) );
OAI22xp33_ASAP7_75t_L g923 ( .A1(n_924), .A2(n_925), .B1(n_927), .B2(n_928), .Y(n_923) );
BUFx2_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
OAI22xp33_ASAP7_75t_L g967 ( .A1(n_926), .A2(n_968), .B1(n_969), .B2(n_970), .Y(n_967) );
INVx1_ASAP7_75t_L g1153 ( .A(n_926), .Y(n_1153) );
OAI22xp33_ASAP7_75t_L g1325 ( .A1(n_926), .A2(n_1034), .B1(n_1299), .B2(n_1326), .Y(n_1325) );
OAI22xp5_ASAP7_75t_L g1332 ( .A1(n_926), .A2(n_1034), .B1(n_1333), .B2(n_1334), .Y(n_1332) );
INVx2_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx2_ASAP7_75t_L g1020 ( .A(n_932), .Y(n_1020) );
INVx2_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
BUFx2_ASAP7_75t_L g1264 ( .A(n_933), .Y(n_1264) );
CKINVDCx5p33_ASAP7_75t_R g936 ( .A(n_937), .Y(n_936) );
INVx2_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g1001 ( .A(n_942), .Y(n_1001) );
XNOR2xp5_ASAP7_75t_L g942 ( .A(n_943), .B(n_944), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_945), .B(n_972), .Y(n_944) );
NOR3xp33_ASAP7_75t_SL g945 ( .A(n_946), .B(n_953), .C(n_954), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_947), .B(n_950), .Y(n_946) );
OAI22xp33_ASAP7_75t_L g1031 ( .A1(n_959), .A2(n_1032), .B1(n_1033), .B2(n_1035), .Y(n_1031) );
INVx3_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
AOI21xp5_ASAP7_75t_L g972 ( .A1(n_973), .A2(n_974), .B(n_975), .Y(n_972) );
INVx1_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
AOI31xp33_ASAP7_75t_L g978 ( .A1(n_979), .A2(n_983), .A3(n_985), .B(n_986), .Y(n_978) );
INVx1_ASAP7_75t_L g1411 ( .A(n_980), .Y(n_1411) );
INVx1_ASAP7_75t_L g1296 ( .A(n_981), .Y(n_1296) );
BUFx2_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVx2_ASAP7_75t_L g1136 ( .A(n_982), .Y(n_1136) );
INVx1_ASAP7_75t_L g1387 ( .A(n_984), .Y(n_1387) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
INVx1_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
BUFx2_ASAP7_75t_SL g1004 ( .A(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1005), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1036), .Y(n_1006) );
NOR3xp33_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1015), .C(n_1017), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1012), .Y(n_1008) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_1020), .A2(n_1027), .B1(n_1028), .B2(n_1030), .Y(n_1026) );
INVx2_ASAP7_75t_L g1436 ( .A(n_1028), .Y(n_1436) );
INVx2_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
INVx2_ASAP7_75t_L g1164 ( .A(n_1029), .Y(n_1164) );
INVx2_ASAP7_75t_L g1235 ( .A(n_1029), .Y(n_1235) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1029), .Y(n_1324) );
OAI22xp33_ASAP7_75t_L g1151 ( .A1(n_1033), .A2(n_1152), .B1(n_1154), .B2(n_1155), .Y(n_1151) );
OAI22xp33_ASAP7_75t_L g1166 ( .A1(n_1033), .A2(n_1152), .B1(n_1167), .B2(n_1168), .Y(n_1166) );
OAI22xp33_ASAP7_75t_L g1257 ( .A1(n_1033), .A2(n_1152), .B1(n_1258), .B2(n_1259), .Y(n_1257) );
BUFx2_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
OAI22xp5_ASAP7_75t_L g1054 ( .A1(n_1055), .A2(n_1284), .B1(n_1285), .B2(n_1440), .Y(n_1054) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1055), .Y(n_1440) );
XNOR2xp5_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1194), .Y(n_1055) );
AO22x2_ASAP7_75t_L g1056 ( .A1(n_1057), .A2(n_1058), .B1(n_1137), .B2(n_1193), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
NAND4xp25_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1067), .C(n_1076), .D(n_1088), .Y(n_1060) );
BUFx2_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
INVx5_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_1068), .A2(n_1069), .B1(n_1072), .B2(n_1073), .Y(n_1067) );
AND2x4_ASAP7_75t_L g1083 ( .A(n_1070), .B(n_1084), .Y(n_1083) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
AND2x4_ASAP7_75t_L g1090 ( .A(n_1074), .B(n_1091), .Y(n_1090) );
INVx1_ASAP7_75t_SL g1074 ( .A(n_1075), .Y(n_1074) );
AOI222xp33_ASAP7_75t_L g1076 ( .A1(n_1077), .A2(n_1078), .B1(n_1081), .B2(n_1082), .C1(n_1086), .C2(n_1087), .Y(n_1076) );
OAI21xp5_ASAP7_75t_SL g1102 ( .A1(n_1077), .A2(n_1103), .B(n_1104), .Y(n_1102) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
BUFx4f_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_1089), .A2(n_1090), .B1(n_1092), .B2(n_1093), .Y(n_1088) );
NAND3xp33_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1115), .C(n_1119), .Y(n_1096) );
NOR3xp33_ASAP7_75t_SL g1097 ( .A(n_1098), .B(n_1100), .C(n_1106), .Y(n_1097) );
INVx2_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1112), .Y(n_1109) );
INVx2_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
OAI22xp5_ASAP7_75t_L g1122 ( .A1(n_1123), .A2(n_1125), .B1(n_1132), .B2(n_1133), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
OAI221xp5_ASAP7_75t_L g1125 ( .A1(n_1126), .A2(n_1127), .B1(n_1128), .B2(n_1130), .C(n_1131), .Y(n_1125) );
INVx2_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1137), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1169), .Y(n_1138) );
NOR3xp33_ASAP7_75t_SL g1139 ( .A(n_1140), .B(n_1148), .C(n_1149), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1145), .Y(n_1140) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
BUFx2_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
HB1xp67_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
INVx2_ASAP7_75t_L g1429 ( .A(n_1164), .Y(n_1429) );
NAND3xp33_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1181), .C(n_1190), .Y(n_1170) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
INVx2_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
XOR2x2_ASAP7_75t_L g1195 ( .A(n_1196), .B(n_1244), .Y(n_1195) );
XNOR2xp5_ASAP7_75t_L g1196 ( .A(n_1197), .B(n_1243), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1223), .Y(n_1197) );
NAND3xp33_ASAP7_75t_SL g1199 ( .A(n_1200), .B(n_1212), .C(n_1219), .Y(n_1199) );
INVx2_ASAP7_75t_SL g1203 ( .A(n_1204), .Y(n_1203) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
AND4x1_ASAP7_75t_L g1223 ( .A(n_1224), .B(n_1227), .C(n_1237), .D(n_1239), .Y(n_1223) );
AOI33xp33_ASAP7_75t_L g1700 ( .A1(n_1228), .A2(n_1701), .A3(n_1702), .B1(n_1703), .B2(n_1705), .B3(n_1706), .Y(n_1700) );
INVx2_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
XNOR2x1_ASAP7_75t_L g1244 ( .A(n_1245), .B(n_1246), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1247), .B(n_1270), .Y(n_1246) );
NOR3xp33_ASAP7_75t_L g1247 ( .A(n_1248), .B(n_1255), .C(n_1256), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1249), .B(n_1252), .Y(n_1248) );
NAND3xp33_ASAP7_75t_L g1271 ( .A(n_1272), .B(n_1276), .C(n_1279), .Y(n_1271) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
OAI22xp5_ASAP7_75t_L g1285 ( .A1(n_1286), .A2(n_1287), .B1(n_1393), .B2(n_1439), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
AOI22xp5_ASAP7_75t_L g1287 ( .A1(n_1288), .A2(n_1336), .B1(n_1390), .B2(n_1391), .Y(n_1287) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1288), .Y(n_1390) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
XNOR2x1_ASAP7_75t_L g1289 ( .A(n_1290), .B(n_1291), .Y(n_1289) );
OAI22xp5_ASAP7_75t_L g1450 ( .A1(n_1290), .A2(n_1451), .B1(n_1458), .B2(n_1459), .Y(n_1450) );
OR2x2_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1314), .Y(n_1291) );
AOI31xp33_ASAP7_75t_SL g1292 ( .A1(n_1293), .A2(n_1302), .A3(n_1307), .B(n_1313), .Y(n_1292) );
INVx2_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
AOI22xp5_ASAP7_75t_L g1307 ( .A1(n_1308), .A2(n_1309), .B1(n_1310), .B2(n_1312), .Y(n_1307) );
INVx2_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
NAND3xp33_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1327), .C(n_1335), .Y(n_1314) );
INVx2_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1330), .Y(n_1435) );
INVx2_ASAP7_75t_L g1392 ( .A(n_1336), .Y(n_1392) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1337), .Y(n_1388) );
NAND3xp33_ASAP7_75t_L g1337 ( .A(n_1338), .B(n_1346), .C(n_1363), .Y(n_1337) );
NOR2xp33_ASAP7_75t_L g1338 ( .A(n_1339), .B(n_1343), .Y(n_1338) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
INVx2_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
NOR2xp33_ASAP7_75t_L g1346 ( .A(n_1347), .B(n_1348), .Y(n_1346) );
AOI22xp33_ASAP7_75t_L g1368 ( .A1(n_1356), .A2(n_1360), .B1(n_1369), .B2(n_1371), .Y(n_1368) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
BUFx2_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
OAI22xp5_ASAP7_75t_L g1374 ( .A1(n_1375), .A2(n_1377), .B1(n_1380), .B2(n_1384), .Y(n_1374) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
BUFx2_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1393), .Y(n_1439) );
HB1xp67_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
NOR2x1_ASAP7_75t_L g1395 ( .A(n_1396), .B(n_1416), .Y(n_1395) );
AOI21xp5_ASAP7_75t_L g1396 ( .A1(n_1397), .A2(n_1406), .B(n_1415), .Y(n_1396) );
AOI221xp5_ASAP7_75t_L g1397 ( .A1(n_1398), .A2(n_1399), .B1(n_1400), .B2(n_1402), .C(n_1405), .Y(n_1397) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1404), .Y(n_1403) );
INVx1_ASAP7_75t_L g1728 ( .A(n_1405), .Y(n_1728) );
HB1xp67_ASAP7_75t_L g1409 ( .A(n_1410), .Y(n_1409) );
NAND4xp25_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1420), .C(n_1423), .D(n_1426), .Y(n_1416) );
OAI221xp5_ASAP7_75t_L g1442 ( .A1(n_1443), .A2(n_1691), .B1(n_1693), .B2(n_1734), .C(n_1740), .Y(n_1442) );
AOI211xp5_ASAP7_75t_L g1443 ( .A1(n_1444), .A2(n_1599), .B(n_1641), .C(n_1673), .Y(n_1443) );
NAND5xp2_ASAP7_75t_L g1444 ( .A(n_1445), .B(n_1541), .C(n_1559), .D(n_1588), .E(n_1591), .Y(n_1444) );
AOI321xp33_ASAP7_75t_L g1445 ( .A1(n_1446), .A2(n_1488), .A3(n_1505), .B1(n_1512), .B2(n_1520), .C(n_1531), .Y(n_1445) );
NAND2xp5_ASAP7_75t_L g1446 ( .A(n_1447), .B(n_1484), .Y(n_1446) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1448), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_1449), .B(n_1471), .Y(n_1448) );
CKINVDCx6p67_ASAP7_75t_R g1487 ( .A(n_1449), .Y(n_1487) );
AND2x2_ASAP7_75t_L g1522 ( .A(n_1449), .B(n_1486), .Y(n_1522) );
AND2x2_ASAP7_75t_L g1533 ( .A(n_1449), .B(n_1534), .Y(n_1533) );
OR2x2_ASAP7_75t_L g1550 ( .A(n_1449), .B(n_1486), .Y(n_1550) );
AND2x2_ASAP7_75t_L g1556 ( .A(n_1449), .B(n_1557), .Y(n_1556) );
AND2x2_ASAP7_75t_L g1594 ( .A(n_1449), .B(n_1584), .Y(n_1594) );
OR2x2_ASAP7_75t_L g1598 ( .A(n_1449), .B(n_1535), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1628 ( .A(n_1449), .B(n_1472), .Y(n_1628) );
A2O1A1Ixp33_ASAP7_75t_SL g1677 ( .A1(n_1449), .A2(n_1678), .B(n_1682), .C(n_1684), .Y(n_1677) );
OR2x6_ASAP7_75t_SL g1449 ( .A(n_1450), .B(n_1461), .Y(n_1449) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
AND2x2_ASAP7_75t_L g1452 ( .A(n_1453), .B(n_1455), .Y(n_1452) );
AND2x4_ASAP7_75t_L g1460 ( .A(n_1453), .B(n_1456), .Y(n_1460) );
AND2x4_ASAP7_75t_L g1500 ( .A(n_1453), .B(n_1455), .Y(n_1500) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1454), .Y(n_1466) );
HB1xp67_ASAP7_75t_L g1753 ( .A(n_1455), .Y(n_1753) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
NAND2xp5_ASAP7_75t_L g1465 ( .A(n_1457), .B(n_1466), .Y(n_1465) );
OAI22xp5_ASAP7_75t_L g1497 ( .A1(n_1459), .A2(n_1498), .B1(n_1499), .B2(n_1501), .Y(n_1497) );
INVx1_ASAP7_75t_SL g1459 ( .A(n_1460), .Y(n_1459) );
INVx2_ASAP7_75t_L g1511 ( .A(n_1460), .Y(n_1511) );
OAI22xp5_ASAP7_75t_L g1461 ( .A1(n_1462), .A2(n_1467), .B1(n_1468), .B2(n_1470), .Y(n_1461) );
OAI22xp33_ASAP7_75t_L g1492 ( .A1(n_1462), .A2(n_1493), .B1(n_1494), .B2(n_1495), .Y(n_1492) );
OAI22xp33_ASAP7_75t_L g1515 ( .A1(n_1462), .A2(n_1468), .B1(n_1516), .B2(n_1517), .Y(n_1515) );
BUFx3_ASAP7_75t_L g1574 ( .A(n_1462), .Y(n_1574) );
BUFx6f_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
OAI22xp5_ASAP7_75t_L g1481 ( .A1(n_1463), .A2(n_1468), .B1(n_1482), .B2(n_1483), .Y(n_1481) );
OR2x2_ASAP7_75t_L g1463 ( .A(n_1464), .B(n_1465), .Y(n_1463) );
OR2x2_ASAP7_75t_L g1468 ( .A(n_1464), .B(n_1469), .Y(n_1468) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1464), .Y(n_1476) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1465), .Y(n_1475) );
HB1xp67_ASAP7_75t_L g1755 ( .A(n_1466), .Y(n_1755) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1468), .Y(n_1496) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1469), .Y(n_1478) );
AND2x2_ASAP7_75t_L g1529 ( .A(n_1471), .B(n_1530), .Y(n_1529) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1471), .Y(n_1536) );
OAI32xp33_ASAP7_75t_L g1603 ( .A1(n_1471), .A2(n_1502), .A3(n_1542), .B1(n_1604), .B2(n_1606), .Y(n_1603) );
AND2x2_ASAP7_75t_L g1635 ( .A(n_1471), .B(n_1487), .Y(n_1635) );
NAND2xp5_ASAP7_75t_L g1653 ( .A(n_1471), .B(n_1546), .Y(n_1653) );
AND2x2_ASAP7_75t_L g1471 ( .A(n_1472), .B(n_1480), .Y(n_1471) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1472), .Y(n_1486) );
OR2x2_ASAP7_75t_L g1535 ( .A(n_1472), .B(n_1480), .Y(n_1535) );
AND2x2_ASAP7_75t_L g1557 ( .A(n_1472), .B(n_1558), .Y(n_1557) );
AND2x2_ASAP7_75t_L g1472 ( .A(n_1473), .B(n_1479), .Y(n_1472) );
AND2x4_ASAP7_75t_L g1474 ( .A(n_1475), .B(n_1476), .Y(n_1474) );
AND2x4_ASAP7_75t_L g1477 ( .A(n_1476), .B(n_1478), .Y(n_1477) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1480), .Y(n_1558) );
AND2x2_ASAP7_75t_L g1565 ( .A(n_1480), .B(n_1487), .Y(n_1565) );
AND2x2_ASAP7_75t_L g1584 ( .A(n_1480), .B(n_1486), .Y(n_1584) );
OAI221xp5_ASAP7_75t_L g1560 ( .A1(n_1484), .A2(n_1519), .B1(n_1561), .B2(n_1563), .C(n_1566), .Y(n_1560) );
O2A1O1Ixp33_ASAP7_75t_L g1622 ( .A1(n_1484), .A2(n_1586), .B(n_1623), .C(n_1624), .Y(n_1622) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
A2O1A1Ixp33_ASAP7_75t_L g1637 ( .A1(n_1485), .A2(n_1506), .B(n_1595), .C(n_1638), .Y(n_1637) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_1486), .B(n_1487), .Y(n_1485) );
AND2x2_ASAP7_75t_L g1546 ( .A(n_1487), .B(n_1507), .Y(n_1546) );
AND2x2_ASAP7_75t_L g1583 ( .A(n_1487), .B(n_1584), .Y(n_1583) );
AND2x2_ASAP7_75t_L g1590 ( .A(n_1487), .B(n_1557), .Y(n_1590) );
NOR2xp33_ASAP7_75t_L g1605 ( .A(n_1487), .B(n_1507), .Y(n_1605) );
OR2x2_ASAP7_75t_L g1608 ( .A(n_1487), .B(n_1558), .Y(n_1608) );
AND2x2_ASAP7_75t_L g1616 ( .A(n_1487), .B(n_1529), .Y(n_1616) );
AND2x2_ASAP7_75t_L g1649 ( .A(n_1487), .B(n_1558), .Y(n_1649) );
NAND2xp5_ASAP7_75t_L g1588 ( .A(n_1488), .B(n_1589), .Y(n_1588) );
INVx1_ASAP7_75t_L g1488 ( .A(n_1489), .Y(n_1488) );
OAI22xp5_ASAP7_75t_SL g1646 ( .A1(n_1489), .A2(n_1555), .B1(n_1647), .B2(n_1648), .Y(n_1646) );
OR2x2_ASAP7_75t_L g1489 ( .A(n_1490), .B(n_1502), .Y(n_1489) );
AND2x2_ASAP7_75t_L g1518 ( .A(n_1490), .B(n_1519), .Y(n_1518) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1490), .Y(n_1525) );
INVx3_ASAP7_75t_L g1587 ( .A(n_1490), .Y(n_1587) );
AND2x2_ASAP7_75t_L g1595 ( .A(n_1490), .B(n_1582), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1633 ( .A(n_1490), .B(n_1552), .Y(n_1633) );
AOI221xp5_ASAP7_75t_L g1650 ( .A1(n_1490), .A2(n_1651), .B1(n_1652), .B2(n_1654), .C(n_1658), .Y(n_1650) );
AND2x2_ASAP7_75t_L g1675 ( .A(n_1490), .B(n_1502), .Y(n_1675) );
AND2x2_ASAP7_75t_L g1684 ( .A(n_1490), .B(n_1540), .Y(n_1684) );
INVx3_ASAP7_75t_L g1490 ( .A(n_1491), .Y(n_1490) );
OR2x2_ASAP7_75t_L g1597 ( .A(n_1491), .B(n_1527), .Y(n_1597) );
AND2x2_ASAP7_75t_L g1661 ( .A(n_1491), .B(n_1502), .Y(n_1661) );
OR2x2_ASAP7_75t_L g1491 ( .A(n_1492), .B(n_1497), .Y(n_1491) );
HB1xp67_ASAP7_75t_L g1576 ( .A(n_1495), .Y(n_1576) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1500), .Y(n_1570) );
INVx2_ASAP7_75t_L g1519 ( .A(n_1502), .Y(n_1519) );
OR2x2_ASAP7_75t_L g1527 ( .A(n_1502), .B(n_1514), .Y(n_1527) );
AND2x2_ASAP7_75t_L g1540 ( .A(n_1502), .B(n_1514), .Y(n_1540) );
NAND2xp5_ASAP7_75t_L g1548 ( .A(n_1502), .B(n_1549), .Y(n_1548) );
OR2x2_ASAP7_75t_L g1554 ( .A(n_1502), .B(n_1552), .Y(n_1554) );
AND2x2_ASAP7_75t_L g1562 ( .A(n_1502), .B(n_1552), .Y(n_1562) );
AND2x4_ASAP7_75t_L g1502 ( .A(n_1503), .B(n_1504), .Y(n_1502) );
NOR2x1_ASAP7_75t_L g1607 ( .A(n_1505), .B(n_1608), .Y(n_1607) );
NAND2xp5_ASAP7_75t_L g1610 ( .A(n_1505), .B(n_1522), .Y(n_1610) );
AND2x2_ASAP7_75t_L g1613 ( .A(n_1505), .B(n_1594), .Y(n_1613) );
OR2x2_ASAP7_75t_L g1624 ( .A(n_1505), .B(n_1554), .Y(n_1624) );
NAND2xp5_ASAP7_75t_L g1647 ( .A(n_1505), .B(n_1612), .Y(n_1647) );
INVx2_ASAP7_75t_L g1505 ( .A(n_1506), .Y(n_1505) );
AND2x2_ASAP7_75t_L g1564 ( .A(n_1506), .B(n_1565), .Y(n_1564) );
NAND2xp5_ASAP7_75t_L g1580 ( .A(n_1506), .B(n_1581), .Y(n_1580) );
NAND2xp5_ASAP7_75t_L g1593 ( .A(n_1506), .B(n_1594), .Y(n_1593) );
AND2x2_ASAP7_75t_L g1686 ( .A(n_1506), .B(n_1687), .Y(n_1686) );
INVx2_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
INVx4_ASAP7_75t_L g1530 ( .A(n_1507), .Y(n_1530) );
NAND2xp5_ASAP7_75t_L g1551 ( .A(n_1507), .B(n_1552), .Y(n_1551) );
OR2x2_ASAP7_75t_L g1602 ( .A(n_1507), .B(n_1535), .Y(n_1602) );
NAND2xp5_ASAP7_75t_L g1623 ( .A(n_1507), .B(n_1582), .Y(n_1623) );
OR2x2_ASAP7_75t_L g1669 ( .A(n_1507), .B(n_1581), .Y(n_1669) );
NAND2xp5_ASAP7_75t_L g1676 ( .A(n_1507), .B(n_1556), .Y(n_1676) );
OR2x2_ASAP7_75t_L g1683 ( .A(n_1507), .B(n_1598), .Y(n_1683) );
AND2x6_ASAP7_75t_L g1507 ( .A(n_1508), .B(n_1509), .Y(n_1507) );
INVx2_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
OAI22xp5_ASAP7_75t_L g1568 ( .A1(n_1511), .A2(n_1569), .B1(n_1570), .B2(n_1571), .Y(n_1568) );
INVx1_ASAP7_75t_L g1692 ( .A(n_1511), .Y(n_1692) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1512), .Y(n_1651) );
NAND2xp5_ASAP7_75t_L g1512 ( .A(n_1513), .B(n_1518), .Y(n_1512) );
INVx1_ASAP7_75t_L g1645 ( .A(n_1513), .Y(n_1645) );
NAND2xp5_ASAP7_75t_L g1648 ( .A(n_1513), .B(n_1649), .Y(n_1648) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1513), .Y(n_1655) );
INVx1_ASAP7_75t_L g1672 ( .A(n_1513), .Y(n_1672) );
HB1xp67_ASAP7_75t_L g1513 ( .A(n_1514), .Y(n_1513) );
INVx2_ASAP7_75t_SL g1552 ( .A(n_1514), .Y(n_1552) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1519), .Y(n_1543) );
OAI22xp5_ASAP7_75t_L g1520 ( .A1(n_1521), .A2(n_1523), .B1(n_1525), .B2(n_1528), .Y(n_1520) );
INVxp67_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
AND2x2_ASAP7_75t_L g1620 ( .A(n_1522), .B(n_1530), .Y(n_1620) );
INVxp67_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
AND2x2_ASAP7_75t_L g1524 ( .A(n_1525), .B(n_1526), .Y(n_1524) );
AOI21xp5_ASAP7_75t_L g1636 ( .A1(n_1525), .A2(n_1544), .B(n_1566), .Y(n_1636) );
AOI22xp5_ASAP7_75t_L g1662 ( .A1(n_1525), .A2(n_1663), .B1(n_1666), .B2(n_1670), .Y(n_1662) );
OAI211xp5_ASAP7_75t_L g1599 ( .A1(n_1526), .A2(n_1600), .B(n_1611), .C(n_1625), .Y(n_1599) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
INVxp67_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1530), .Y(n_1539) );
NAND2xp5_ASAP7_75t_L g1561 ( .A(n_1530), .B(n_1562), .Y(n_1561) );
AND2x2_ASAP7_75t_L g1589 ( .A(n_1530), .B(n_1590), .Y(n_1589) );
AOI21xp5_ASAP7_75t_L g1531 ( .A1(n_1532), .A2(n_1536), .B(n_1537), .Y(n_1531) );
AND2x2_ASAP7_75t_L g1664 ( .A(n_1532), .B(n_1665), .Y(n_1664) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
OAI31xp33_ASAP7_75t_L g1685 ( .A1(n_1533), .A2(n_1564), .A3(n_1686), .B(n_1688), .Y(n_1685) );
NAND2xp5_ASAP7_75t_L g1545 ( .A(n_1534), .B(n_1546), .Y(n_1545) );
NAND2xp5_ASAP7_75t_L g1657 ( .A(n_1534), .B(n_1605), .Y(n_1657) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
INVx1_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
AND2x2_ASAP7_75t_L g1538 ( .A(n_1539), .B(n_1540), .Y(n_1538) );
NAND2xp5_ASAP7_75t_L g1627 ( .A(n_1539), .B(n_1628), .Y(n_1627) );
AND2x2_ASAP7_75t_L g1638 ( .A(n_1539), .B(n_1557), .Y(n_1638) );
INVx1_ASAP7_75t_L g1640 ( .A(n_1540), .Y(n_1640) );
AOI211xp5_ASAP7_75t_SL g1541 ( .A1(n_1542), .A2(n_1544), .B(n_1547), .C(n_1553), .Y(n_1541) );
OAI22xp5_ASAP7_75t_L g1626 ( .A1(n_1542), .A2(n_1627), .B1(n_1629), .B2(n_1630), .Y(n_1626) );
AOI21xp5_ASAP7_75t_L g1642 ( .A1(n_1542), .A2(n_1643), .B(n_1646), .Y(n_1642) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1543), .Y(n_1542) );
NAND2xp5_ASAP7_75t_L g1644 ( .A(n_1544), .B(n_1645), .Y(n_1644) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
OR2x2_ASAP7_75t_L g1671 ( .A(n_1545), .B(n_1672), .Y(n_1671) );
INVxp67_ASAP7_75t_SL g1547 ( .A(n_1548), .Y(n_1547) );
INVxp33_ASAP7_75t_L g1659 ( .A(n_1549), .Y(n_1659) );
NOR2xp33_ASAP7_75t_L g1549 ( .A(n_1550), .B(n_1551), .Y(n_1549) );
INVx1_ASAP7_75t_L g1687 ( .A(n_1550), .Y(n_1687) );
INVx2_ASAP7_75t_SL g1582 ( .A(n_1552), .Y(n_1582) );
NOR2xp33_ASAP7_75t_L g1553 ( .A(n_1554), .B(n_1555), .Y(n_1553) );
INVx2_ASAP7_75t_L g1612 ( .A(n_1554), .Y(n_1612) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1556), .Y(n_1555) );
OAI21xp33_ASAP7_75t_SL g1619 ( .A1(n_1556), .A2(n_1620), .B(n_1621), .Y(n_1619) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1557), .Y(n_1680) );
OAI21xp5_ASAP7_75t_L g1559 ( .A1(n_1560), .A2(n_1577), .B(n_1585), .Y(n_1559) );
INVx1_ASAP7_75t_L g1629 ( .A(n_1562), .Y(n_1629) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
INVxp67_ASAP7_75t_L g1630 ( .A(n_1565), .Y(n_1630) );
NAND2xp5_ASAP7_75t_L g1585 ( .A(n_1566), .B(n_1586), .Y(n_1585) );
CKINVDCx5p33_ASAP7_75t_R g1566 ( .A(n_1567), .Y(n_1566) );
OR2x6_ASAP7_75t_SL g1567 ( .A(n_1568), .B(n_1572), .Y(n_1567) );
OAI22xp5_ASAP7_75t_L g1572 ( .A1(n_1573), .A2(n_1574), .B1(n_1575), .B2(n_1576), .Y(n_1572) );
INVxp67_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
NAND2xp5_ASAP7_75t_L g1578 ( .A(n_1579), .B(n_1583), .Y(n_1578) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
AOI221xp5_ASAP7_75t_L g1600 ( .A1(n_1582), .A2(n_1587), .B1(n_1601), .B2(n_1603), .C(n_1609), .Y(n_1600) );
NOR2xp33_ASAP7_75t_L g1609 ( .A(n_1582), .B(n_1610), .Y(n_1609) );
NAND2xp5_ASAP7_75t_L g1618 ( .A(n_1582), .B(n_1602), .Y(n_1618) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1582), .Y(n_1690) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1584), .Y(n_1681) );
AOI211xp5_ASAP7_75t_L g1625 ( .A1(n_1586), .A2(n_1626), .B(n_1631), .C(n_1639), .Y(n_1625) );
NOR2xp33_ASAP7_75t_L g1668 ( .A(n_1586), .B(n_1669), .Y(n_1668) );
INVx1_ASAP7_75t_SL g1586 ( .A(n_1587), .Y(n_1586) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1590), .Y(n_1665) );
AOI21xp5_ASAP7_75t_L g1591 ( .A1(n_1592), .A2(n_1595), .B(n_1596), .Y(n_1591) );
INVx1_ASAP7_75t_L g1592 ( .A(n_1593), .Y(n_1592) );
NOR2xp33_ASAP7_75t_L g1596 ( .A(n_1597), .B(n_1598), .Y(n_1596) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1597), .Y(n_1621) );
NOR2xp33_ASAP7_75t_L g1639 ( .A(n_1598), .B(n_1640), .Y(n_1639) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1602), .Y(n_1601) );
INVx1_ASAP7_75t_L g1604 ( .A(n_1605), .Y(n_1604) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1607), .Y(n_1606) );
AOI211xp5_ASAP7_75t_L g1611 ( .A1(n_1612), .A2(n_1613), .B(n_1614), .C(n_1622), .Y(n_1611) );
OAI21xp33_ASAP7_75t_L g1614 ( .A1(n_1615), .A2(n_1617), .B(n_1619), .Y(n_1614) );
INVx1_ASAP7_75t_L g1615 ( .A(n_1616), .Y(n_1615) );
INVxp67_ASAP7_75t_SL g1617 ( .A(n_1618), .Y(n_1617) );
NAND2xp5_ASAP7_75t_L g1666 ( .A(n_1624), .B(n_1667), .Y(n_1666) );
OAI211xp5_ASAP7_75t_L g1631 ( .A1(n_1632), .A2(n_1634), .B(n_1636), .C(n_1637), .Y(n_1631) );
INVx1_ASAP7_75t_L g1632 ( .A(n_1633), .Y(n_1632) );
AOI21xp33_ASAP7_75t_SL g1658 ( .A1(n_1634), .A2(n_1659), .B(n_1660), .Y(n_1658) );
INVx1_ASAP7_75t_L g1634 ( .A(n_1635), .Y(n_1634) );
NAND3xp33_ASAP7_75t_L g1641 ( .A(n_1642), .B(n_1650), .C(n_1662), .Y(n_1641) );
INVxp67_ASAP7_75t_SL g1643 ( .A(n_1644), .Y(n_1643) );
INVx1_ASAP7_75t_L g1652 ( .A(n_1653), .Y(n_1652) );
AND2x2_ASAP7_75t_L g1654 ( .A(n_1655), .B(n_1656), .Y(n_1654) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1657), .Y(n_1656) );
INVx1_ASAP7_75t_L g1660 ( .A(n_1661), .Y(n_1660) );
INVxp67_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
INVxp67_ASAP7_75t_SL g1667 ( .A(n_1668), .Y(n_1667) );
INVx1_ASAP7_75t_L g1670 ( .A(n_1671), .Y(n_1670) );
OAI211xp5_ASAP7_75t_L g1673 ( .A1(n_1674), .A2(n_1676), .B(n_1677), .C(n_1685), .Y(n_1673) );
INVx1_ASAP7_75t_L g1674 ( .A(n_1675), .Y(n_1674) );
NAND2xp5_ASAP7_75t_L g1689 ( .A(n_1675), .B(n_1690), .Y(n_1689) );
INVx1_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_1680), .B(n_1681), .Y(n_1679) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1683), .Y(n_1682) );
INVx1_ASAP7_75t_L g1688 ( .A(n_1689), .Y(n_1688) );
INVx1_ASAP7_75t_L g1691 ( .A(n_1692), .Y(n_1691) );
INVx1_ASAP7_75t_L g1693 ( .A(n_1694), .Y(n_1693) );
HB1xp67_ASAP7_75t_L g1748 ( .A(n_1695), .Y(n_1748) );
NAND3xp33_ASAP7_75t_L g1695 ( .A(n_1696), .B(n_1709), .C(n_1716), .Y(n_1695) );
AND3x1_ASAP7_75t_L g1696 ( .A(n_1697), .B(n_1700), .C(n_1707), .Y(n_1696) );
AND2x2_ASAP7_75t_L g1709 ( .A(n_1710), .B(n_1713), .Y(n_1709) );
OAI211xp5_ASAP7_75t_L g1724 ( .A1(n_1712), .A2(n_1725), .B(n_1726), .C(n_1727), .Y(n_1724) );
NAND3xp33_ASAP7_75t_L g1718 ( .A(n_1719), .B(n_1724), .C(n_1728), .Y(n_1718) );
OAI211xp5_ASAP7_75t_L g1719 ( .A1(n_1720), .A2(n_1721), .B(n_1722), .C(n_1723), .Y(n_1719) );
CKINVDCx14_ASAP7_75t_R g1734 ( .A(n_1735), .Y(n_1734) );
INVx4_ASAP7_75t_L g1735 ( .A(n_1736), .Y(n_1735) );
INVx1_ASAP7_75t_L g1736 ( .A(n_1737), .Y(n_1736) );
INVx1_ASAP7_75t_L g1737 ( .A(n_1738), .Y(n_1737) );
INVx1_ASAP7_75t_L g1738 ( .A(n_1739), .Y(n_1738) );
HB1xp67_ASAP7_75t_SL g1741 ( .A(n_1742), .Y(n_1741) );
A2O1A1Ixp33_ASAP7_75t_L g1751 ( .A1(n_1743), .A2(n_1752), .B(n_1754), .C(n_1756), .Y(n_1751) );
INVxp33_ASAP7_75t_SL g1744 ( .A(n_1745), .Y(n_1744) );
INVx1_ASAP7_75t_L g1747 ( .A(n_1748), .Y(n_1747) );
BUFx2_ASAP7_75t_L g1749 ( .A(n_1750), .Y(n_1749) );
HB1xp67_ASAP7_75t_L g1750 ( .A(n_1751), .Y(n_1750) );
INVx1_ASAP7_75t_L g1752 ( .A(n_1753), .Y(n_1752) );
INVx1_ASAP7_75t_L g1754 ( .A(n_1755), .Y(n_1754) );
endmodule