module fake_jpeg_20396_n_214 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_214);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_214;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_SL g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_31),
.Y(n_55)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_31),
.Y(n_47)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_25),
.B1(n_30),
.B2(n_29),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_44),
.A2(n_33),
.B1(n_26),
.B2(n_23),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_56),
.Y(n_73)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

NAND3xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_28),
.C(n_14),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_21),
.B(n_18),
.C(n_17),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_22),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_22),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_25),
.B1(n_30),
.B2(n_27),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_64),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_16),
.Y(n_59)
);

OR2x2_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_33),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_38),
.Y(n_74)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_22),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_36),
.A2(n_27),
.B1(n_21),
.B2(n_18),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_18),
.B1(n_26),
.B2(n_23),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_68),
.B(n_79),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_37),
.B1(n_33),
.B2(n_38),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_69),
.A2(n_62),
.B1(n_49),
.B2(n_58),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_43),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_76),
.Y(n_115)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_71),
.A2(n_77),
.B(n_6),
.C(n_7),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_78),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_43),
.Y(n_76)
);

AO22x1_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_33),
.B1(n_18),
.B2(n_23),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_63),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_81),
.Y(n_120)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_17),
.B(n_33),
.C(n_3),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_84),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_118)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_1),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_46),
.B(n_1),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_61),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_9),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_20),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_95),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_49),
.A2(n_26),
.B1(n_20),
.B2(n_16),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_16),
.B1(n_2),
.B2(n_4),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_54),
.B(n_20),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_54),
.Y(n_96)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_50),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_105),
.Y(n_132)
);

MAJx2_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_46),
.C(n_62),
.Y(n_103)
);

XNOR2x1_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_69),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_58),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_111),
.B1(n_117),
.B2(n_116),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_5),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_122),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_85),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_SL g126 ( 
.A(n_118),
.B(n_79),
.C(n_68),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_88),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_86),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_93),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_84),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_137),
.C(n_123),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_127),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_126),
.B(n_130),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_72),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_128),
.B(n_134),
.Y(n_156)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_135),
.A2(n_138),
.B1(n_111),
.B2(n_117),
.Y(n_152)
);

AO22x1_ASAP7_75t_SL g136 ( 
.A1(n_103),
.A2(n_69),
.B1(n_77),
.B2(n_93),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_140),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_68),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_99),
.A2(n_69),
.B1(n_83),
.B2(n_77),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_88),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_139),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_141),
.A2(n_142),
.B(n_96),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_99),
.A2(n_104),
.B(n_118),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_101),
.B(n_67),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_143),
.B(n_145),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_110),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_109),
.B(n_112),
.C(n_106),
.D(n_115),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_146),
.A2(n_147),
.B(n_159),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_115),
.B(n_106),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_152),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_108),
.B1(n_120),
.B2(n_122),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_153),
.A2(n_157),
.B1(n_158),
.B2(n_138),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_113),
.Y(n_155)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_112),
.B1(n_115),
.B2(n_119),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_119),
.B1(n_97),
.B2(n_121),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_67),
.C(n_121),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_161),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_144),
.Y(n_162)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_154),
.B(n_133),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_164),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_159),
.A2(n_126),
.B(n_131),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_172),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_140),
.C(n_133),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_173),
.B(n_148),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_171),
.Y(n_185)
);

OAI322xp33_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_124),
.A3(n_131),
.B1(n_141),
.B2(n_136),
.C1(n_132),
.C2(n_135),
.Y(n_172)
);

AO21x1_ASAP7_75t_L g173 ( 
.A1(n_151),
.A2(n_136),
.B(n_102),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

OAI322xp33_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_114),
.C2(n_134),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_179),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_149),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_151),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_183),
.Y(n_195)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_153),
.B1(n_158),
.B2(n_157),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_184),
.A2(n_167),
.B1(n_168),
.B2(n_165),
.Y(n_193)
);

NOR3xp33_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_147),
.C(n_146),
.Y(n_190)
);

AO21x1_ASAP7_75t_L g188 ( 
.A1(n_181),
.A2(n_173),
.B(n_169),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_190),
.A2(n_192),
.B1(n_193),
.B2(n_196),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_177),
.A2(n_164),
.B(n_169),
.Y(n_191)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_168),
.B(n_160),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_185),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_195),
.A2(n_152),
.B1(n_185),
.B2(n_186),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_200),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_179),
.C(n_180),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_196),
.A2(n_155),
.B1(n_162),
.B2(n_178),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_10),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_189),
.C(n_190),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_206),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_201),
.A2(n_197),
.B(n_188),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

A2O1A1O1Ixp25_ASAP7_75t_L g207 ( 
.A1(n_205),
.A2(n_202),
.B(n_199),
.C(n_198),
.D(n_12),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_10),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_211),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_209),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_212),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_211),
.Y(n_214)
);


endmodule