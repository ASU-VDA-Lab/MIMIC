module fake_jpeg_31384_n_211 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_211);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_211;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_118;
wire n_128;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_13),
.B(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_18),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_17),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_40),
.A2(n_50),
.B1(n_51),
.B2(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_1),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_2),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_48),
.Y(n_58)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_6),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_6),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_22),
.A2(n_15),
.B1(n_11),
.B2(n_12),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_23),
.B(n_10),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_54),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_22),
.B(n_10),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_24),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_27),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_24),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_62),
.B(n_59),
.Y(n_99)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_65),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_27),
.B1(n_36),
.B2(n_16),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_69),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_74),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_32),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_73),
.B(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_30),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_76),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_30),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_41),
.B(n_23),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_79),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_34),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_37),
.B(n_34),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_88),
.Y(n_115)
);

BUFx8_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_86),
.Y(n_89)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_32),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_40),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_98),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_86),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_94),
.B(n_95),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_86),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_100),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_67),
.A2(n_47),
.B1(n_44),
.B2(n_54),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_60),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_19),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_102),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_20),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_20),
.C(n_25),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_25),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_59),
.Y(n_128)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_58),
.B(n_36),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_128),
.B(n_136),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_80),
.C(n_72),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_130),
.B(n_93),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_131),
.Y(n_157)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_116),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_95),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_134),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_97),
.B1(n_113),
.B2(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_84),
.B(n_65),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_69),
.Y(n_149)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_124),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_140),
.B(n_144),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_142),
.B(n_104),
.Y(n_169)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_106),
.B(n_129),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g146 ( 
.A(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_153),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_100),
.B1(n_99),
.B2(n_112),
.Y(n_147)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_149),
.A2(n_68),
.B(n_122),
.Y(n_166)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_131),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_96),
.B1(n_111),
.B2(n_115),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_123),
.B1(n_130),
.B2(n_137),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_135),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_138),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_152),
.B(n_108),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_160),
.Y(n_176)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_119),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_168),
.C(n_141),
.Y(n_175)
);

A2O1A1O1Ixp25_ASAP7_75t_L g165 ( 
.A1(n_149),
.A2(n_122),
.B(n_119),
.C(n_110),
.D(n_98),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_169),
.Y(n_177)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_90),
.C(n_129),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_151),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_127),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_172),
.A2(n_156),
.B1(n_163),
.B2(n_167),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_150),
.C(n_154),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_179),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_178),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_145),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_141),
.C(n_157),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_158),
.A2(n_156),
.B(n_73),
.Y(n_180)
);

AO21x1_ASAP7_75t_L g187 ( 
.A1(n_180),
.A2(n_161),
.B(n_171),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_181),
.A2(n_139),
.B1(n_127),
.B2(n_125),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_126),
.C(n_125),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_182),
.Y(n_186)
);

AOI322xp5_ASAP7_75t_L g185 ( 
.A1(n_183),
.A2(n_166),
.A3(n_164),
.B1(n_171),
.B2(n_165),
.C1(n_172),
.C2(n_170),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_176),
.C(n_182),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_188),
.Y(n_193)
);

O2A1O1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_173),
.A2(n_121),
.B(n_143),
.C(n_126),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_139),
.B(n_89),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_184),
.B(n_175),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_191),
.B(n_143),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_194),
.B(n_198),
.Y(n_199)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_186),
.C(n_192),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_189),
.B1(n_186),
.B2(n_191),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_94),
.Y(n_198)
);

AOI322xp5_ASAP7_75t_L g205 ( 
.A1(n_200),
.A2(n_202),
.A3(n_197),
.B1(n_105),
.B2(n_89),
.C1(n_69),
.C2(n_61),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_190),
.C(n_177),
.Y(n_204)
);

OAI31xp33_ASAP7_75t_L g202 ( 
.A1(n_193),
.A2(n_177),
.A3(n_190),
.B(n_134),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_204),
.A2(n_205),
.B(n_206),
.Y(n_208)
);

AOI322xp5_ASAP7_75t_L g206 ( 
.A1(n_203),
.A2(n_87),
.A3(n_61),
.B1(n_16),
.B2(n_26),
.C1(n_114),
.C2(n_82),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_199),
.A2(n_26),
.A3(n_60),
.B1(n_71),
.B2(n_82),
.C1(n_202),
.C2(n_201),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_207),
.A2(n_71),
.B(n_26),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_209),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_208),
.C(n_26),
.Y(n_211)
);


endmodule