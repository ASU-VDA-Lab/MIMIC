module fake_jpeg_21602_n_154 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_154);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_28),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_32),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_59),
.B(n_21),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_64),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_81),
.Y(n_85)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

NOR2xp67_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_67),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_84),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_81),
.A2(n_74),
.B1(n_55),
.B2(n_66),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_87),
.A2(n_50),
.B1(n_52),
.B2(n_71),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_48),
.B1(n_63),
.B2(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_52),
.Y(n_96)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_85),
.B(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_94),
.B(n_96),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_53),
.B1(n_70),
.B2(n_65),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_56),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_98),
.B(n_54),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_101),
.B(n_60),
.Y(n_112)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_91),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_104),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_108),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_105),
.A2(n_83),
.B1(n_84),
.B2(n_92),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_115),
.B1(n_117),
.B2(n_102),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_95),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_97),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_111),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_112),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_83),
.B1(n_62),
.B2(n_71),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_119),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_73),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_124),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_69),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_72),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_120),
.C(n_113),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_61),
.B1(n_1),
.B2(n_2),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_5),
.C(n_6),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_126),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_134),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_125),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_138),
.Y(n_141)
);

NAND3xp33_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_31),
.C(n_40),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_136),
.A2(n_137),
.B(n_139),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_131),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_140),
.A2(n_132),
.B1(n_131),
.B2(n_128),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_141),
.Y(n_145)
);

AOI322xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_142),
.A3(n_136),
.B1(n_121),
.B2(n_113),
.C1(n_17),
.C2(n_19),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_121),
.C(n_37),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_147),
.A2(n_36),
.B1(n_47),
.B2(n_45),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_24),
.B(n_44),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_23),
.B(n_41),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_16),
.C(n_26),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_38),
.B(n_9),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_120),
.B1(n_9),
.B2(n_10),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_7),
.Y(n_154)
);


endmodule