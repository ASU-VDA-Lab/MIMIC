module real_jpeg_31905_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_0),
.Y(n_169)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_0),
.Y(n_294)
);

NAND2xp33_ASAP7_75t_SL g285 ( 
.A(n_1),
.B(n_96),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_1),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_1),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_2),
.B(n_182),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_2),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_2),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_2),
.B(n_374),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

AND2x4_ASAP7_75t_L g200 ( 
.A(n_4),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_4),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_4),
.B(n_312),
.Y(n_311)
);

NAND2xp33_ASAP7_75t_SL g322 ( 
.A(n_4),
.B(n_323),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_4),
.B(n_346),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_5),
.Y(n_96)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_6),
.Y(n_81)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_7),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_7),
.Y(n_186)
);

AND2x4_ASAP7_75t_L g40 ( 
.A(n_8),
.B(n_41),
.Y(n_40)
);

NAND2xp33_ASAP7_75t_SL g44 ( 
.A(n_8),
.B(n_45),
.Y(n_44)
);

AND2x4_ASAP7_75t_L g57 ( 
.A(n_8),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_8),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_8),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_8),
.B(n_63),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_8),
.B(n_185),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_8),
.B(n_169),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_9),
.B(n_182),
.Y(n_181)
);

AND2x2_ASAP7_75t_SL g230 ( 
.A(n_9),
.B(n_231),
.Y(n_230)
);

NAND2xp33_ASAP7_75t_SL g287 ( 
.A(n_9),
.B(n_288),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_9),
.B(n_348),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_9),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_10),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_10),
.B(n_50),
.Y(n_49)
);

NAND2x1_ASAP7_75t_SL g92 ( 
.A(n_10),
.B(n_93),
.Y(n_92)
);

NAND2xp67_ASAP7_75t_SL g135 ( 
.A(n_10),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_10),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_10),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_10),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_10),
.B(n_292),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_19),
.B(n_20),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_12),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_13),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_14),
.B(n_51),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_14),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_14),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_14),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_14),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_14),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_14),
.B(n_327),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_14),
.Y(n_342)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_15),
.Y(n_245)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_15),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_16),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_16),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_24),
.Y(n_23)
);

AND2x4_ASAP7_75t_SL g62 ( 
.A(n_17),
.B(n_63),
.Y(n_62)
);

NAND2x1p5_ASAP7_75t_L g65 ( 
.A(n_17),
.B(n_66),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g77 ( 
.A(n_17),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_17),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_17),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_17),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_17),
.B(n_169),
.Y(n_168)
);

AO31x2_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_28),
.A3(n_268),
.B(n_417),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_22),
.B(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_26),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_23),
.B(n_57),
.C(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_23),
.A2(n_56),
.B1(n_57),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_23),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1O1Ixp25_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_170),
.B(n_254),
.C(n_255),
.D(n_266),
.Y(n_28)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_29),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_110),
.Y(n_29)
);

NOR2x1_ASAP7_75t_L g254 ( 
.A(n_30),
.B(n_110),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_84),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_31),
.B(n_86),
.C(n_88),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_61),
.C(n_69),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_32),
.A2(n_33),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_47),
.Y(n_33)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_40),
.C(n_44),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_35),
.A2(n_36),
.B1(n_40),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_40),
.Y(n_160)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_40),
.B(n_198),
.C(n_200),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_40),
.A2(n_160),
.B1(n_200),
.B2(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_42),
.Y(n_313)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_42),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_43),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_44),
.B(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_44),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_44),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_56),
.B2(n_57),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_57),
.C(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_51),
.B(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_55),
.Y(n_201)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_55),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_56),
.B(n_197),
.C(n_202),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_56),
.A2(n_57),
.B1(n_202),
.B2(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_61),
.B(n_69),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.C(n_68),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_62),
.A2(n_65),
.B1(n_82),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_62),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_62),
.B(n_119),
.C(n_124),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_62),
.B(n_120),
.Y(n_144)
);

MAJx2_ASAP7_75t_L g344 ( 
.A(n_62),
.B(n_345),
.C(n_347),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_62),
.A2(n_117),
.B1(n_347),
.B2(n_363),
.Y(n_362)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_65),
.A2(n_77),
.B1(n_82),
.B2(n_83),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_65),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_70),
.C(n_77),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_65),
.B(n_150),
.C(n_284),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_67),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_67),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_67),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_68),
.B(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_76),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_77),
.A2(n_83),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_77),
.B(n_230),
.Y(n_333)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_82),
.B(n_283),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_83),
.B(n_157),
.C(n_229),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_83),
.B(n_104),
.C(n_261),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_100),
.B2(n_101),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_92),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_96),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_96),
.Y(n_203)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_97),
.B(n_98),
.C(n_100),
.Y(n_265)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_129),
.C(n_133),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_156),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g237 ( 
.A(n_106),
.B(n_238),
.C(n_243),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_L g260 ( 
.A1(n_106),
.A2(n_164),
.B1(n_190),
.B2(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_106),
.Y(n_261)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_107),
.B(n_243),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_109),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_114),
.C(n_139),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_111),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_114),
.B(n_140),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_128),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_115),
.B(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_118),
.B(n_128),
.Y(n_206)
);

INVxp33_ASAP7_75t_SL g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_125),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_164),
.C(n_168),
.Y(n_163)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_125),
.B(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_126),
.Y(n_310)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_134),
.B1(n_135),
.B2(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_129),
.A2(n_157),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_130),
.Y(n_346)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_158),
.C(n_161),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_142),
.B(n_209),
.Y(n_208)
);

MAJx2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.C(n_155),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_143),
.Y(n_219)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_146),
.B(n_155),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_152),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_152),
.Y(n_178)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_150),
.A2(n_151),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_161),
.Y(n_209)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_164),
.Y(n_190)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_184),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_189),
.Y(n_188)
);

XNOR2x1_ASAP7_75t_L g224 ( 
.A(n_168),
.B(n_225),
.Y(n_224)
);

INVx4_ASAP7_75t_SL g343 ( 
.A(n_169),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_212),
.B(n_253),
.Y(n_170)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_171),
.Y(n_271)
);

NOR2x1_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_210),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_172),
.B(n_210),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_204),
.C(n_207),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_173),
.B(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_191),
.C(n_195),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2x1_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.C(n_188),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_177),
.B(n_179),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_183),
.B(n_187),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_180),
.A2(n_181),
.B1(n_184),
.B2(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_184),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_R g340 ( 
.A(n_184),
.B(n_341),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_184),
.A2(n_226),
.B1(n_341),
.B2(n_378),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_187),
.B(n_298),
.C(n_300),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_188),
.B(n_407),
.Y(n_406)
);

NOR3xp33_ASAP7_75t_L g418 ( 
.A(n_190),
.B(n_261),
.C(n_262),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_191),
.A2(n_192),
.B1(n_195),
.B2(n_196),
.Y(n_216)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_197),
.B(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_234),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_200),
.Y(n_235)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_201),
.Y(n_308)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_205),
.B(n_208),
.Y(n_252)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_251),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_213),
.B(n_251),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.C(n_221),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_215),
.B(n_218),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2x1_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_221),
.B(n_415),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_236),
.C(n_246),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_222),
.B(n_405),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_227),
.C(n_233),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_224),
.B(n_228),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_233),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_236),
.A2(n_237),
.B1(n_247),
.B2(n_248),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_237),
.Y(n_236)
);

XOR2x2_ASAP7_75t_L g391 ( 
.A(n_238),
.B(n_392),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.C(n_242),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_239),
.B(n_241),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_242),
.B(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_255),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_257),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_265),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_264),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_260),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_264),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_275),
.Y(n_268)
);

NOR3xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_273),
.C(n_274),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

INVxp33_ASAP7_75t_SL g275 ( 
.A(n_276),
.Y(n_275)
);

A2O1A1O1Ixp25_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_396),
.B(n_410),
.C(n_411),
.D(n_416),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_379),
.C(n_394),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_351),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_318),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_302),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_281),
.B(n_318),
.C(n_395),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_286),
.C(n_296),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_282),
.B(n_286),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_285),
.Y(n_284)
);

OA21x2_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_291),
.B(n_295),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_291),
.Y(n_295)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx8_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_295),
.A2(n_304),
.B1(n_314),
.B2(n_315),
.Y(n_303)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_297),
.B(n_354),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_302),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_316),
.Y(n_302)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_309),
.C(n_311),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_305),
.A2(n_306),
.B1(n_309),
.B2(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_305),
.B(n_309),
.C(n_311),
.Y(n_388)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_309),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_311),
.B(n_337),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

MAJx2_ASAP7_75t_L g387 ( 
.A(n_314),
.B(n_316),
.C(n_388),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_335),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_332),
.Y(n_319)
);

MAJx2_ASAP7_75t_L g393 ( 
.A(n_320),
.B(n_332),
.C(n_335),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_331),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_325),
.B1(n_326),
.B2(n_330),
.Y(n_321)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_322),
.Y(n_330)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_324),
.Y(n_369)
);

MAJx2_ASAP7_75t_L g390 ( 
.A(n_325),
.B(n_330),
.C(n_331),
.Y(n_390)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_339),
.C(n_344),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_336),
.B(n_357),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_339),
.A2(n_340),
.B1(n_344),
.B2(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_341),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_344),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_345),
.B(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_347),
.Y(n_363)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_355),
.C(n_359),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_364),
.C(n_376),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_370),
.C(n_372),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

XOR2x2_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_393),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_382),
.B1(n_385),
.B2(n_386),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_398),
.C(n_399),
.Y(n_397)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

XNOR2x1_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_386),
.Y(n_399)
);

XNOR2x1_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_389),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_387),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_390),
.B(n_391),
.C(n_402),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_393),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_400),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_400),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_403),
.Y(n_400)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_401),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_406),
.B1(n_408),
.B2(n_409),
.Y(n_403)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_404),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_404),
.B(n_406),
.C(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_406),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_414),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_412),
.B(n_414),
.Y(n_416)
);


endmodule