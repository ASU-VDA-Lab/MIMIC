module fake_jpeg_22057_n_198 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_198);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx4_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_12),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_10),
.B(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_48),
.Y(n_52)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_38),
.B(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_2),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_46),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_34),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_23),
.B(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_16),
.B(n_3),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_55),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_57),
.B(n_65),
.Y(n_101)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

CKINVDCx6p67_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_69),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_61),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_25),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_28),
.B1(n_21),
.B2(n_33),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_66),
.A2(n_81),
.B1(n_70),
.B2(n_64),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_21),
.B1(n_27),
.B2(n_34),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_72),
.B1(n_75),
.B2(n_79),
.Y(n_88)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_38),
.B(n_50),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_71),
.B(n_14),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_39),
.A2(n_24),
.B1(n_16),
.B2(n_29),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_29),
.B1(n_24),
.B2(n_32),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_80),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_32),
.B1(n_18),
.B2(n_19),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_36),
.A2(n_22),
.B1(n_19),
.B2(n_26),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_17),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_86),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_17),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_22),
.B1(n_30),
.B2(n_5),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_92),
.B1(n_94),
.B2(n_70),
.Y(n_115)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

AO21x1_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_91),
.B(n_93),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_3),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_80),
.Y(n_127)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_63),
.A2(n_8),
.B1(n_9),
.B2(n_14),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_64),
.B1(n_73),
.B2(n_62),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_9),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_53),
.Y(n_124)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_52),
.B(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_103),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_112),
.Y(n_143)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_116),
.B1(n_94),
.B2(n_88),
.Y(n_132)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_120),
.Y(n_131)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_76),
.B(n_80),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_92),
.B(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_86),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_126),
.C(n_129),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_60),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_127),
.B(n_68),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_60),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_136),
.B1(n_137),
.B2(n_142),
.Y(n_156)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_101),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_133),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_93),
.B(n_85),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_130),
.B(n_124),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_129),
.A2(n_87),
.B1(n_102),
.B2(n_108),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_128),
.A2(n_102),
.B1(n_108),
.B2(n_91),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_145),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_128),
.A2(n_105),
.B1(n_82),
.B2(n_83),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_101),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_147),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_83),
.C(n_89),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_148),
.B(n_126),
.C(n_145),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_153),
.C(n_160),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_141),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_117),
.C(n_125),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_SL g168 ( 
.A1(n_154),
.A2(n_155),
.B(n_138),
.C(n_135),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_115),
.B1(n_118),
.B2(n_113),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_122),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_159),
.Y(n_164)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_117),
.C(n_121),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_111),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_163),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_134),
.B(n_110),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_152),
.B(n_150),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_167),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_148),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_175),
.B1(n_136),
.B2(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_139),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_174),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_111),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_144),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_160),
.C(n_146),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_179),
.C(n_181),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_154),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_134),
.C(n_161),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_182),
.A2(n_168),
.B(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

AOI31xp67_ASAP7_75t_L g185 ( 
.A1(n_181),
.A2(n_161),
.A3(n_155),
.B(n_172),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_186),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_118),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_183),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_188),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_177),
.A2(n_174),
.B(n_164),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_176),
.C(n_178),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_137),
.C(n_142),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_192),
.A2(n_170),
.B1(n_179),
.B2(n_178),
.Y(n_194)
);

INVxp33_ASAP7_75t_L g196 ( 
.A(n_194),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_191),
.B(n_190),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_195),
.Y(n_198)
);


endmodule