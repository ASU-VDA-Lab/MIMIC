module real_aes_16115_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_1797;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_1034;
wire n_571;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1845;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_1441;
wire n_951;
wire n_875;
wire n_1199;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_1883;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_346;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1853;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_1172;
wire n_459;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1827;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1855;
wire n_1056;
wire n_1802;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_1226;
wire n_525;
wire n_1790;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_1192;
wire n_518;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_372;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_559;
wire n_1584;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_430;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_1430;
wire n_907;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1877;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1868;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_1352;
wire n_729;
wire n_394;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g1099 ( .A(n_0), .Y(n_1099) );
INVx1_ASAP7_75t_L g783 ( .A(n_1), .Y(n_783) );
OAI211xp5_ASAP7_75t_L g823 ( .A1(n_1), .A2(n_824), .B(n_825), .C(n_832), .Y(n_823) );
INVx1_ASAP7_75t_L g359 ( .A(n_2), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_2), .B(n_369), .Y(n_449) );
AND2x2_ASAP7_75t_L g558 ( .A(n_2), .B(n_517), .Y(n_558) );
AND2x2_ASAP7_75t_L g575 ( .A(n_2), .B(n_263), .Y(n_575) );
OAI211xp5_ASAP7_75t_SL g1119 ( .A1(n_3), .A2(n_847), .B(n_896), .C(n_1120), .Y(n_1119) );
INVx1_ASAP7_75t_L g1134 ( .A(n_3), .Y(n_1134) );
INVx1_ASAP7_75t_L g496 ( .A(n_4), .Y(n_496) );
INVx1_ASAP7_75t_L g1420 ( .A(n_5), .Y(n_1420) );
INVx1_ASAP7_75t_L g1145 ( .A(n_6), .Y(n_1145) );
AOI22xp5_ASAP7_75t_L g1579 ( .A1(n_7), .A2(n_69), .B1(n_1562), .B2(n_1580), .Y(n_1579) );
OAI211xp5_ASAP7_75t_L g482 ( .A1(n_8), .A2(n_483), .B(n_486), .C(n_490), .Y(n_482) );
INVx1_ASAP7_75t_L g539 ( .A(n_8), .Y(n_539) );
INVx1_ASAP7_75t_L g1512 ( .A(n_9), .Y(n_1512) );
AOI22xp33_ASAP7_75t_L g1418 ( .A1(n_10), .A2(n_81), .B1(n_642), .B2(n_806), .Y(n_1418) );
AOI221xp5_ASAP7_75t_L g1435 ( .A1(n_10), .A2(n_21), .B1(n_985), .B2(n_1436), .C(n_1438), .Y(n_1435) );
INVx1_ASAP7_75t_L g1462 ( .A(n_11), .Y(n_1462) );
OAI22xp5_ASAP7_75t_L g1534 ( .A1(n_12), .A2(n_46), .B1(n_475), .B2(n_1535), .Y(n_1534) );
OAI22xp5_ASAP7_75t_L g1543 ( .A1(n_12), .A2(n_46), .B1(n_1032), .B2(n_1544), .Y(n_1543) );
INVx1_ASAP7_75t_L g691 ( .A(n_13), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_14), .A2(n_183), .B1(n_813), .B2(n_815), .Y(n_812) );
INVx1_ASAP7_75t_L g826 ( .A(n_14), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g1364 ( .A1(n_15), .A2(n_28), .B1(n_766), .B2(n_1365), .Y(n_1364) );
INVx1_ASAP7_75t_L g1398 ( .A(n_15), .Y(n_1398) );
OAI211xp5_ASAP7_75t_L g947 ( .A1(n_16), .A2(n_867), .B(n_948), .C(n_950), .Y(n_947) );
INVx1_ASAP7_75t_L g958 ( .A(n_16), .Y(n_958) );
INVx1_ASAP7_75t_L g1192 ( .A(n_17), .Y(n_1192) );
INVx1_ASAP7_75t_L g1174 ( .A(n_18), .Y(n_1174) );
OAI211xp5_ASAP7_75t_L g1181 ( .A1(n_18), .A2(n_867), .B(n_1182), .C(n_1183), .Y(n_1181) );
INVx1_ASAP7_75t_L g1248 ( .A(n_19), .Y(n_1248) );
INVx1_ASAP7_75t_L g1148 ( .A(n_20), .Y(n_1148) );
AOI22xp33_ASAP7_75t_SL g1427 ( .A1(n_21), .A2(n_250), .B1(n_643), .B2(n_1365), .Y(n_1427) );
INVx1_ASAP7_75t_L g930 ( .A(n_22), .Y(n_930) );
INVx2_ASAP7_75t_L g420 ( .A(n_23), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_24), .A2(n_343), .B1(n_749), .B2(n_750), .Y(n_748) );
INVx1_ASAP7_75t_L g761 ( .A(n_24), .Y(n_761) );
OAI22xp33_ASAP7_75t_L g1215 ( .A1(n_25), .A2(n_291), .B1(n_361), .B2(n_859), .Y(n_1215) );
OAI22xp5_ASAP7_75t_L g1224 ( .A1(n_25), .A2(n_291), .B1(n_1225), .B2(n_1226), .Y(n_1224) );
INVx1_ASAP7_75t_L g621 ( .A(n_26), .Y(n_621) );
INVx1_ASAP7_75t_L g1102 ( .A(n_27), .Y(n_1102) );
AOI221xp5_ASAP7_75t_L g1378 ( .A1(n_28), .A2(n_45), .B1(n_750), .B2(n_1379), .C(n_1381), .Y(n_1378) );
INVx1_ASAP7_75t_L g1424 ( .A(n_29), .Y(n_1424) );
INVx1_ASAP7_75t_L g1476 ( .A(n_30), .Y(n_1476) );
AOI22xp5_ASAP7_75t_L g1589 ( .A1(n_31), .A2(n_234), .B1(n_1569), .B2(n_1572), .Y(n_1589) );
INVx1_ASAP7_75t_L g1156 ( .A(n_32), .Y(n_1156) );
OA222x2_ASAP7_75t_L g1280 ( .A1(n_33), .A2(n_90), .B1(n_257), .B2(n_1281), .C1(n_1283), .C2(n_1287), .Y(n_1280) );
INVx1_ASAP7_75t_L g1337 ( .A(n_33), .Y(n_1337) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_34), .Y(n_354) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_34), .B(n_352), .Y(n_1563) );
AOI22xp5_ASAP7_75t_L g1578 ( .A1(n_35), .A2(n_211), .B1(n_1569), .B2(n_1572), .Y(n_1578) );
AOI22xp33_ASAP7_75t_L g1849 ( .A1(n_36), .A2(n_325), .B1(n_556), .B2(n_831), .Y(n_1849) );
INVxp67_ASAP7_75t_SL g1866 ( .A(n_36), .Y(n_1866) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_37), .A2(n_218), .B1(n_728), .B2(n_729), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_37), .A2(n_277), .B1(n_773), .B2(n_775), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g1366 ( .A1(n_38), .A2(n_226), .B1(n_645), .B2(n_1006), .Y(n_1366) );
INVx1_ASAP7_75t_L g1383 ( .A(n_38), .Y(n_1383) );
AOI22xp5_ASAP7_75t_L g1614 ( .A1(n_39), .A2(n_283), .B1(n_1569), .B2(n_1572), .Y(n_1614) );
INVx1_ASAP7_75t_L g700 ( .A(n_40), .Y(n_700) );
INVx1_ASAP7_75t_L g1513 ( .A(n_41), .Y(n_1513) );
INVx1_ASAP7_75t_L g1200 ( .A(n_42), .Y(n_1200) );
XNOR2xp5_ASAP7_75t_L g917 ( .A(n_43), .B(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g1039 ( .A(n_44), .Y(n_1039) );
AOI22xp33_ASAP7_75t_SL g1370 ( .A1(n_45), .A2(n_319), .B1(n_656), .B2(n_1365), .Y(n_1370) );
INVxp67_ASAP7_75t_SL g1423 ( .A(n_47), .Y(n_1423) );
OAI22xp5_ASAP7_75t_L g1443 ( .A1(n_47), .A2(n_182), .B1(n_465), .B2(n_1444), .Y(n_1443) );
AOI22xp5_ASAP7_75t_L g1585 ( .A1(n_48), .A2(n_124), .B1(n_1569), .B2(n_1572), .Y(n_1585) );
INVx1_ASAP7_75t_L g382 ( .A(n_49), .Y(n_382) );
INVx1_ASAP7_75t_L g1471 ( .A(n_50), .Y(n_1471) );
INVx1_ASAP7_75t_L g1048 ( .A(n_51), .Y(n_1048) );
OAI211xp5_ASAP7_75t_L g844 ( .A1(n_52), .A2(n_845), .B(n_847), .C(n_848), .Y(n_844) );
INVx1_ASAP7_75t_L g870 ( .A(n_52), .Y(n_870) );
INVx1_ASAP7_75t_L g1244 ( .A(n_53), .Y(n_1244) );
OAI211xp5_ASAP7_75t_L g1216 ( .A1(n_54), .A2(n_956), .B(n_1026), .C(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1229 ( .A(n_54), .Y(n_1229) );
CKINVDCx5p33_ASAP7_75t_R g1305 ( .A(n_55), .Y(n_1305) );
INVx1_ASAP7_75t_L g1431 ( .A(n_56), .Y(n_1431) );
INVx1_ASAP7_75t_L g800 ( .A(n_57), .Y(n_800) );
AOI21xp33_ASAP7_75t_L g833 ( .A1(n_57), .A2(n_564), .B(n_603), .Y(n_833) );
AOI22xp5_ASAP7_75t_L g1583 ( .A1(n_58), .A2(n_188), .B1(n_1562), .B2(n_1584), .Y(n_1583) );
NAND5xp2_ASAP7_75t_L g1788 ( .A(n_58), .B(n_1789), .C(n_1804), .D(n_1815), .E(n_1817), .Y(n_1788) );
INVx1_ASAP7_75t_L g1823 ( .A(n_58), .Y(n_1823) );
AOI22xp33_ASAP7_75t_L g1833 ( .A1(n_58), .A2(n_1834), .B1(n_1837), .B2(n_1886), .Y(n_1833) );
AOI22xp33_ASAP7_75t_SL g1854 ( .A1(n_59), .A2(n_272), .B1(n_831), .B2(n_1855), .Y(n_1854) );
AOI22xp33_ASAP7_75t_L g1867 ( .A1(n_59), .A2(n_253), .B1(n_1327), .B2(n_1811), .Y(n_1867) );
OAI22xp33_ASAP7_75t_L g501 ( .A1(n_60), .A2(n_148), .B1(n_502), .B2(n_504), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_60), .A2(n_148), .B1(n_541), .B2(n_543), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g1422 ( .A(n_61), .Y(n_1422) );
INVx1_ASAP7_75t_L g1453 ( .A(n_62), .Y(n_1453) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_63), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g1367 ( .A1(n_64), .A2(n_76), .B1(n_651), .B2(n_1368), .Y(n_1367) );
INVx1_ASAP7_75t_L g1382 ( .A(n_64), .Y(n_1382) );
INVx1_ASAP7_75t_L g887 ( .A(n_65), .Y(n_887) );
OAI22xp33_ASAP7_75t_SL g1845 ( .A1(n_66), .A2(n_260), .B1(n_894), .B2(n_1304), .Y(n_1845) );
INVx1_ASAP7_75t_L g1878 ( .A(n_66), .Y(n_1878) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_67), .A2(n_114), .B1(n_568), .B2(n_572), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_67), .A2(n_243), .B1(n_645), .B2(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g792 ( .A(n_68), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_68), .A2(n_313), .B1(n_821), .B2(n_822), .Y(n_820) );
XNOR2xp5_ASAP7_75t_L g1457 ( .A(n_69), .B(n_1458), .Y(n_1457) );
AOI21xp33_ASAP7_75t_L g993 ( .A1(n_70), .A2(n_726), .B(n_994), .Y(n_993) );
AOI221xp5_ASAP7_75t_L g1012 ( .A1(n_70), .A2(n_279), .B1(n_1006), .B2(n_1013), .C(n_1015), .Y(n_1012) );
CKINVDCx5p33_ASAP7_75t_R g1358 ( .A(n_71), .Y(n_1358) );
XOR2x2_ASAP7_75t_L g550 ( .A(n_72), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g1195 ( .A(n_73), .Y(n_1195) );
OAI222xp33_ASAP7_75t_L g971 ( .A1(n_74), .A2(n_87), .B1(n_95), .B2(n_628), .C1(n_972), .C2(n_973), .Y(n_971) );
AOI21xp33_ASAP7_75t_L g745 ( .A1(n_75), .A2(n_746), .B(n_747), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_75), .A2(n_218), .B1(n_763), .B2(n_766), .Y(n_762) );
INVx1_ASAP7_75t_L g1402 ( .A(n_76), .Y(n_1402) );
AOI22xp33_ASAP7_75t_L g1693 ( .A1(n_77), .A2(n_252), .B1(n_1562), .B2(n_1580), .Y(n_1693) );
INVx1_ASAP7_75t_L g1496 ( .A(n_78), .Y(n_1496) );
OAI211xp5_ASAP7_75t_L g1504 ( .A1(n_78), .A2(n_521), .B(n_1026), .C(n_1505), .Y(n_1504) );
INVx1_ASAP7_75t_L g1265 ( .A(n_79), .Y(n_1265) );
OAI211xp5_ASAP7_75t_L g1269 ( .A1(n_79), .A2(n_486), .B(n_1010), .C(n_1270), .Y(n_1269) );
AOI221xp5_ASAP7_75t_L g1793 ( .A1(n_80), .A2(n_186), .B1(n_528), .B2(n_603), .C(n_829), .Y(n_1793) );
AOI22xp33_ASAP7_75t_L g1809 ( .A1(n_80), .A2(n_245), .B1(n_645), .B2(n_771), .Y(n_1809) );
INVx1_ASAP7_75t_L g1452 ( .A(n_81), .Y(n_1452) );
AOI22xp33_ASAP7_75t_L g1794 ( .A1(n_82), .A2(n_245), .B1(n_750), .B2(n_1795), .Y(n_1794) );
AOI22xp33_ASAP7_75t_L g1808 ( .A1(n_82), .A2(n_186), .B1(n_771), .B2(n_1347), .Y(n_1808) );
OAI22xp33_ASAP7_75t_L g1033 ( .A1(n_83), .A2(n_89), .B1(n_1034), .B2(n_1035), .Y(n_1033) );
OAI22xp33_ASAP7_75t_L g1081 ( .A1(n_83), .A2(n_89), .B1(n_873), .B2(n_1082), .Y(n_1081) );
CKINVDCx5p33_ASAP7_75t_R g978 ( .A(n_84), .Y(n_978) );
CKINVDCx5p33_ASAP7_75t_R g718 ( .A(n_85), .Y(n_718) );
INVx1_ASAP7_75t_L g1243 ( .A(n_86), .Y(n_1243) );
AOI22xp5_ASAP7_75t_L g1838 ( .A1(n_88), .A2(n_1839), .B1(n_1884), .B2(n_1885), .Y(n_1838) );
CKINVDCx5p33_ASAP7_75t_R g1884 ( .A(n_88), .Y(n_1884) );
OAI221xp5_ASAP7_75t_L g1320 ( .A1(n_90), .A2(n_206), .B1(n_1321), .B2(n_1323), .C(n_1325), .Y(n_1320) );
OAI22xp5_ASAP7_75t_L g1391 ( .A1(n_91), .A2(n_306), .B1(n_442), .B2(n_465), .Y(n_1391) );
INVx1_ASAP7_75t_L g1404 ( .A(n_91), .Y(n_1404) );
INVx1_ASAP7_75t_L g1293 ( .A(n_92), .Y(n_1293) );
AOI22xp33_ASAP7_75t_L g1353 ( .A1(n_92), .A2(n_145), .B1(n_648), .B2(n_773), .Y(n_1353) );
CKINVDCx5p33_ASAP7_75t_R g1800 ( .A(n_93), .Y(n_1800) );
INVx1_ASAP7_75t_L g1057 ( .A(n_94), .Y(n_1057) );
OAI22xp5_ASAP7_75t_L g1001 ( .A1(n_95), .A2(n_338), .B1(n_822), .B2(n_1002), .Y(n_1001) );
OAI22xp5_ASAP7_75t_L g1221 ( .A1(n_96), .A2(n_180), .B1(n_541), .B2(n_1222), .Y(n_1221) );
OAI22xp33_ASAP7_75t_L g1230 ( .A1(n_96), .A2(n_180), .B1(n_502), .B2(n_1231), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g1598 ( .A1(n_97), .A2(n_189), .B1(n_1562), .B2(n_1569), .Y(n_1598) );
INVx1_ASAP7_75t_L g1094 ( .A(n_98), .Y(n_1094) );
INVx1_ASAP7_75t_L g1121 ( .A(n_99), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g1597 ( .A1(n_100), .A2(n_305), .B1(n_1572), .B2(n_1580), .Y(n_1597) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_101), .A2(n_169), .B1(n_729), .B2(n_749), .Y(n_995) );
INVx1_ASAP7_75t_L g1008 ( .A(n_101), .Y(n_1008) );
INVx1_ASAP7_75t_L g1469 ( .A(n_102), .Y(n_1469) );
XNOR2xp5_ASAP7_75t_L g1233 ( .A(n_103), .B(n_1234), .Y(n_1233) );
AOI22xp5_ASAP7_75t_L g1561 ( .A1(n_103), .A2(n_167), .B1(n_1562), .B2(n_1566), .Y(n_1561) );
XNOR2xp5_ASAP7_75t_L g377 ( .A(n_104), .B(n_378), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g1430 ( .A(n_105), .Y(n_1430) );
AOI22xp33_ASAP7_75t_L g1426 ( .A1(n_106), .A2(n_324), .B1(n_646), .B2(n_1368), .Y(n_1426) );
AOI221xp5_ASAP7_75t_L g1449 ( .A1(n_106), .A2(n_222), .B1(n_750), .B2(n_831), .C(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g400 ( .A(n_107), .Y(n_400) );
OAI211xp5_ASAP7_75t_L g1798 ( .A1(n_108), .A2(n_998), .B(n_1063), .C(n_1799), .Y(n_1798) );
INVx1_ASAP7_75t_L g1819 ( .A(n_108), .Y(n_1819) );
AOI22xp33_ASAP7_75t_L g1694 ( .A1(n_109), .A2(n_330), .B1(n_1569), .B2(n_1572), .Y(n_1694) );
INVx1_ASAP7_75t_L g1406 ( .A(n_110), .Y(n_1406) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_111), .A2(n_154), .B1(n_1031), .B2(n_1032), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_111), .A2(n_154), .B1(n_1074), .B2(n_1076), .Y(n_1073) );
OAI22xp33_ASAP7_75t_L g1167 ( .A1(n_112), .A2(n_120), .B1(n_514), .B2(n_1127), .Y(n_1167) );
OAI22xp33_ASAP7_75t_L g1178 ( .A1(n_112), .A2(n_120), .B1(n_1074), .B2(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g1218 ( .A(n_113), .Y(n_1218) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_114), .A2(n_135), .B1(n_384), .B2(n_651), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g953 ( .A1(n_115), .A2(n_194), .B1(n_478), .B2(n_873), .Y(n_953) );
OAI22xp5_ASAP7_75t_L g960 ( .A1(n_115), .A2(n_233), .B1(n_541), .B2(n_961), .Y(n_960) );
INVx1_ASAP7_75t_L g811 ( .A(n_116), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_116), .A2(n_264), .B1(n_556), .B2(n_831), .Y(n_830) );
CKINVDCx5p33_ASAP7_75t_R g716 ( .A(n_117), .Y(n_716) );
INVx1_ASAP7_75t_L g352 ( .A(n_118), .Y(n_352) );
INVx1_ASAP7_75t_L g1468 ( .A(n_119), .Y(n_1468) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_121), .A2(n_178), .B1(n_623), .B2(n_628), .Y(n_622) );
INVx1_ASAP7_75t_L g926 ( .A(n_122), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_123), .A2(n_340), .B1(n_854), .B2(n_856), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_123), .A2(n_134), .B1(n_862), .B2(n_863), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g1266 ( .A1(n_125), .A2(n_165), .B1(n_541), .B2(n_1222), .Y(n_1266) );
OAI22xp33_ASAP7_75t_L g1272 ( .A1(n_125), .A2(n_165), .B1(n_502), .B2(n_504), .Y(n_1272) );
INVxp67_ASAP7_75t_SL g599 ( .A(n_126), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_126), .A2(n_284), .B1(n_642), .B2(n_656), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g1844 ( .A1(n_127), .A2(n_159), .B1(n_1294), .B2(n_1295), .Y(n_1844) );
NOR2xp33_ASAP7_75t_L g1882 ( .A(n_127), .B(n_863), .Y(n_1882) );
INVx1_ASAP7_75t_L g1107 ( .A(n_128), .Y(n_1107) );
CKINVDCx5p33_ASAP7_75t_R g1375 ( .A(n_129), .Y(n_1375) );
INVx1_ASAP7_75t_L g1104 ( .A(n_130), .Y(n_1104) );
INVx1_ASAP7_75t_L g1106 ( .A(n_131), .Y(n_1106) );
OAI22xp5_ASAP7_75t_L g1125 ( .A1(n_132), .A2(n_142), .B1(n_542), .B2(n_856), .Y(n_1125) );
OAI22xp33_ASAP7_75t_L g1135 ( .A1(n_132), .A2(n_142), .B1(n_946), .B2(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g1196 ( .A(n_133), .Y(n_1196) );
OAI22xp33_ASAP7_75t_L g858 ( .A1(n_134), .A2(n_323), .B1(n_361), .B2(n_859), .Y(n_858) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_135), .A2(n_243), .B1(n_564), .B2(n_601), .C(n_603), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g1175 ( .A1(n_136), .A2(n_295), .B1(n_541), .B2(n_856), .Y(n_1175) );
OAI22xp5_ASAP7_75t_L g1180 ( .A1(n_136), .A2(n_295), .B1(n_504), .B2(n_1082), .Y(n_1180) );
INVx1_ASAP7_75t_L g1173 ( .A(n_137), .Y(n_1173) );
INVx1_ASAP7_75t_L g1124 ( .A(n_138), .Y(n_1124) );
OAI211xp5_ASAP7_75t_L g1130 ( .A1(n_138), .A2(n_867), .B(n_1131), .C(n_1133), .Y(n_1130) );
INVx1_ASAP7_75t_L g1095 ( .A(n_139), .Y(n_1095) );
INVx1_ASAP7_75t_L g1139 ( .A(n_140), .Y(n_1139) );
AOI22xp33_ASAP7_75t_SL g1613 ( .A1(n_140), .A2(n_225), .B1(n_1562), .B2(n_1580), .Y(n_1613) );
AOI22xp33_ASAP7_75t_SL g804 ( .A1(n_141), .A2(n_285), .B1(n_805), .B2(n_806), .Y(n_804) );
AOI21xp33_ASAP7_75t_L g828 ( .A1(n_141), .A2(n_747), .B(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g1264 ( .A(n_143), .Y(n_1264) );
INVx1_ASAP7_75t_L g1539 ( .A(n_144), .Y(n_1539) );
OAI211xp5_ASAP7_75t_L g1546 ( .A1(n_144), .A2(n_890), .B(n_1547), .C(n_1548), .Y(n_1546) );
AOI22xp33_ASAP7_75t_L g1306 ( .A1(n_145), .A2(n_191), .B1(n_568), .B2(n_572), .Y(n_1306) );
INVx1_ASAP7_75t_L g1239 ( .A(n_146), .Y(n_1239) );
AOI221xp5_ASAP7_75t_L g560 ( .A1(n_147), .A2(n_284), .B1(n_561), .B2(n_562), .C(n_566), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_147), .A2(n_247), .B1(n_640), .B2(n_643), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g1312 ( .A1(n_149), .A2(n_206), .B1(n_624), .B2(n_1313), .Y(n_1312) );
INVx1_ASAP7_75t_L g1338 ( .A(n_149), .Y(n_1338) );
INVx1_ASAP7_75t_L g1518 ( .A(n_150), .Y(n_1518) );
OAI22xp33_ASAP7_75t_L g1126 ( .A1(n_151), .A2(n_254), .B1(n_859), .B2(n_1127), .Y(n_1126) );
OAI22xp33_ASAP7_75t_L g1129 ( .A1(n_151), .A2(n_254), .B1(n_477), .B2(n_1076), .Y(n_1129) );
INVx1_ASAP7_75t_L g1051 ( .A(n_152), .Y(n_1051) );
INVx1_ASAP7_75t_L g934 ( .A(n_153), .Y(n_934) );
OAI221xp5_ASAP7_75t_L g1858 ( .A1(n_155), .A2(n_326), .B1(n_1859), .B2(n_1860), .C(n_1861), .Y(n_1858) );
INVx1_ASAP7_75t_L g1875 ( .A(n_155), .Y(n_1875) );
INVx1_ASAP7_75t_L g1847 ( .A(n_156), .Y(n_1847) );
AOI22xp33_ASAP7_75t_L g1871 ( .A1(n_156), .A2(n_272), .B1(n_1327), .B2(n_1807), .Y(n_1871) );
INVx1_ASAP7_75t_L g436 ( .A(n_157), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g1851 ( .A(n_158), .Y(n_1851) );
INVx1_ASAP7_75t_L g1877 ( .A(n_159), .Y(n_1877) );
INVx1_ASAP7_75t_L g422 ( .A(n_160), .Y(n_422) );
INVx1_ASAP7_75t_L g952 ( .A(n_161), .Y(n_952) );
OAI211xp5_ASAP7_75t_SL g955 ( .A1(n_161), .A2(n_847), .B(n_956), .C(n_957), .Y(n_955) );
INVx1_ASAP7_75t_L g1152 ( .A(n_162), .Y(n_1152) );
OAI22xp33_ASAP7_75t_L g1497 ( .A1(n_163), .A2(n_266), .B1(n_862), .B2(n_1179), .Y(n_1497) );
OAI22xp5_ASAP7_75t_L g1499 ( .A1(n_163), .A2(n_266), .B1(n_1032), .B2(n_1500), .Y(n_1499) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_164), .A2(n_233), .B1(n_862), .B2(n_946), .Y(n_945) );
OAI22xp33_ASAP7_75t_L g963 ( .A1(n_164), .A2(n_194), .B1(n_361), .B2(n_514), .Y(n_963) );
INVx1_ASAP7_75t_L g1466 ( .A(n_166), .Y(n_1466) );
INVx1_ASAP7_75t_L g1473 ( .A(n_168), .Y(n_1473) );
INVxp67_ASAP7_75t_SL g1016 ( .A(n_169), .Y(n_1016) );
INVx1_ASAP7_75t_L g1816 ( .A(n_170), .Y(n_1816) );
INVx1_ASAP7_75t_L g424 ( .A(n_171), .Y(n_424) );
OAI22xp33_ASAP7_75t_L g474 ( .A1(n_172), .A2(n_334), .B1(n_475), .B2(n_478), .Y(n_474) );
OAI22xp33_ASAP7_75t_L g513 ( .A1(n_172), .A2(n_334), .B1(n_361), .B2(n_514), .Y(n_513) );
OAI22xp33_ASAP7_75t_L g1491 ( .A1(n_173), .A2(n_203), .B1(n_502), .B2(n_873), .Y(n_1491) );
OAI22xp33_ASAP7_75t_L g1501 ( .A1(n_173), .A2(n_203), .B1(n_854), .B2(n_1502), .Y(n_1501) );
INVx1_ASAP7_75t_L g1203 ( .A(n_174), .Y(n_1203) );
OAI211xp5_ASAP7_75t_L g1168 ( .A1(n_175), .A2(n_890), .B(n_1169), .C(n_1172), .Y(n_1168) );
INVx1_ASAP7_75t_L g1184 ( .A(n_175), .Y(n_1184) );
INVx1_ASAP7_75t_L g1251 ( .A(n_176), .Y(n_1251) );
INVx1_ASAP7_75t_L g392 ( .A(n_177), .Y(n_392) );
OAI211xp5_ASAP7_75t_L g553 ( .A1(n_178), .A2(n_554), .B(n_559), .C(n_576), .Y(n_553) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_179), .A2(n_332), .B1(n_723), .B2(n_725), .C(n_726), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_179), .A2(n_343), .B1(n_770), .B2(n_771), .Y(n_769) );
XOR2x2_ASAP7_75t_L g1507 ( .A(n_181), .B(n_1508), .Y(n_1507) );
INVxp67_ASAP7_75t_SL g1433 ( .A(n_182), .Y(n_1433) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_183), .A2(n_285), .B1(n_556), .B2(n_831), .Y(n_834) );
CKINVDCx5p33_ASAP7_75t_R g1301 ( .A(n_184), .Y(n_1301) );
INVx1_ASAP7_75t_L g1538 ( .A(n_185), .Y(n_1538) );
INVx1_ASAP7_75t_L g1522 ( .A(n_187), .Y(n_1522) );
INVx1_ASAP7_75t_L g882 ( .A(n_190), .Y(n_882) );
INVx1_ASAP7_75t_L g1349 ( .A(n_191), .Y(n_1349) );
XNOR2xp5_ASAP7_75t_L g1186 ( .A(n_192), .B(n_1187), .Y(n_1186) );
INVx1_ASAP7_75t_L g849 ( .A(n_193), .Y(n_849) );
INVx1_ASAP7_75t_L g1250 ( .A(n_195), .Y(n_1250) );
INVx1_ASAP7_75t_L g992 ( .A(n_196), .Y(n_992) );
AOI221x1_ASAP7_75t_SL g1005 ( .A1(n_196), .A2(n_275), .B1(n_384), .B2(n_1006), .C(n_1007), .Y(n_1005) );
INVx1_ASAP7_75t_L g1144 ( .A(n_197), .Y(n_1144) );
AOI221x1_ASAP7_75t_SL g1289 ( .A1(n_198), .A2(n_269), .B1(n_1290), .B2(n_1291), .C(n_1292), .Y(n_1289) );
AOI21xp33_ASAP7_75t_L g1351 ( .A1(n_198), .A2(n_677), .B(n_1352), .Y(n_1351) );
OAI211xp5_ASAP7_75t_L g1790 ( .A1(n_199), .A2(n_822), .B(n_1791), .C(n_1797), .Y(n_1790) );
NOR2xp33_ASAP7_75t_L g1803 ( .A(n_199), .B(n_628), .Y(n_1803) );
INVx1_ASAP7_75t_L g577 ( .A(n_200), .Y(n_577) );
OAI22xp33_ASAP7_75t_L g669 ( .A1(n_200), .A2(n_309), .B1(n_670), .B2(n_674), .Y(n_669) );
AOI21xp33_ASAP7_75t_L g999 ( .A1(n_201), .A2(n_746), .B(n_747), .Y(n_999) );
INVx1_ASAP7_75t_L g1017 ( .A(n_201), .Y(n_1017) );
OAI221xp5_ASAP7_75t_L g584 ( .A1(n_202), .A2(n_270), .B1(n_585), .B2(n_589), .C(n_594), .Y(n_584) );
INVx1_ASAP7_75t_L g659 ( .A(n_202), .Y(n_659) );
INVx2_ASAP7_75t_L g1565 ( .A(n_204), .Y(n_1565) );
AND2x2_ASAP7_75t_L g1567 ( .A(n_204), .B(n_303), .Y(n_1567) );
AND2x2_ASAP7_75t_L g1573 ( .A(n_204), .B(n_1571), .Y(n_1573) );
INVx1_ASAP7_75t_L g889 ( .A(n_205), .Y(n_889) );
OAI22xp33_ASAP7_75t_L g1540 ( .A1(n_207), .A2(n_268), .B1(n_1136), .B2(n_1541), .Y(n_1540) );
OAI22xp33_ASAP7_75t_L g1550 ( .A1(n_207), .A2(n_268), .B1(n_541), .B2(n_1035), .Y(n_1550) );
INVx1_ASAP7_75t_L g895 ( .A(n_208), .Y(n_895) );
INVx1_ASAP7_75t_L g1028 ( .A(n_209), .Y(n_1028) );
AOI22xp5_ASAP7_75t_L g1591 ( .A1(n_210), .A2(n_261), .B1(n_1562), .B2(n_1572), .Y(n_1591) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_212), .A2(n_689), .B1(n_776), .B2(n_777), .Y(n_688) );
INVxp67_ASAP7_75t_L g777 ( .A(n_212), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g1297 ( .A(n_213), .Y(n_1297) );
AOI22xp33_ASAP7_75t_L g1592 ( .A1(n_214), .A2(n_219), .B1(n_1566), .B2(n_1569), .Y(n_1592) );
INVx1_ASAP7_75t_L g902 ( .A(n_215), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g1792 ( .A1(n_216), .A2(n_287), .B1(n_750), .B2(n_831), .Y(n_1792) );
AOI22xp33_ASAP7_75t_SL g1810 ( .A1(n_216), .A2(n_302), .B1(n_1365), .B2(n_1811), .Y(n_1810) );
OAI211xp5_ASAP7_75t_L g1025 ( .A1(n_217), .A2(n_928), .B(n_1026), .C(n_1027), .Y(n_1025) );
INVx1_ASAP7_75t_L g1080 ( .A(n_217), .Y(n_1080) );
INVx1_ASAP7_75t_L g1191 ( .A(n_220), .Y(n_1191) );
OAI221xp5_ASAP7_75t_SL g710 ( .A1(n_221), .A2(n_296), .B1(n_711), .B2(n_713), .C(n_715), .Y(n_710) );
INVx1_ASAP7_75t_L g737 ( .A(n_221), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g1417 ( .A1(n_222), .A2(n_310), .B1(n_384), .B2(n_651), .Y(n_1417) );
XNOR2xp5_ASAP7_75t_L g841 ( .A(n_223), .B(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g1515 ( .A(n_224), .Y(n_1515) );
INVx1_ASAP7_75t_L g1400 ( .A(n_226), .Y(n_1400) );
CKINVDCx5p33_ASAP7_75t_R g1801 ( .A(n_227), .Y(n_1801) );
INVx1_ASAP7_75t_L g1516 ( .A(n_228), .Y(n_1516) );
INVx2_ASAP7_75t_L g419 ( .A(n_229), .Y(n_419) );
INVx1_ASAP7_75t_L g431 ( .A(n_229), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_229), .B(n_420), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g1568 ( .A1(n_230), .A2(n_335), .B1(n_1569), .B2(n_1572), .Y(n_1568) );
INVx1_ASAP7_75t_L g405 ( .A(n_231), .Y(n_405) );
INVx1_ASAP7_75t_L g1157 ( .A(n_232), .Y(n_1157) );
INVx1_ASAP7_75t_L g951 ( .A(n_235), .Y(n_951) );
INVx1_ASAP7_75t_L g969 ( .A(n_236), .Y(n_969) );
OAI22xp5_ASAP7_75t_L g1802 ( .A1(n_237), .A2(n_308), .B1(n_928), .B2(n_1063), .Y(n_1802) );
INVx1_ASAP7_75t_L g1818 ( .A(n_237), .Y(n_1818) );
INVx1_ASAP7_75t_L g905 ( .A(n_238), .Y(n_905) );
INVx1_ASAP7_75t_L g1149 ( .A(n_239), .Y(n_1149) );
INVx1_ASAP7_75t_L g933 ( .A(n_240), .Y(n_933) );
OAI22xp33_ASAP7_75t_L g1261 ( .A1(n_241), .A2(n_265), .B1(n_361), .B2(n_859), .Y(n_1261) );
OAI22xp5_ASAP7_75t_L g1268 ( .A1(n_241), .A2(n_265), .B1(n_1179), .B2(n_1225), .Y(n_1268) );
BUFx3_ASAP7_75t_L g391 ( .A(n_242), .Y(n_391) );
INVx1_ASAP7_75t_L g694 ( .A(n_244), .Y(n_694) );
INVx1_ASAP7_75t_L g1524 ( .A(n_246), .Y(n_1524) );
INVxp67_ASAP7_75t_SL g597 ( .A(n_247), .Y(n_597) );
INVx1_ASAP7_75t_L g1198 ( .A(n_248), .Y(n_1198) );
OAI22xp5_ASAP7_75t_SL g980 ( .A1(n_249), .A2(n_286), .B1(n_613), .B2(n_626), .Y(n_980) );
CKINVDCx5p33_ASAP7_75t_R g990 ( .A(n_249), .Y(n_990) );
INVx1_ASAP7_75t_L g1451 ( .A(n_250), .Y(n_1451) );
INVx1_ASAP7_75t_L g1220 ( .A(n_251), .Y(n_1220) );
OAI211xp5_ASAP7_75t_SL g1227 ( .A1(n_251), .A2(n_867), .B(n_1010), .C(n_1228), .Y(n_1227) );
AOI21xp33_ASAP7_75t_L g1848 ( .A1(n_253), .A2(n_746), .B(n_747), .Y(n_1848) );
INVx1_ASAP7_75t_L g1047 ( .A(n_255), .Y(n_1047) );
INVx1_ASAP7_75t_L g931 ( .A(n_256), .Y(n_931) );
INVx1_ASAP7_75t_L g1326 ( .A(n_257), .Y(n_1326) );
INVx1_ASAP7_75t_L g788 ( .A(n_258), .Y(n_788) );
INVx1_ASAP7_75t_L g1475 ( .A(n_259), .Y(n_1475) );
INVx1_ASAP7_75t_L g1881 ( .A(n_260), .Y(n_1881) );
INVx1_ASAP7_75t_L g878 ( .A(n_262), .Y(n_878) );
BUFx3_ASAP7_75t_L g369 ( .A(n_263), .Y(n_369) );
INVx1_ASAP7_75t_L g517 ( .A(n_263), .Y(n_517) );
INVx1_ASAP7_75t_L g803 ( .A(n_264), .Y(n_803) );
XNOR2xp5_ASAP7_75t_L g1088 ( .A(n_267), .B(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g1348 ( .A(n_269), .Y(n_1348) );
INVx1_ASAP7_75t_L g664 ( .A(n_270), .Y(n_664) );
INVx1_ASAP7_75t_L g923 ( .A(n_271), .Y(n_923) );
INVx1_ASAP7_75t_L g1278 ( .A(n_273), .Y(n_1278) );
INVx1_ASAP7_75t_L g924 ( .A(n_274), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_275), .A2(n_279), .B1(n_729), .B2(n_749), .Y(n_1000) );
INVx1_ASAP7_75t_L g1100 ( .A(n_276), .Y(n_1100) );
INVx1_ASAP7_75t_L g744 ( .A(n_277), .Y(n_744) );
INVx1_ASAP7_75t_L g1029 ( .A(n_278), .Y(n_1029) );
OAI211xp5_ASAP7_75t_L g1077 ( .A1(n_278), .A2(n_406), .B(n_486), .C(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g1246 ( .A(n_280), .Y(n_1246) );
INVx1_ASAP7_75t_L g1052 ( .A(n_281), .Y(n_1052) );
CKINVDCx5p33_ASAP7_75t_R g1376 ( .A(n_282), .Y(n_1376) );
INVx1_ASAP7_75t_L g984 ( .A(n_286), .Y(n_984) );
AOI22xp33_ASAP7_75t_SL g1806 ( .A1(n_287), .A2(n_342), .B1(n_1365), .B2(n_1807), .Y(n_1806) );
INVx1_ASAP7_75t_L g389 ( .A(n_288), .Y(n_389) );
INVx1_ASAP7_75t_L g398 ( .A(n_288), .Y(n_398) );
INVx1_ASAP7_75t_L g500 ( .A(n_289), .Y(n_500) );
OAI211xp5_ASAP7_75t_L g520 ( .A1(n_289), .A2(n_521), .B(n_525), .C(n_530), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_290), .A2(n_779), .B1(n_780), .B2(n_839), .Y(n_778) );
INVxp67_ASAP7_75t_L g839 ( .A(n_290), .Y(n_839) );
INVxp67_ASAP7_75t_SL g784 ( .A(n_292), .Y(n_784) );
OAI221xp5_ASAP7_75t_L g836 ( .A1(n_292), .A2(n_333), .B1(n_590), .B2(n_620), .C(n_837), .Y(n_836) );
OAI211xp5_ASAP7_75t_L g1262 ( .A1(n_293), .A2(n_956), .B(n_1026), .C(n_1263), .Y(n_1262) );
INVx1_ASAP7_75t_L g1271 ( .A(n_293), .Y(n_1271) );
INVx1_ASAP7_75t_L g997 ( .A(n_294), .Y(n_997) );
INVx1_ASAP7_75t_L g753 ( .A(n_296), .Y(n_753) );
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_297), .Y(n_789) );
INVx1_ASAP7_75t_L g1495 ( .A(n_298), .Y(n_1495) );
INVx1_ASAP7_75t_L g1520 ( .A(n_299), .Y(n_1520) );
AOI22xp5_ASAP7_75t_L g1021 ( .A1(n_300), .A2(n_1022), .B1(n_1023), .B2(n_1083), .Y(n_1021) );
INVxp67_ASAP7_75t_SL g1083 ( .A(n_300), .Y(n_1083) );
AOI22xp5_ASAP7_75t_SL g1588 ( .A1(n_300), .A2(n_339), .B1(n_1562), .B2(n_1566), .Y(n_1588) );
CKINVDCx5p33_ASAP7_75t_R g1372 ( .A(n_301), .Y(n_1372) );
AOI221xp5_ASAP7_75t_SL g1796 ( .A1(n_302), .A2(n_342), .B1(n_528), .B2(n_564), .C(n_747), .Y(n_1796) );
AND2x2_ASAP7_75t_L g1564 ( .A(n_303), .B(n_1565), .Y(n_1564) );
INVx1_ASAP7_75t_L g1571 ( .A(n_303), .Y(n_1571) );
OAI211xp5_ASAP7_75t_SL g1492 ( .A1(n_304), .A2(n_486), .B(n_1493), .C(n_1494), .Y(n_1492) );
INVx1_ASAP7_75t_L g1506 ( .A(n_304), .Y(n_1506) );
INVx1_ASAP7_75t_L g1361 ( .A(n_306), .Y(n_1361) );
OAI211xp5_ASAP7_75t_L g1536 ( .A1(n_307), .A2(n_867), .B(n_1018), .C(n_1537), .Y(n_1536) );
INVx1_ASAP7_75t_L g1549 ( .A(n_307), .Y(n_1549) );
INVx1_ASAP7_75t_L g1814 ( .A(n_308), .Y(n_1814) );
INVx1_ASAP7_75t_L g580 ( .A(n_309), .Y(n_580) );
INVx1_ASAP7_75t_L g1440 ( .A(n_310), .Y(n_1440) );
INVx1_ASAP7_75t_L g897 ( .A(n_311), .Y(n_897) );
INVx1_ASAP7_75t_L g852 ( .A(n_312), .Y(n_852) );
OAI211xp5_ASAP7_75t_L g864 ( .A1(n_312), .A2(n_865), .B(n_867), .C(n_868), .Y(n_864) );
INVx1_ASAP7_75t_L g794 ( .A(n_313), .Y(n_794) );
INVx1_ASAP7_75t_L g1857 ( .A(n_314), .Y(n_1857) );
INVx1_ASAP7_75t_L g1240 ( .A(n_315), .Y(n_1240) );
INVx1_ASAP7_75t_L g434 ( .A(n_316), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g809 ( .A(n_317), .Y(n_809) );
INVx1_ASAP7_75t_L g927 ( .A(n_318), .Y(n_927) );
AOI211xp5_ASAP7_75t_SL g1395 ( .A1(n_319), .A2(n_1396), .B(n_1397), .C(n_1399), .Y(n_1395) );
INVx1_ASAP7_75t_L g1154 ( .A(n_320), .Y(n_1154) );
AOI21xp5_ASAP7_75t_SL g1852 ( .A1(n_321), .A2(n_746), .B(n_1853), .Y(n_1852) );
INVx1_ASAP7_75t_L g1865 ( .A(n_321), .Y(n_1865) );
INVx1_ASAP7_75t_L g1204 ( .A(n_322), .Y(n_1204) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_323), .A2(n_340), .B1(n_872), .B2(n_873), .Y(n_871) );
INVx1_ASAP7_75t_L g1439 ( .A(n_324), .Y(n_1439) );
INVxp67_ASAP7_75t_L g1870 ( .A(n_325), .Y(n_1870) );
INVxp67_ASAP7_75t_SL g1880 ( .A(n_326), .Y(n_1880) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_327), .Y(n_365) );
INVx1_ASAP7_75t_L g1042 ( .A(n_328), .Y(n_1042) );
INVx1_ASAP7_75t_L g1058 ( .A(n_329), .Y(n_1058) );
CKINVDCx5p33_ASAP7_75t_R g1317 ( .A(n_331), .Y(n_1317) );
INVx1_ASAP7_75t_L g760 ( .A(n_332), .Y(n_760) );
INVx1_ASAP7_75t_L g787 ( .A(n_333), .Y(n_787) );
INVx1_ASAP7_75t_L g417 ( .A(n_336), .Y(n_417) );
INVx1_ASAP7_75t_L g430 ( .A(n_336), .Y(n_430) );
INVx2_ASAP7_75t_L g448 ( .A(n_336), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g1318 ( .A(n_337), .Y(n_1318) );
INVx1_ASAP7_75t_L g979 ( .A(n_338), .Y(n_979) );
CKINVDCx5p33_ASAP7_75t_R g1362 ( .A(n_341), .Y(n_1362) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_370), .B(n_1554), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx4f_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_355), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g1832 ( .A(n_349), .B(n_358), .Y(n_1832) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g1836 ( .A(n_351), .B(n_354), .Y(n_1836) );
INVx1_ASAP7_75t_L g1888 ( .A(n_351), .Y(n_1888) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g1890 ( .A(n_354), .B(n_1888), .Y(n_1890) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_357), .B(n_360), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_L g547 ( .A(n_358), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x4_ASAP7_75t_L g470 ( .A(n_359), .B(n_369), .Y(n_470) );
AND2x4_ASAP7_75t_L g604 ( .A(n_359), .B(n_368), .Y(n_604) );
INVx1_ASAP7_75t_L g1031 ( .A(n_360), .Y(n_1031) );
INVxp67_ASAP7_75t_SL g1500 ( .A(n_360), .Y(n_1500) );
AND2x4_ASAP7_75t_SL g1831 ( .A(n_360), .B(n_1832), .Y(n_1831) );
INVx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x6_ASAP7_75t_L g361 ( .A(n_362), .B(n_367), .Y(n_361) );
BUFx4f_ASAP7_75t_L g439 ( .A(n_362), .Y(n_439) );
OR2x6_ASAP7_75t_L g542 ( .A(n_362), .B(n_516), .Y(n_542) );
INVx1_ASAP7_75t_L g1489 ( .A(n_362), .Y(n_1489) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx3_ASAP7_75t_L g465 ( .A(n_363), .Y(n_465) );
BUFx4f_ASAP7_75t_L g881 ( .A(n_363), .Y(n_881) );
INVx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx2_ASAP7_75t_L g444 ( .A(n_365), .Y(n_444) );
INVx2_ASAP7_75t_L g455 ( .A(n_365), .Y(n_455) );
NAND2x1_ASAP7_75t_L g459 ( .A(n_365), .B(n_366), .Y(n_459) );
AND2x2_ASAP7_75t_L g518 ( .A(n_365), .B(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g529 ( .A(n_365), .B(n_366), .Y(n_529) );
INVx1_ASAP7_75t_L g538 ( .A(n_365), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_366), .B(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g454 ( .A(n_366), .B(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g519 ( .A(n_366), .Y(n_519) );
BUFx2_ASAP7_75t_L g533 ( .A(n_366), .Y(n_533) );
AND2x2_ASAP7_75t_L g557 ( .A(n_366), .B(n_444), .Y(n_557) );
INVx1_ASAP7_75t_L g571 ( .A(n_366), .Y(n_571) );
OR2x6_ASAP7_75t_L g1127 ( .A(n_367), .B(n_465), .Y(n_1127) );
INVxp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g527 ( .A(n_368), .Y(n_527) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g532 ( .A(n_369), .Y(n_532) );
AND2x4_ASAP7_75t_L g536 ( .A(n_369), .B(n_537), .Y(n_536) );
OAI22xp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B1(n_1410), .B2(n_1411), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_1085), .B1(n_1407), .B2(n_1409), .Y(n_372) );
XNOR2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_684), .Y(n_373) );
XNOR2xp5_ASAP7_75t_L g1408 ( .A(n_374), .B(n_684), .Y(n_1408) );
AOI22xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_550), .B1(n_682), .B2(n_683), .Y(n_374) );
INVx1_ASAP7_75t_L g682 ( .A(n_375), .Y(n_682) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND3xp33_ASAP7_75t_L g378 ( .A(n_379), .B(n_473), .C(n_512), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_380), .B(n_437), .Y(n_379) );
OAI33xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_399), .A3(n_412), .B1(n_421), .B2(n_425), .B3(n_432), .Y(n_380) );
OAI22xp33_ASAP7_75t_SL g381 ( .A1(n_382), .A2(n_383), .B1(n_392), .B2(n_393), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_382), .A2(n_434), .B1(n_451), .B2(n_456), .Y(n_450) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g940 ( .A(n_384), .Y(n_940) );
INVx8_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx3_ASAP7_75t_L g433 ( .A(n_385), .Y(n_433) );
INVx5_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_SL g938 ( .A(n_386), .Y(n_938) );
INVx3_ASAP7_75t_L g1335 ( .A(n_386), .Y(n_1335) );
INVx2_ASAP7_75t_SL g1369 ( .A(n_386), .Y(n_1369) );
AOI22xp33_ASAP7_75t_L g1876 ( .A1(n_386), .A2(n_1365), .B1(n_1877), .B2(n_1878), .Y(n_1876) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_387), .Y(n_481) );
BUFx8_ASAP7_75t_L g677 ( .A(n_387), .Y(n_677) );
INVx2_ASAP7_75t_L g705 ( .A(n_387), .Y(n_705) );
AND2x4_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g404 ( .A(n_389), .Y(n_404) );
AND2x4_ASAP7_75t_L g630 ( .A(n_390), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_391), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g403 ( .A(n_391), .B(n_404), .Y(n_403) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_391), .Y(n_411) );
AND2x4_ASAP7_75t_L g488 ( .A(n_391), .B(n_489), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_392), .A2(n_436), .B1(n_464), .B2(n_466), .Y(n_463) );
OAI221xp5_ASAP7_75t_L g758 ( .A1(n_393), .A2(n_759), .B1(n_760), .B2(n_761), .C(n_762), .Y(n_758) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g941 ( .A(n_395), .Y(n_941) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx3_ASAP7_75t_L g435 ( .A(n_396), .Y(n_435) );
OR2x6_ASAP7_75t_L g506 ( .A(n_396), .B(n_428), .Y(n_506) );
BUFx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g615 ( .A(n_397), .Y(n_615) );
INVx1_ASAP7_75t_L g410 ( .A(n_398), .Y(n_410) );
INVx2_ASAP7_75t_L g489 ( .A(n_398), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_405), .B2(n_406), .Y(n_399) );
OAI22xp33_ASAP7_75t_L g438 ( .A1(n_400), .A2(n_422), .B1(n_439), .B2(n_440), .Y(n_438) );
BUFx4f_ASAP7_75t_SL g1009 ( .A(n_401), .Y(n_1009) );
OAI22xp33_ASAP7_75t_L g1105 ( .A1(n_401), .A2(n_1045), .B1(n_1106), .B2(n_1107), .Y(n_1105) );
OAI22xp33_ASAP7_75t_L g1527 ( .A1(n_401), .A2(n_1512), .B1(n_1518), .B2(n_1528), .Y(n_1527) );
OAI22xp33_ASAP7_75t_L g1531 ( .A1(n_401), .A2(n_1096), .B1(n_1513), .B2(n_1520), .Y(n_1531) );
INVx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_SL g671 ( .A(n_402), .Y(n_671) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx3_ASAP7_75t_L g423 ( .A(n_403), .Y(n_423) );
OR2x4_ASAP7_75t_L g477 ( .A(n_403), .B(n_428), .Y(n_477) );
OR2x4_ASAP7_75t_L g503 ( .A(n_403), .B(n_480), .Y(n_503) );
BUFx4f_ASAP7_75t_L g914 ( .A(n_403), .Y(n_914) );
BUFx3_ASAP7_75t_L g1465 ( .A(n_403), .Y(n_1465) );
INVx1_ASAP7_75t_L g631 ( .A(n_404), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_405), .A2(n_424), .B1(n_461), .B2(n_462), .Y(n_460) );
OAI22xp33_ASAP7_75t_L g421 ( .A1(n_406), .A2(n_422), .B1(n_423), .B2(n_424), .Y(n_421) );
OAI22xp33_ASAP7_75t_L g907 ( .A1(n_406), .A2(n_671), .B1(n_878), .B2(n_895), .Y(n_907) );
OAI22xp5_ASAP7_75t_L g1056 ( .A1(n_406), .A2(n_1040), .B1(n_1057), .B2(n_1058), .Y(n_1056) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g1182 ( .A(n_407), .Y(n_1182) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx6f_ASAP7_75t_L g915 ( .A(n_408), .Y(n_915) );
HB1xp67_ASAP7_75t_L g1241 ( .A(n_408), .Y(n_1241) );
HB1xp67_ASAP7_75t_L g1252 ( .A(n_408), .Y(n_1252) );
BUFx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx2_ASAP7_75t_L g485 ( .A(n_409), .Y(n_485) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_409), .Y(n_627) );
NAND2x1p5_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
BUFx2_ASAP7_75t_L g499 ( .A(n_410), .Y(n_499) );
BUFx2_ASAP7_75t_L g495 ( .A(n_411), .Y(n_495) );
AND2x4_ASAP7_75t_L g648 ( .A(n_411), .B(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g662 ( .A(n_411), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_412), .A2(n_798), .B1(n_807), .B2(n_817), .Y(n_797) );
OAI33xp33_ASAP7_75t_L g1037 ( .A1(n_412), .A2(n_1038), .A3(n_1046), .B1(n_1050), .B2(n_1053), .B3(n_1056), .Y(n_1037) );
OAI22xp33_ASAP7_75t_L g1862 ( .A1(n_412), .A2(n_942), .B1(n_1863), .B2(n_1868), .Y(n_1862) );
BUFx3_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx4f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx4f_ASAP7_75t_L g767 ( .A(n_414), .Y(n_767) );
BUFx2_ASAP7_75t_L g1092 ( .A(n_414), .Y(n_1092) );
BUFx8_ASAP7_75t_L g1237 ( .A(n_414), .Y(n_1237) );
OR2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_418), .Y(n_414) );
INVx1_ASAP7_75t_L g472 ( .A(n_415), .Y(n_472) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_415), .Y(n_511) );
OR2x2_ASAP7_75t_L g616 ( .A(n_415), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_SL g1116 ( .A(n_415), .B(n_470), .Y(n_1116) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx2_ASAP7_75t_L g549 ( .A(n_416), .Y(n_549) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx2_ASAP7_75t_L g1352 ( .A(n_418), .Y(n_1352) );
NAND2xp33_ASAP7_75t_SL g418 ( .A(n_419), .B(n_420), .Y(n_418) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_419), .Y(n_509) );
INVx1_ASAP7_75t_L g633 ( .A(n_419), .Y(n_633) );
AND3x4_ASAP7_75t_L g638 ( .A(n_419), .B(n_494), .C(n_609), .Y(n_638) );
INVx3_ASAP7_75t_L g428 ( .A(n_420), .Y(n_428) );
BUFx3_ASAP7_75t_L g494 ( .A(n_420), .Y(n_494) );
OAI22xp33_ASAP7_75t_L g1155 ( .A1(n_423), .A2(n_1156), .B1(n_1157), .B2(n_1158), .Y(n_1155) );
OAI22xp33_ASAP7_75t_L g1190 ( .A1(n_423), .A2(n_1191), .B1(n_1192), .B2(n_1193), .Y(n_1190) );
OAI22xp33_ASAP7_75t_L g1238 ( .A1(n_423), .A2(n_1239), .B1(n_1240), .B2(n_1241), .Y(n_1238) );
OAI22xp33_ASAP7_75t_L g1249 ( .A1(n_423), .A2(n_1250), .B1(n_1251), .B2(n_1252), .Y(n_1249) );
OAI221xp5_ASAP7_75t_L g1343 ( .A1(n_423), .A2(n_1132), .B1(n_1297), .B2(n_1305), .C(n_1344), .Y(n_1343) );
OAI33xp33_ASAP7_75t_L g1189 ( .A1(n_425), .A2(n_767), .A3(n_1190), .B1(n_1194), .B2(n_1197), .B3(n_1202), .Y(n_1189) );
OAI33xp33_ASAP7_75t_L g1236 ( .A1(n_425), .A2(n_1237), .A3(n_1238), .B1(n_1242), .B2(n_1245), .B3(n_1249), .Y(n_1236) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_426), .Y(n_425) );
NAND3xp33_ASAP7_75t_L g768 ( .A(n_426), .B(n_769), .C(n_772), .Y(n_768) );
INVx2_ASAP7_75t_L g817 ( .A(n_426), .Y(n_817) );
INVx2_ASAP7_75t_L g942 ( .A(n_426), .Y(n_942) );
AOI221xp5_ASAP7_75t_L g1004 ( .A1(n_426), .A2(n_680), .B1(n_1005), .B2(n_1012), .C(n_1019), .Y(n_1004) );
INVx3_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx3_ASAP7_75t_L g1055 ( .A(n_427), .Y(n_1055) );
NAND3x1_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .C(n_431), .Y(n_427) );
INVx1_ASAP7_75t_L g480 ( .A(n_428), .Y(n_480) );
AND2x4_ASAP7_75t_L g487 ( .A(n_428), .B(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g632 ( .A(n_428), .B(n_633), .Y(n_632) );
NAND2x1p5_ASAP7_75t_L g654 ( .A(n_428), .B(n_431), .Y(n_654) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g619 ( .A(n_430), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_430), .B(n_558), .Y(n_1286) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B1(n_435), .B2(n_436), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g1242 ( .A1(n_433), .A2(n_801), .B1(n_1243), .B2(n_1244), .Y(n_1242) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_435), .A2(n_887), .B1(n_902), .B2(n_909), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_435), .A2(n_926), .B1(n_933), .B2(n_938), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g1245 ( .A1(n_435), .A2(n_1246), .B1(n_1247), .B2(n_1248), .Y(n_1245) );
OAI22xp5_ASAP7_75t_L g1467 ( .A1(n_435), .A2(n_940), .B1(n_1468), .B2(n_1469), .Y(n_1467) );
OAI33xp33_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_445), .A3(n_450), .B1(n_460), .B2(n_463), .B3(n_468), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g1117 ( .A1(n_439), .A2(n_598), .B1(n_1100), .B2(n_1104), .Y(n_1117) );
OAI22xp5_ASAP7_75t_L g1164 ( .A1(n_439), .A2(n_598), .B1(n_1149), .B2(n_1154), .Y(n_1164) );
OAI22xp33_ASAP7_75t_L g1511 ( .A1(n_439), .A2(n_1295), .B1(n_1512), .B2(n_1513), .Y(n_1511) );
OAI22xp33_ASAP7_75t_L g1254 ( .A1(n_440), .A2(n_1239), .B1(n_1250), .B2(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_441), .Y(n_467) );
INVx2_ASAP7_75t_SL g885 ( .A(n_441), .Y(n_885) );
INVx1_ASAP7_75t_L g904 ( .A(n_441), .Y(n_904) );
INVx4_ASAP7_75t_L g1066 ( .A(n_441), .Y(n_1066) );
INVx2_ASAP7_75t_L g1296 ( .A(n_441), .Y(n_1296) );
INVx2_ASAP7_75t_L g1444 ( .A(n_441), .Y(n_1444) );
INVx2_ASAP7_75t_L g1525 ( .A(n_441), .Y(n_1525) );
INVx8_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g545 ( .A(n_442), .B(n_532), .Y(n_545) );
BUFx2_ASAP7_75t_L g598 ( .A(n_442), .Y(n_598) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI33xp33_ASAP7_75t_L g876 ( .A1(n_445), .A2(n_877), .A3(n_886), .B1(n_891), .B2(n_898), .B3(n_901), .Y(n_876) );
OAI33xp33_ASAP7_75t_L g1059 ( .A1(n_445), .A2(n_898), .A3(n_1060), .B1(n_1067), .B2(n_1070), .B3(n_1071), .Y(n_1059) );
INVx1_ASAP7_75t_L g1298 ( .A(n_445), .Y(n_1298) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx4_ASAP7_75t_L g921 ( .A(n_446), .Y(n_921) );
INVx2_ASAP7_75t_L g1161 ( .A(n_446), .Y(n_1161) );
INVx2_ASAP7_75t_L g1207 ( .A(n_446), .Y(n_1207) );
INVx1_ASAP7_75t_L g1478 ( .A(n_446), .Y(n_1478) );
AND2x4_ASAP7_75t_L g446 ( .A(n_447), .B(n_449), .Y(n_446) );
OR2x6_ASAP7_75t_L g653 ( .A(n_447), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g756 ( .A(n_447), .Y(n_756) );
BUFx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g609 ( .A(n_448), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_448), .B(n_575), .Y(n_1311) );
OAI22xp5_ASAP7_75t_L g1165 ( .A1(n_451), .A2(n_896), .B1(n_1145), .B2(n_1157), .Y(n_1165) );
OAI22xp5_ASAP7_75t_L g1514 ( .A1(n_451), .A2(n_456), .B1(n_1515), .B2(n_1516), .Y(n_1514) );
INVx4_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g461 ( .A(n_452), .Y(n_461) );
INVx2_ASAP7_75t_L g888 ( .A(n_452), .Y(n_888) );
INVx2_ASAP7_75t_L g1519 ( .A(n_452), .Y(n_1519) );
INVx4_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx3_ASAP7_75t_L g894 ( .A(n_454), .Y(n_894) );
INVx2_ASAP7_75t_L g1069 ( .A(n_454), .Y(n_1069) );
BUFx2_ASAP7_75t_L g1113 ( .A(n_454), .Y(n_1113) );
INVx1_ASAP7_75t_L g1303 ( .A(n_454), .Y(n_1303) );
AND2x2_ASAP7_75t_L g570 ( .A(n_455), .B(n_571), .Y(n_570) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_455), .Y(n_735) );
OAI211xp5_ASAP7_75t_L g743 ( .A1(n_456), .A2(n_744), .B(n_745), .C(n_748), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_456), .A2(n_892), .B1(n_930), .B2(n_931), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g1209 ( .A1(n_456), .A2(n_1195), .B1(n_1198), .B2(n_1210), .Y(n_1209) );
OAI22xp5_ASAP7_75t_L g1256 ( .A1(n_456), .A2(n_1210), .B1(n_1243), .B2(n_1246), .Y(n_1256) );
OAI22xp5_ASAP7_75t_L g1480 ( .A1(n_456), .A2(n_1468), .B1(n_1471), .B2(n_1481), .Y(n_1480) );
OAI22xp33_ASAP7_75t_L g1483 ( .A1(n_456), .A2(n_1466), .B1(n_1476), .B2(n_1484), .Y(n_1483) );
INVx5_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_SL g462 ( .A(n_458), .Y(n_462) );
BUFx3_ASAP7_75t_L g827 ( .A(n_458), .Y(n_827) );
OR2x2_ASAP7_75t_L g1287 ( .A(n_458), .B(n_1286), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1393 ( .A(n_458), .B(n_1394), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1446 ( .A(n_458), .B(n_1447), .Y(n_1446) );
BUFx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_459), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_461), .A2(n_462), .B1(n_1240), .B2(n_1251), .Y(n_1257) );
OAI22xp5_ASAP7_75t_L g1212 ( .A1(n_462), .A2(n_1192), .B1(n_1204), .B2(n_1210), .Y(n_1212) );
BUFx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_SL g596 ( .A(n_465), .Y(n_596) );
BUFx6f_ASAP7_75t_L g1163 ( .A(n_465), .Y(n_1163) );
BUFx3_ASAP7_75t_L g1294 ( .A(n_465), .Y(n_1294) );
OAI22xp5_ASAP7_75t_L g1208 ( .A1(n_466), .A2(n_1061), .B1(n_1191), .B2(n_1203), .Y(n_1208) );
OAI22xp5_ASAP7_75t_L g1213 ( .A1(n_466), .A2(n_1063), .B1(n_1196), .B2(n_1200), .Y(n_1213) );
OAI22xp5_ASAP7_75t_L g1258 ( .A1(n_466), .A2(n_1244), .B1(n_1248), .B2(n_1259), .Y(n_1258) );
OAI22xp33_ASAP7_75t_L g1479 ( .A1(n_466), .A2(n_1259), .B1(n_1462), .B2(n_1475), .Y(n_1479) );
INVx6_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OAI33xp33_ASAP7_75t_L g1205 ( .A1(n_468), .A2(n_1206), .A3(n_1208), .B1(n_1209), .B2(n_1212), .B3(n_1213), .Y(n_1205) );
OAI33xp33_ASAP7_75t_L g1253 ( .A1(n_468), .A2(n_1206), .A3(n_1254), .B1(n_1256), .B2(n_1257), .B3(n_1258), .Y(n_1253) );
OAI33xp33_ASAP7_75t_L g1477 ( .A1(n_468), .A2(n_1478), .A3(n_1479), .B1(n_1480), .B2(n_1483), .B3(n_1485), .Y(n_1477) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g1307 ( .A(n_469), .Y(n_1307) );
AND2x4_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx1_ASAP7_75t_SL g566 ( .A(n_470), .Y(n_566) );
INVx4_ASAP7_75t_L g747 ( .A(n_470), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_470), .B(n_471), .Y(n_900) );
OAI21xp33_ASAP7_75t_L g1397 ( .A1(n_470), .A2(n_894), .B(n_1398), .Y(n_1397) );
OAI221xp5_ASAP7_75t_L g1450 ( .A1(n_470), .A2(n_524), .B1(n_894), .B2(n_1451), .C(n_1452), .Y(n_1450) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OAI31xp33_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_482), .A3(n_501), .B(n_507), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_SL g793 ( .A(n_477), .Y(n_793) );
INVx2_ASAP7_75t_SL g1075 ( .A(n_477), .Y(n_1075) );
HB1xp67_ASAP7_75t_L g1225 ( .A(n_477), .Y(n_1225) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_479), .A2(n_783), .B1(n_784), .B2(n_785), .Y(n_782) );
INVx1_ASAP7_75t_L g872 ( .A(n_479), .Y(n_872) );
INVx2_ASAP7_75t_L g1076 ( .A(n_479), .Y(n_1076) );
INVx1_ASAP7_75t_L g1179 ( .A(n_479), .Y(n_1179) );
INVx1_ASAP7_75t_L g1226 ( .A(n_479), .Y(n_1226) );
INVxp67_ASAP7_75t_L g1535 ( .A(n_479), .Y(n_1535) );
AND2x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_481), .Y(n_645) );
INVx2_ASAP7_75t_L g759 ( .A(n_481), .Y(n_759) );
INVx1_ASAP7_75t_L g1199 ( .A(n_481), .Y(n_1199) );
BUFx6f_ASAP7_75t_L g1347 ( .A(n_481), .Y(n_1347) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVxp67_ASAP7_75t_SL g949 ( .A(n_484), .Y(n_949) );
INVxp67_ASAP7_75t_SL g1158 ( .A(n_484), .Y(n_1158) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g1097 ( .A(n_485), .Y(n_1097) );
NAND4xp25_ASAP7_75t_L g781 ( .A(n_486), .B(n_782), .C(n_786), .D(n_791), .Y(n_781) );
CKINVDCx8_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
CKINVDCx8_ASAP7_75t_R g867 ( .A(n_487), .Y(n_867) );
OAI31xp33_ASAP7_75t_L g1872 ( .A1(n_487), .A2(n_1873), .A3(n_1882), .B(n_1883), .Y(n_1872) );
BUFx2_ASAP7_75t_L g643 ( .A(n_488), .Y(n_643) );
INVx2_ASAP7_75t_L g657 ( .A(n_488), .Y(n_657) );
BUFx2_ASAP7_75t_L g681 ( .A(n_488), .Y(n_681) );
BUFx2_ASAP7_75t_L g766 ( .A(n_488), .Y(n_766) );
BUFx2_ASAP7_75t_L g790 ( .A(n_488), .Y(n_790) );
BUFx3_ASAP7_75t_L g1328 ( .A(n_488), .Y(n_1328) );
BUFx2_ASAP7_75t_L g1807 ( .A(n_488), .Y(n_1807) );
INVx1_ASAP7_75t_L g649 ( .A(n_489), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_496), .B1(n_497), .B2(n_500), .Y(n_490) );
AOI222xp33_ASAP7_75t_L g786 ( .A1(n_491), .A2(n_497), .B1(n_787), .B2(n_788), .C1(n_789), .C2(n_790), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g1270 ( .A1(n_491), .A2(n_497), .B1(n_1264), .B2(n_1271), .Y(n_1270) );
BUFx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx3_ASAP7_75t_L g1079 ( .A(n_492), .Y(n_1079) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_495), .Y(n_492) );
AND2x4_ASAP7_75t_L g498 ( .A(n_493), .B(n_499), .Y(n_498) );
AND2x4_ASAP7_75t_L g869 ( .A(n_493), .B(n_495), .Y(n_869) );
A2O1A1Ixp33_ASAP7_75t_L g1873 ( .A1(n_493), .A2(n_1874), .B(n_1876), .C(n_1879), .Y(n_1873) );
INVx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_496), .A2(n_531), .B1(n_534), .B2(n_539), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_497), .A2(n_1028), .B1(n_1079), .B2(n_1080), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g1228 ( .A1(n_497), .A2(n_1079), .B1(n_1218), .B2(n_1229), .Y(n_1228) );
AOI22xp33_ASAP7_75t_L g1494 ( .A1(n_497), .A2(n_1079), .B1(n_1495), .B2(n_1496), .Y(n_1494) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_498), .A2(n_849), .B1(n_869), .B2(n_870), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_498), .A2(n_869), .B1(n_951), .B2(n_952), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_498), .A2(n_869), .B1(n_1121), .B2(n_1134), .Y(n_1133) );
AOI22xp33_ASAP7_75t_SL g1183 ( .A1(n_498), .A2(n_869), .B1(n_1173), .B2(n_1184), .Y(n_1183) );
AOI22xp33_ASAP7_75t_L g1537 ( .A1(n_498), .A2(n_869), .B1(n_1538), .B2(n_1539), .Y(n_1537) );
AOI22xp5_ASAP7_75t_L g1879 ( .A1(n_498), .A2(n_869), .B1(n_1880), .B2(n_1881), .Y(n_1879) );
BUFx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_SL g795 ( .A(n_503), .Y(n_795) );
BUFx2_ASAP7_75t_L g863 ( .A(n_503), .Y(n_863) );
BUFx3_ASAP7_75t_L g1541 ( .A(n_503), .Y(n_1541) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g785 ( .A(n_506), .Y(n_785) );
BUFx3_ASAP7_75t_L g873 ( .A(n_506), .Y(n_873) );
INVx1_ASAP7_75t_L g1232 ( .A(n_506), .Y(n_1232) );
OAI31xp33_ASAP7_75t_L g1490 ( .A1(n_507), .A2(n_1491), .A3(n_1492), .B(n_1497), .Y(n_1490) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_510), .Y(n_507) );
AND2x4_ASAP7_75t_L g796 ( .A(n_508), .B(n_510), .Y(n_796) );
AND2x2_ASAP7_75t_SL g874 ( .A(n_508), .B(n_510), .Y(n_874) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_508), .B(n_510), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1883 ( .A(n_508), .B(n_510), .Y(n_1883) );
INVx1_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
OAI31xp33_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_520), .A3(n_540), .B(n_546), .Y(n_512) );
CKINVDCx16_ASAP7_75t_R g514 ( .A(n_515), .Y(n_514) );
INVx4_ASAP7_75t_L g859 ( .A(n_515), .Y(n_859) );
INVx3_ASAP7_75t_SL g1032 ( .A(n_515), .Y(n_1032) );
AND2x4_ASAP7_75t_L g515 ( .A(n_516), .B(n_518), .Y(n_515) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g565 ( .A(n_518), .Y(n_565) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_518), .Y(n_583) );
BUFx3_ASAP7_75t_L g994 ( .A(n_518), .Y(n_994) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g1160 ( .A1(n_523), .A2(n_1113), .B1(n_1148), .B2(n_1152), .Y(n_1160) );
OAI22xp5_ASAP7_75t_L g1517 ( .A1(n_523), .A2(n_1518), .B1(n_1519), .B2(n_1520), .Y(n_1517) );
BUFx4f_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx4_ASAP7_75t_L g846 ( .A(n_524), .Y(n_846) );
BUFx4f_ASAP7_75t_L g890 ( .A(n_524), .Y(n_890) );
BUFx4f_ASAP7_75t_L g928 ( .A(n_524), .Y(n_928) );
BUFx4f_ASAP7_75t_L g1304 ( .A(n_524), .Y(n_1304) );
OR2x6_ASAP7_75t_L g1308 ( .A(n_524), .B(n_1309), .Y(n_1308) );
BUFx6f_ASAP7_75t_L g1861 ( .A(n_524), .Y(n_1861) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx3_ASAP7_75t_L g847 ( .A(n_526), .Y(n_847) );
INVx1_ASAP7_75t_L g1026 ( .A(n_526), .Y(n_1026) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_527), .B(n_1171), .Y(n_1170) );
BUFx3_ASAP7_75t_L g561 ( .A(n_528), .Y(n_561) );
AND2x6_ASAP7_75t_L g574 ( .A(n_528), .B(n_575), .Y(n_574) );
AND2x4_ASAP7_75t_SL g588 ( .A(n_528), .B(n_558), .Y(n_588) );
INVx1_ASAP7_75t_L g602 ( .A(n_528), .Y(n_602) );
BUFx6f_ASAP7_75t_L g725 ( .A(n_528), .Y(n_725) );
BUFx3_ASAP7_75t_L g1396 ( .A(n_528), .Y(n_1396) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g740 ( .A(n_529), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_531), .A2(n_1121), .B1(n_1122), .B2(n_1124), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_531), .A2(n_1122), .B1(n_1173), .B2(n_1174), .Y(n_1172) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_531), .A2(n_1218), .B1(n_1219), .B2(n_1220), .Y(n_1217) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
AND2x4_ASAP7_75t_L g851 ( .A(n_532), .B(n_533), .Y(n_851) );
INVx1_ASAP7_75t_L g592 ( .A(n_533), .Y(n_592) );
BUFx2_ASAP7_75t_L g989 ( .A(n_533), .Y(n_989) );
INVx1_ASAP7_75t_L g1315 ( .A(n_533), .Y(n_1315) );
AOI22xp33_ASAP7_75t_L g1394 ( .A1(n_533), .A2(n_734), .B1(n_1358), .B2(n_1375), .Y(n_1394) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_534), .A2(n_849), .B1(n_850), .B2(n_852), .Y(n_848) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx3_ASAP7_75t_L g959 ( .A(n_536), .Y(n_959) );
INVx2_ASAP7_75t_L g1123 ( .A(n_536), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1263 ( .A1(n_536), .A2(n_851), .B1(n_1264), .B2(n_1265), .Y(n_1263) );
AOI22xp33_ASAP7_75t_L g1548 ( .A1(n_536), .A2(n_851), .B1(n_1538), .B2(n_1549), .Y(n_1548) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_537), .B(n_575), .Y(n_625) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g855 ( .A(n_542), .Y(n_855) );
HB1xp67_ASAP7_75t_L g1034 ( .A(n_542), .Y(n_1034) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g1035 ( .A(n_544), .Y(n_1035) );
INVx2_ASAP7_75t_L g1222 ( .A(n_544), .Y(n_1222) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g857 ( .A(n_545), .Y(n_857) );
BUFx2_ASAP7_75t_L g962 ( .A(n_545), .Y(n_962) );
OAI31xp33_ASAP7_75t_L g843 ( .A1(n_546), .A2(n_844), .A3(n_853), .B(n_858), .Y(n_843) );
OAI31xp33_ASAP7_75t_L g1214 ( .A1(n_546), .A2(n_1215), .A3(n_1216), .B(n_1221), .Y(n_1214) );
BUFx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx2_ASAP7_75t_SL g964 ( .A(n_547), .Y(n_964) );
OAI31xp33_ASAP7_75t_L g1024 ( .A1(n_547), .A2(n_1025), .A3(n_1030), .B(n_1033), .Y(n_1024) );
OAI31xp33_ASAP7_75t_L g1118 ( .A1(n_547), .A2(n_1119), .A3(n_1125), .B(n_1126), .Y(n_1118) );
BUFx2_ASAP7_75t_L g1176 ( .A(n_547), .Y(n_1176) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g624 ( .A(n_549), .B(n_625), .Y(n_624) );
INVxp67_ASAP7_75t_L g634 ( .A(n_549), .Y(n_634) );
INVx1_ASAP7_75t_L g698 ( .A(n_549), .Y(n_698) );
INVx1_ASAP7_75t_L g683 ( .A(n_550), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_610), .C(n_635), .Y(n_551) );
OAI21xp33_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_584), .B(n_605), .Y(n_552) );
INVx2_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
INVx1_ASAP7_75t_L g1437 ( .A(n_556), .Y(n_1437) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g573 ( .A(n_557), .Y(n_573) );
BUFx3_ASAP7_75t_L g729 ( .A(n_557), .Y(n_729) );
BUFx3_ASAP7_75t_L g750 ( .A(n_557), .Y(n_750) );
AND2x2_ASAP7_75t_L g579 ( .A(n_558), .B(n_570), .Y(n_579) );
AND2x4_ASAP7_75t_L g582 ( .A(n_558), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g708 ( .A(n_558), .B(n_583), .Y(n_708) );
AND2x2_ASAP7_75t_L g752 ( .A(n_558), .B(n_572), .Y(n_752) );
BUFx2_ASAP7_75t_L g1387 ( .A(n_558), .Y(n_1387) );
AOI21xp5_ASAP7_75t_SL g559 ( .A1(n_560), .A2(n_567), .B(n_574), .Y(n_559) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g1290 ( .A(n_563), .Y(n_1290) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g829 ( .A(n_565), .Y(n_829) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g728 ( .A(n_569), .Y(n_728) );
INVx2_ASAP7_75t_SL g732 ( .A(n_569), .Y(n_732) );
INVx1_ASAP7_75t_L g749 ( .A(n_569), .Y(n_749) );
INVx2_ASAP7_75t_L g1795 ( .A(n_569), .Y(n_1795) );
INVx3_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_570), .B(n_575), .Y(n_620) );
BUFx6f_ASAP7_75t_L g831 ( .A(n_570), .Y(n_831) );
AND2x4_ASAP7_75t_L g1284 ( .A(n_572), .B(n_1285), .Y(n_1284) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g1855 ( .A(n_573), .Y(n_1855) );
AOI211xp5_ASAP7_75t_SL g835 ( .A1(n_574), .A2(n_754), .B(n_788), .C(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g593 ( .A(n_575), .Y(n_593) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_575), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B1(n_580), .B2(n_581), .Y(n_576) );
INVx1_ASAP7_75t_L g821 ( .A(n_578), .Y(n_821) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x4_ASAP7_75t_L g697 ( .A(n_579), .B(n_698), .Y(n_697) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g824 ( .A(n_582), .Y(n_824) );
INVx1_ASAP7_75t_L g724 ( .A(n_583), .Y(n_724) );
BUFx6f_ASAP7_75t_L g746 ( .A(n_583), .Y(n_746) );
INVx2_ASAP7_75t_L g1390 ( .A(n_583), .Y(n_1390) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g1002 ( .A(n_586), .Y(n_1002) );
INVx4_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
BUFx3_ASAP7_75t_L g754 ( .A(n_588), .Y(n_754) );
BUFx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2x1_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_L g736 ( .A(n_592), .Y(n_736) );
INVx1_ASAP7_75t_L g1448 ( .A(n_593), .Y(n_1448) );
OAI221xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_597), .B1(n_598), .B2(n_599), .C(n_600), .Y(n_594) );
OAI22xp33_ASAP7_75t_L g1111 ( .A1(n_595), .A2(n_1066), .B1(n_1094), .B2(n_1106), .Y(n_1111) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx3_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g726 ( .A(n_604), .Y(n_726) );
OAI221xp5_ASAP7_75t_L g1381 ( .A1(n_604), .A2(n_998), .B1(n_1382), .B2(n_1383), .C(n_1384), .Y(n_1381) );
OAI221xp5_ASAP7_75t_L g1438 ( .A1(n_604), .A2(n_998), .B1(n_1068), .B2(n_1439), .C(n_1440), .Y(n_1438) );
INVx1_ASAP7_75t_L g1853 ( .A(n_604), .Y(n_1853) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AOI21xp33_ASAP7_75t_L g818 ( .A1(n_606), .A2(n_819), .B(n_835), .Y(n_818) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
HB1xp67_ASAP7_75t_L g1003 ( .A(n_607), .Y(n_1003) );
BUFx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OAI31xp33_ASAP7_75t_L g1377 ( .A1(n_608), .A2(n_1378), .A3(n_1385), .B(n_1395), .Y(n_1377) );
OAI31xp33_ASAP7_75t_L g1434 ( .A1(n_608), .A2(n_1435), .A3(n_1441), .B(n_1449), .Y(n_1434) );
AOI21x1_ASAP7_75t_L g1789 ( .A1(n_608), .A2(n_1790), .B(n_1803), .Y(n_1789) );
HB1xp67_ASAP7_75t_L g1841 ( .A(n_608), .Y(n_1841) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AOI21xp33_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_621), .B(n_622), .Y(n_610) );
INVx8_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x4_ASAP7_75t_L g612 ( .A(n_613), .B(n_618), .Y(n_612) );
INVx1_ASAP7_75t_L g717 ( .A(n_613), .Y(n_717) );
OR2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
BUFx3_ASAP7_75t_L g1103 ( .A(n_614), .Y(n_1103) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
BUFx6f_ASAP7_75t_L g802 ( .A(n_615), .Y(n_802) );
OR2x2_ASAP7_75t_L g626 ( .A(n_616), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g673 ( .A(n_616), .Y(n_673) );
INVx1_ASAP7_75t_L g676 ( .A(n_616), .Y(n_676) );
INVx1_ASAP7_75t_L g1341 ( .A(n_617), .Y(n_1341) );
INVx1_ASAP7_75t_L g1282 ( .A(n_618), .Y(n_1282) );
OR2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
AND2x4_ASAP7_75t_L g663 ( .A(n_619), .B(n_632), .Y(n_663) );
AND2x4_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
INVx1_ASAP7_75t_L g838 ( .A(n_625), .Y(n_838) );
INVx2_ASAP7_75t_L g719 ( .A(n_626), .Y(n_719) );
INVx3_ASAP7_75t_L g866 ( .A(n_627), .Y(n_866) );
INVx4_ASAP7_75t_L g1011 ( .A(n_627), .Y(n_1011) );
BUFx6f_ASAP7_75t_L g1045 ( .A(n_627), .Y(n_1045) );
INVx3_ASAP7_75t_L g692 ( .A(n_628), .Y(n_692) );
INVx5_ASAP7_75t_L g1405 ( .A(n_628), .Y(n_1405) );
OR2x6_ASAP7_75t_L g628 ( .A(n_629), .B(n_634), .Y(n_628) );
NAND2x1p5_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
BUFx3_ASAP7_75t_L g642 ( .A(n_630), .Y(n_642) );
BUFx3_ASAP7_75t_L g765 ( .A(n_630), .Y(n_765) );
INVx8_ASAP7_75t_L g774 ( .A(n_630), .Y(n_774) );
HB1xp67_ASAP7_75t_L g1333 ( .A(n_630), .Y(n_1333) );
AND2x6_ASAP7_75t_L g1322 ( .A(n_632), .B(n_661), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_632), .B(n_668), .Y(n_1324) );
INVx1_ASAP7_75t_L g1330 ( .A(n_632), .Y(n_1330) );
NOR3xp33_ASAP7_75t_L g635 ( .A(n_636), .B(n_669), .C(n_678), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_637), .B(n_658), .Y(n_636) );
AOI33xp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .A3(n_644), .B1(n_650), .B2(n_652), .B3(n_655), .Y(n_637) );
BUFx3_ASAP7_75t_L g1019 ( .A(n_638), .Y(n_1019) );
AOI33xp33_ASAP7_75t_L g1363 ( .A1(n_638), .A2(n_652), .A3(n_1364), .B1(n_1366), .B2(n_1367), .B3(n_1370), .Y(n_1363) );
NAND3xp33_ASAP7_75t_L g1416 ( .A(n_638), .B(n_1417), .C(n_1418), .Y(n_1416) );
AOI33xp33_ASAP7_75t_L g1805 ( .A1(n_638), .A2(n_1806), .A3(n_1808), .B1(n_1809), .B2(n_1810), .B3(n_1812), .Y(n_1805) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
BUFx3_ASAP7_75t_L g805 ( .A(n_642), .Y(n_805) );
INVx1_ASAP7_75t_L g814 ( .A(n_642), .Y(n_814) );
INVx1_ASAP7_75t_L g1530 ( .A(n_645), .Y(n_1530) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx5_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
BUFx3_ASAP7_75t_L g651 ( .A(n_648), .Y(n_651) );
BUFx12f_ASAP7_75t_L g771 ( .A(n_648), .Y(n_771) );
BUFx3_ASAP7_75t_L g1006 ( .A(n_648), .Y(n_1006) );
INVx1_ASAP7_75t_L g668 ( .A(n_649), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g1425 ( .A(n_652), .B(n_1426), .C(n_1427), .Y(n_1425) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI33xp33_ASAP7_75t_L g1091 ( .A1(n_653), .A2(n_1092), .A3(n_1093), .B1(n_1098), .B2(n_1101), .B3(n_1105), .Y(n_1091) );
OAI33xp33_ASAP7_75t_L g1142 ( .A1(n_653), .A2(n_1092), .A3(n_1143), .B1(n_1147), .B2(n_1151), .B3(n_1155), .Y(n_1142) );
OAI33xp33_ASAP7_75t_L g1526 ( .A1(n_653), .A2(n_1237), .A3(n_1527), .B1(n_1529), .B2(n_1531), .B3(n_1532), .Y(n_1526) );
INVx1_ASAP7_75t_L g1812 ( .A(n_653), .Y(n_1812) );
INVx3_ASAP7_75t_L g1344 ( .A(n_654), .Y(n_1344) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g775 ( .A(n_657), .Y(n_775) );
INVx1_ASAP7_75t_L g806 ( .A(n_657), .Y(n_806) );
INVx2_ASAP7_75t_L g1811 ( .A(n_657), .Y(n_1811) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B1(n_664), .B2(n_665), .Y(n_658) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
AND2x4_ASAP7_75t_SL g712 ( .A(n_661), .B(n_663), .Y(n_712) );
NAND2x1_ASAP7_75t_L g977 ( .A(n_661), .B(n_663), .Y(n_977) );
INVx3_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x4_ASAP7_75t_L g665 ( .A(n_663), .B(n_666), .Y(n_665) );
AND2x4_ASAP7_75t_L g680 ( .A(n_663), .B(n_681), .Y(n_680) );
AND2x4_ASAP7_75t_SL g714 ( .A(n_663), .B(n_666), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g975 ( .A1(n_665), .A2(n_976), .B1(n_978), .B2(n_979), .C(n_980), .Y(n_975) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
OR2x6_ASAP7_75t_L g699 ( .A(n_671), .B(n_672), .Y(n_699) );
OAI22xp33_ASAP7_75t_L g936 ( .A1(n_671), .A2(n_915), .B1(n_923), .B2(n_930), .Y(n_936) );
OAI22xp33_ASAP7_75t_L g943 ( .A1(n_671), .A2(n_865), .B1(n_924), .B2(n_931), .Y(n_943) );
INVx2_ASAP7_75t_SL g1041 ( .A(n_671), .Y(n_1041) );
INVxp67_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g703 ( .A(n_673), .B(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g1371 ( .A(n_675), .B(n_1372), .Y(n_1371) );
NAND2xp5_ASAP7_75t_L g1419 ( .A(n_675), .B(n_1420), .Y(n_1419) );
AND2x4_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
AND2x4_ASAP7_75t_L g1359 ( .A(n_676), .B(n_1360), .Y(n_1359) );
INVx3_ASAP7_75t_L g909 ( .A(n_677), .Y(n_909) );
INVx3_ASAP7_75t_L g911 ( .A(n_677), .Y(n_911) );
INVx2_ASAP7_75t_SL g1014 ( .A(n_677), .Y(n_1014) );
INVx2_ASAP7_75t_SL g1153 ( .A(n_677), .Y(n_1153) );
INVx2_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
OAI211xp5_ASAP7_75t_SL g757 ( .A1(n_679), .A2(n_758), .B(n_767), .C(n_768), .Y(n_757) );
INVx3_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g1374 ( .A1(n_680), .A2(n_712), .B1(n_714), .B2(n_1375), .C(n_1376), .Y(n_1374) );
AOI221xp5_ASAP7_75t_L g1429 ( .A1(n_680), .A2(n_712), .B1(n_714), .B2(n_1430), .C(n_1431), .Y(n_1429) );
AOI221xp5_ASAP7_75t_L g1813 ( .A1(n_680), .A2(n_712), .B1(n_714), .B2(n_1800), .C(n_1814), .Y(n_1813) );
XOR2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_967), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .B1(n_840), .B2(n_966), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
XOR2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_778), .Y(n_687) );
INVx1_ASAP7_75t_L g776 ( .A(n_689), .Y(n_776) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_693), .C(n_709), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_691), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B1(n_700), .B2(n_701), .Y(n_693) );
INVxp67_ASAP7_75t_L g972 ( .A(n_695), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_696), .B(n_699), .Y(n_695) );
INVx3_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g1316 ( .A1(n_697), .A2(n_707), .B1(n_1317), .B2(n_1318), .Y(n_1316) );
AND2x4_ASAP7_75t_L g707 ( .A(n_698), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g973 ( .A(n_701), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g1815 ( .A(n_701), .B(n_1816), .Y(n_1815) );
NAND2x1_ASAP7_75t_L g701 ( .A(n_702), .B(n_706), .Y(n_701) );
INVx2_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g1869 ( .A(n_704), .Y(n_1869) );
INVx3_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g770 ( .A(n_705), .Y(n_770) );
BUFx2_ASAP7_75t_L g808 ( .A(n_705), .Y(n_808) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NOR3xp33_ASAP7_75t_SL g709 ( .A(n_710), .B(n_720), .C(n_757), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B1(n_718), .B2(n_719), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_716), .B(n_732), .Y(n_731) );
AOI222xp33_ASAP7_75t_L g1357 ( .A1(n_717), .A2(n_719), .B1(n_1358), .B2(n_1359), .C1(n_1361), .C2(n_1362), .Y(n_1357) );
AOI222xp33_ASAP7_75t_L g1421 ( .A1(n_717), .A2(n_719), .B1(n_1359), .B2(n_1422), .C1(n_1423), .C2(n_1424), .Y(n_1421) );
AOI222xp33_ASAP7_75t_L g1817 ( .A1(n_717), .A2(n_719), .B1(n_1359), .B2(n_1801), .C1(n_1818), .C2(n_1819), .Y(n_1817) );
AOI221xp5_ASAP7_75t_L g733 ( .A1(n_718), .A2(n_734), .B1(n_736), .B2(n_737), .C(n_738), .Y(n_733) );
AOI31xp33_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_743), .A3(n_751), .B(n_755), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_727), .B(n_730), .Y(n_721) );
INVx2_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
BUFx2_ASAP7_75t_L g1291 ( .A(n_725), .Y(n_1291) );
AOI221xp5_ASAP7_75t_L g1388 ( .A1(n_725), .A2(n_1372), .B1(n_1376), .B2(n_1389), .C(n_1391), .Y(n_1388) );
AOI221xp5_ASAP7_75t_L g1442 ( .A1(n_725), .A2(n_1389), .B1(n_1420), .B2(n_1431), .C(n_1443), .Y(n_1442) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_733), .B(n_741), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_734), .A2(n_978), .B1(n_989), .B2(n_990), .Y(n_988) );
AOI22xp5_ASAP7_75t_L g1447 ( .A1(n_734), .A2(n_989), .B1(n_1422), .B2(n_1430), .Y(n_1447) );
AOI22xp5_ASAP7_75t_L g1799 ( .A1(n_734), .A2(n_989), .B1(n_1800), .B2(n_1801), .Y(n_1799) );
INVx1_ASAP7_75t_L g1860 ( .A(n_734), .Y(n_1860) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g1859 ( .A(n_736), .Y(n_1859) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
BUFx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g1171 ( .A(n_740), .Y(n_1171) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
A2O1A1Ixp33_ASAP7_75t_L g983 ( .A1(n_742), .A2(n_984), .B(n_985), .C(n_986), .Y(n_983) );
A2O1A1Ixp33_ASAP7_75t_L g1392 ( .A1(n_742), .A2(n_831), .B(n_1362), .C(n_1393), .Y(n_1392) );
A2O1A1Ixp33_ASAP7_75t_SL g1856 ( .A1(n_742), .A2(n_985), .B(n_1857), .C(n_1858), .Y(n_1856) );
INVx2_ASAP7_75t_L g822 ( .A(n_752), .Y(n_822) );
OAI31xp67_ASAP7_75t_L g1319 ( .A1(n_755), .A2(n_1320), .A3(n_1331), .B(n_1342), .Y(n_1319) );
BUFx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g1532 ( .A1(n_759), .A2(n_801), .B1(n_1516), .B2(n_1524), .Y(n_1532) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g1336 ( .A1(n_766), .A2(n_1006), .B1(n_1337), .B2(n_1338), .Y(n_1336) );
OAI33xp33_ASAP7_75t_L g906 ( .A1(n_767), .A2(n_817), .A3(n_907), .B1(n_908), .B2(n_910), .B3(n_912), .Y(n_906) );
OAI33xp33_ASAP7_75t_L g935 ( .A1(n_767), .A2(n_936), .A3(n_937), .B1(n_939), .B2(n_942), .B3(n_943), .Y(n_935) );
OAI33xp33_ASAP7_75t_L g1460 ( .A1(n_767), .A2(n_817), .A3(n_1461), .B1(n_1467), .B2(n_1470), .B3(n_1474), .Y(n_1460) );
INVx1_ASAP7_75t_L g799 ( .A(n_770), .Y(n_799) );
INVx1_ASAP7_75t_L g1247 ( .A(n_770), .Y(n_1247) );
AOI22xp33_ASAP7_75t_L g1874 ( .A1(n_771), .A2(n_1328), .B1(n_1857), .B2(n_1875), .Y(n_1874) );
INVx3_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
CKINVDCx5p33_ASAP7_75t_R g1327 ( .A(n_774), .Y(n_1327) );
INVx2_ASAP7_75t_L g1360 ( .A(n_774), .Y(n_1360) );
INVx8_ASAP7_75t_L g1365 ( .A(n_774), .Y(n_1365) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
AOI211xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_796), .B(n_797), .C(n_818), .Y(n_780) );
INVx2_ASAP7_75t_L g1136 ( .A(n_785), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_789), .B(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g816 ( .A(n_790), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_793), .B1(n_794), .B2(n_795), .Y(n_791) );
INVx2_ASAP7_75t_L g862 ( .A(n_793), .Y(n_862) );
INVx2_ASAP7_75t_L g946 ( .A(n_795), .Y(n_946) );
INVx1_ASAP7_75t_L g1082 ( .A(n_795), .Y(n_1082) );
OAI31xp33_ASAP7_75t_L g944 ( .A1(n_796), .A2(n_945), .A3(n_947), .B(n_953), .Y(n_944) );
OAI221xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_800), .B1(n_801), .B2(n_803), .C(n_804), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g1194 ( .A1(n_801), .A2(n_938), .B1(n_1195), .B2(n_1196), .Y(n_1194) );
OAI22xp5_ASAP7_75t_L g1345 ( .A1(n_801), .A2(n_1346), .B1(n_1348), .B2(n_1349), .Y(n_1345) );
OAI221xp5_ASAP7_75t_L g1863 ( .A1(n_801), .A2(n_1864), .B1(n_1865), .B2(n_1866), .C(n_1867), .Y(n_1863) );
OAI221xp5_ASAP7_75t_L g1868 ( .A1(n_801), .A2(n_1851), .B1(n_1869), .B2(n_1870), .C(n_1871), .Y(n_1868) );
CKINVDCx8_ASAP7_75t_R g801 ( .A(n_802), .Y(n_801) );
INVx3_ASAP7_75t_L g810 ( .A(n_802), .Y(n_810) );
INVx3_ASAP7_75t_L g1049 ( .A(n_802), .Y(n_1049) );
INVx1_ASAP7_75t_L g1150 ( .A(n_802), .Y(n_1150) );
INVx3_ASAP7_75t_L g1201 ( .A(n_802), .Y(n_1201) );
OAI221xp5_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_809), .B1(n_810), .B2(n_811), .C(n_812), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g1098 ( .A1(n_808), .A2(n_810), .B1(n_1099), .B2(n_1100), .Y(n_1098) );
OAI22xp5_ASAP7_75t_L g1101 ( .A1(n_808), .A2(n_1102), .B1(n_1103), .B2(n_1104), .Y(n_1101) );
OAI22xp5_ASAP7_75t_L g1147 ( .A1(n_808), .A2(n_1148), .B1(n_1149), .B2(n_1150), .Y(n_1147) );
OAI211xp5_ASAP7_75t_SL g832 ( .A1(n_809), .A2(n_827), .B(n_833), .C(n_834), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g910 ( .A1(n_810), .A2(n_889), .B1(n_905), .B2(n_911), .Y(n_910) );
OAI22xp5_ASAP7_75t_L g1151 ( .A1(n_810), .A2(n_1152), .B1(n_1153), .B2(n_1154), .Y(n_1151) );
OAI22xp5_ASAP7_75t_L g1529 ( .A1(n_810), .A2(n_1515), .B1(n_1522), .B2(n_1530), .Y(n_1529) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_820), .B(n_823), .Y(n_819) );
OAI211xp5_ASAP7_75t_L g825 ( .A1(n_826), .A2(n_827), .B(n_828), .C(n_830), .Y(n_825) );
BUFx2_ASAP7_75t_L g956 ( .A(n_827), .Y(n_956) );
OAI22xp5_ASAP7_75t_L g1112 ( .A1(n_827), .A2(n_1099), .B1(n_1102), .B2(n_1113), .Y(n_1112) );
OAI22xp5_ASAP7_75t_L g1114 ( .A1(n_827), .A2(n_1095), .B1(n_1107), .B2(n_1113), .Y(n_1114) );
BUFx6f_ASAP7_75t_L g985 ( .A(n_831), .Y(n_985) );
INVx3_ASAP7_75t_L g1380 ( .A(n_831), .Y(n_1380) );
A2O1A1Ixp33_ASAP7_75t_L g1445 ( .A1(n_831), .A2(n_1424), .B(n_1446), .C(n_1448), .Y(n_1445) );
INVx1_ASAP7_75t_L g966 ( .A(n_840), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_916), .B1(n_917), .B2(n_965), .Y(n_840) );
INVx1_ASAP7_75t_L g965 ( .A(n_841), .Y(n_965) );
NAND3xp33_ASAP7_75t_SL g842 ( .A(n_843), .B(n_860), .C(n_875), .Y(n_842) );
OAI211xp5_ASAP7_75t_L g991 ( .A1(n_845), .A2(n_992), .B(n_993), .C(n_995), .Y(n_991) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx2_ASAP7_75t_L g896 ( .A(n_846), .Y(n_896) );
INVx1_ASAP7_75t_L g987 ( .A(n_846), .Y(n_987) );
INVx2_ASAP7_75t_L g998 ( .A(n_846), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_850), .A2(n_951), .B1(n_958), .B2(n_959), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_850), .A2(n_959), .B1(n_1028), .B2(n_1029), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1505 ( .A1(n_850), .A2(n_1219), .B1(n_1495), .B2(n_1506), .Y(n_1505) );
BUFx3_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx2_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
OAI31xp33_ASAP7_75t_SL g860 ( .A1(n_861), .A2(n_864), .A3(n_871), .B(n_874), .Y(n_860) );
OAI22xp33_ASAP7_75t_L g1202 ( .A1(n_865), .A2(n_1009), .B1(n_1203), .B2(n_1204), .Y(n_1202) );
INVx2_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx2_ASAP7_75t_L g1018 ( .A(n_866), .Y(n_1018) );
OAI31xp33_ASAP7_75t_L g1072 ( .A1(n_874), .A2(n_1073), .A3(n_1077), .B(n_1081), .Y(n_1072) );
OAI31xp33_ASAP7_75t_L g1223 ( .A1(n_874), .A2(n_1224), .A3(n_1227), .B(n_1230), .Y(n_1223) );
OAI31xp33_ASAP7_75t_L g1267 ( .A1(n_874), .A2(n_1268), .A3(n_1269), .B(n_1272), .Y(n_1267) );
NOR2xp33_ASAP7_75t_SL g875 ( .A(n_876), .B(n_906), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_878), .A2(n_879), .B1(n_882), .B2(n_883), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_879), .A2(n_902), .B1(n_903), .B2(n_905), .Y(n_901) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_879), .A2(n_883), .B1(n_923), .B2(n_924), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_879), .A2(n_903), .B1(n_933), .B2(n_934), .Y(n_932) );
INVx2_ASAP7_75t_SL g879 ( .A(n_880), .Y(n_879) );
INVx2_ASAP7_75t_L g1255 ( .A(n_880), .Y(n_1255) );
INVx2_ASAP7_75t_L g1259 ( .A(n_880), .Y(n_1259) );
INVx3_ASAP7_75t_L g1523 ( .A(n_880), .Y(n_1523) );
BUFx6f_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx3_ASAP7_75t_L g1063 ( .A(n_881), .Y(n_1063) );
INVx4_ASAP7_75t_L g1401 ( .A(n_881), .Y(n_1401) );
OAI22xp33_ASAP7_75t_L g912 ( .A1(n_882), .A2(n_897), .B1(n_913), .B2(n_915), .Y(n_912) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_887), .A2(n_888), .B1(n_889), .B2(n_890), .Y(n_886) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_888), .A2(n_926), .B1(n_927), .B2(n_928), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_890), .A2(n_1047), .B1(n_1051), .B2(n_1068), .Y(n_1067) );
OAI22xp5_ASAP7_75t_L g1070 ( .A1(n_890), .A2(n_1042), .B1(n_1058), .B2(n_1068), .Y(n_1070) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_892), .A2(n_895), .B1(n_896), .B2(n_897), .Y(n_891) );
INVx3_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
INVx2_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
HB1xp67_ASAP7_75t_L g1484 ( .A(n_894), .Y(n_1484) );
INVx2_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
OAI33xp33_ASAP7_75t_L g920 ( .A1(n_900), .A2(n_921), .A3(n_922), .B1(n_925), .B2(n_929), .B3(n_932), .Y(n_920) );
OAI22xp5_ASAP7_75t_L g1485 ( .A1(n_903), .A2(n_1469), .B1(n_1473), .B2(n_1486), .Y(n_1485) );
BUFx3_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_911), .A2(n_1049), .B1(n_1051), .B2(n_1052), .Y(n_1050) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g1015 ( .A1(n_914), .A2(n_1016), .B1(n_1017), .B2(n_1018), .Y(n_1015) );
OAI22xp33_ASAP7_75t_L g1461 ( .A1(n_915), .A2(n_1462), .B1(n_1463), .B2(n_1466), .Y(n_1461) );
OAI22xp33_ASAP7_75t_L g1474 ( .A1(n_915), .A2(n_1463), .B1(n_1475), .B2(n_1476), .Y(n_1474) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
NAND3xp33_ASAP7_75t_L g918 ( .A(n_919), .B(n_944), .C(n_954), .Y(n_918) );
NOR2xp33_ASAP7_75t_L g919 ( .A(n_920), .B(n_935), .Y(n_919) );
INVx2_ASAP7_75t_SL g1110 ( .A(n_921), .Y(n_1110) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_927), .A2(n_934), .B1(n_940), .B2(n_941), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_940), .A2(n_1047), .B1(n_1048), .B2(n_1049), .Y(n_1046) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
OAI31xp33_ASAP7_75t_L g954 ( .A1(n_955), .A2(n_960), .A3(n_963), .B(n_964), .Y(n_954) );
HB1xp67_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
INVx2_ASAP7_75t_SL g1503 ( .A(n_962), .Y(n_1503) );
OAI31xp33_ASAP7_75t_L g1260 ( .A1(n_964), .A2(n_1261), .A3(n_1262), .B(n_1266), .Y(n_1260) );
OAI31xp33_ASAP7_75t_SL g1498 ( .A1(n_964), .A2(n_1499), .A3(n_1501), .B(n_1504), .Y(n_1498) );
AO22x2_ASAP7_75t_L g967 ( .A1(n_968), .A2(n_1020), .B1(n_1021), .B2(n_1084), .Y(n_967) );
INVx1_ASAP7_75t_SL g1084 ( .A(n_968), .Y(n_1084) );
XNOR2x1_ASAP7_75t_L g968 ( .A(n_969), .B(n_970), .Y(n_968) );
NOR2x1_ASAP7_75t_L g970 ( .A(n_971), .B(n_974), .Y(n_970) );
NAND3xp33_ASAP7_75t_SL g974 ( .A(n_975), .B(n_981), .C(n_1004), .Y(n_974) );
INVx2_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
OAI21xp5_ASAP7_75t_L g981 ( .A1(n_982), .A2(n_1001), .B(n_1003), .Y(n_981) );
NAND3xp33_ASAP7_75t_L g982 ( .A(n_983), .B(n_991), .C(n_996), .Y(n_982) );
NAND2xp5_ASAP7_75t_SL g986 ( .A(n_987), .B(n_988), .Y(n_986) );
OAI211xp5_ASAP7_75t_L g996 ( .A1(n_997), .A2(n_998), .B(n_999), .C(n_1000), .Y(n_996) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_997), .A2(n_1008), .B1(n_1009), .B2(n_1010), .Y(n_1007) );
OAI22xp33_ASAP7_75t_L g1093 ( .A1(n_1009), .A2(n_1094), .B1(n_1095), .B2(n_1096), .Y(n_1093) );
OAI22xp33_ASAP7_75t_L g1143 ( .A1(n_1009), .A2(n_1144), .B1(n_1145), .B2(n_1146), .Y(n_1143) );
INVx2_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
INVx2_ASAP7_75t_L g1132 ( .A(n_1011), .Y(n_1132) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1011), .Y(n_1528) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
OAI211xp5_ASAP7_75t_L g1350 ( .A1(n_1018), .A2(n_1301), .B(n_1351), .C(n_1353), .Y(n_1350) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
NAND3xp33_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1036), .C(n_1072), .Y(n_1023) );
NOR2xp33_ASAP7_75t_SL g1036 ( .A(n_1037), .B(n_1059), .Y(n_1036) );
OAI22xp5_ASAP7_75t_L g1038 ( .A1(n_1039), .A2(n_1040), .B1(n_1042), .B2(n_1043), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g1060 ( .A1(n_1039), .A2(n_1057), .B1(n_1061), .B2(n_1064), .Y(n_1060) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
INVx2_ASAP7_75t_SL g1043 ( .A(n_1044), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
HB1xp67_ASAP7_75t_L g1193 ( .A(n_1045), .Y(n_1193) );
OAI22xp5_ASAP7_75t_L g1071 ( .A1(n_1048), .A2(n_1052), .B1(n_1061), .B2(n_1064), .Y(n_1071) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
BUFx2_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
INVx2_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
INVx2_ASAP7_75t_SL g1062 ( .A(n_1063), .Y(n_1062) );
INVx2_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
INVx2_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
OAI22xp33_ASAP7_75t_L g1162 ( .A1(n_1066), .A2(n_1144), .B1(n_1156), .B2(n_1163), .Y(n_1162) );
OAI22xp5_ASAP7_75t_L g1399 ( .A1(n_1066), .A2(n_1400), .B1(n_1401), .B2(n_1402), .Y(n_1399) );
INVx1_ASAP7_75t_L g1482 ( .A(n_1068), .Y(n_1482) );
INVx2_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
BUFx2_ASAP7_75t_L g1211 ( .A(n_1069), .Y(n_1211) );
INVx2_ASAP7_75t_L g1384 ( .A(n_1069), .Y(n_1384) );
INVx2_ASAP7_75t_SL g1074 ( .A(n_1075), .Y(n_1074) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1085), .Y(n_1409) );
XOR2xp5_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1275), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1086 ( .A1(n_1087), .A2(n_1185), .B1(n_1273), .B2(n_1274), .Y(n_1086) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1087), .Y(n_1274) );
XOR2xp5_ASAP7_75t_L g1087 ( .A(n_1088), .B(n_1138), .Y(n_1087) );
NAND3xp33_ASAP7_75t_L g1089 ( .A(n_1090), .B(n_1118), .C(n_1128), .Y(n_1089) );
NOR2xp33_ASAP7_75t_L g1090 ( .A(n_1091), .B(n_1108), .Y(n_1090) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1097), .Y(n_1146) );
INVxp67_ASAP7_75t_L g1493 ( .A(n_1097), .Y(n_1493) );
OAI33xp33_ASAP7_75t_L g1108 ( .A1(n_1109), .A2(n_1111), .A3(n_1112), .B1(n_1114), .B2(n_1115), .B3(n_1117), .Y(n_1108) );
OAI33xp33_ASAP7_75t_L g1510 ( .A1(n_1109), .A2(n_1307), .A3(n_1511), .B1(n_1514), .B2(n_1517), .B3(n_1521), .Y(n_1510) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
OAI33xp33_ASAP7_75t_L g1159 ( .A1(n_1115), .A2(n_1160), .A3(n_1161), .B1(n_1162), .B2(n_1164), .B3(n_1165), .Y(n_1159) );
INVx2_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
INVx2_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
INVx2_ASAP7_75t_L g1219 ( .A(n_1123), .Y(n_1219) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1127), .Y(n_1545) );
OAI31xp33_ASAP7_75t_L g1128 ( .A1(n_1129), .A2(n_1130), .A3(n_1135), .B(n_1137), .Y(n_1128) );
HB1xp67_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
OAI31xp33_ASAP7_75t_SL g1177 ( .A1(n_1137), .A2(n_1178), .A3(n_1180), .B(n_1181), .Y(n_1177) );
OAI31xp33_ASAP7_75t_L g1533 ( .A1(n_1137), .A2(n_1534), .A3(n_1536), .B(n_1540), .Y(n_1533) );
XNOR2xp5_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1140), .Y(n_1138) );
AND3x1_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1166), .C(n_1177), .Y(n_1140) );
NOR2xp33_ASAP7_75t_SL g1141 ( .A(n_1142), .B(n_1159), .Y(n_1141) );
OAI31xp33_ASAP7_75t_L g1166 ( .A1(n_1167), .A2(n_1168), .A3(n_1175), .B(n_1176), .Y(n_1166) );
INVx2_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
INVx2_ASAP7_75t_L g1547 ( .A(n_1170), .Y(n_1547) );
OAI31xp33_ASAP7_75t_SL g1542 ( .A1(n_1176), .A2(n_1543), .A3(n_1546), .B(n_1550), .Y(n_1542) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1185), .Y(n_1273) );
XOR2x2_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1233), .Y(n_1185) );
AND3x1_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1214), .C(n_1223), .Y(n_1187) );
NOR2xp33_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1205), .Y(n_1188) );
OAI22xp5_ASAP7_75t_L g1197 ( .A1(n_1198), .A2(n_1199), .B1(n_1200), .B2(n_1201), .Y(n_1197) );
OAI22xp5_ASAP7_75t_L g1470 ( .A1(n_1201), .A2(n_1471), .B1(n_1472), .B2(n_1473), .Y(n_1470) );
BUFx6f_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
INVx4_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
AND3x1_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1260), .C(n_1267), .Y(n_1234) );
NOR2xp33_ASAP7_75t_L g1235 ( .A(n_1236), .B(n_1253), .Y(n_1235) );
HB1xp67_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
XOR2xp5_ASAP7_75t_L g1276 ( .A(n_1277), .B(n_1354), .Y(n_1276) );
XNOR2x1_ASAP7_75t_L g1277 ( .A(n_1278), .B(n_1279), .Y(n_1277) );
NAND4xp75_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1288), .C(n_1316), .D(n_1319), .Y(n_1279) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
AOI211x1_ASAP7_75t_L g1288 ( .A1(n_1289), .A2(n_1298), .B(n_1299), .C(n_1312), .Y(n_1288) );
OAI22xp5_ASAP7_75t_L g1292 ( .A1(n_1293), .A2(n_1294), .B1(n_1295), .B2(n_1297), .Y(n_1292) );
BUFx6f_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
OAI21xp5_ASAP7_75t_L g1299 ( .A1(n_1300), .A2(n_1307), .B(n_1308), .Y(n_1299) );
OAI221xp5_ASAP7_75t_L g1300 ( .A1(n_1301), .A2(n_1302), .B1(n_1304), .B2(n_1305), .C(n_1306), .Y(n_1300) );
INVx2_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
OAI211xp5_ASAP7_75t_SL g1846 ( .A1(n_1304), .A2(n_1847), .B(n_1848), .C(n_1849), .Y(n_1846) );
OAI211xp5_ASAP7_75t_SL g1850 ( .A1(n_1304), .A2(n_1851), .B(n_1852), .C(n_1854), .Y(n_1850) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
NAND2x2_ASAP7_75t_L g1313 ( .A(n_1310), .B(n_1314), .Y(n_1313) );
INVx2_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
INVx2_ASAP7_75t_SL g1314 ( .A(n_1315), .Y(n_1314) );
AOI22xp33_ASAP7_75t_L g1332 ( .A1(n_1317), .A2(n_1318), .B1(n_1333), .B2(n_1334), .Y(n_1332) );
INVx4_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
INVx2_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
A2O1A1Ixp33_ASAP7_75t_L g1325 ( .A1(n_1326), .A2(n_1327), .B(n_1328), .C(n_1329), .Y(n_1325) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
AOI21xp33_ASAP7_75t_L g1331 ( .A1(n_1332), .A2(n_1336), .B(n_1339), .Y(n_1331) );
INVx2_ASAP7_75t_L g1472 ( .A(n_1334), .Y(n_1472) );
INVx2_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1340), .Y(n_1339) );
HB1xp67_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
OAI21xp5_ASAP7_75t_SL g1342 ( .A1(n_1343), .A2(n_1345), .B(n_1350), .Y(n_1342) );
INVx2_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
INVx2_ASAP7_75t_SL g1864 ( .A(n_1347), .Y(n_1864) );
XNOR2x1_ASAP7_75t_L g1354 ( .A(n_1355), .B(n_1406), .Y(n_1354) );
OR2x2_ASAP7_75t_L g1355 ( .A(n_1356), .B(n_1373), .Y(n_1355) );
NAND3xp33_ASAP7_75t_L g1356 ( .A(n_1357), .B(n_1363), .C(n_1371), .Y(n_1356) );
INVx2_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
NAND3xp33_ASAP7_75t_SL g1373 ( .A(n_1374), .B(n_1377), .C(n_1403), .Y(n_1373) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
OAI21xp33_ASAP7_75t_L g1385 ( .A1(n_1386), .A2(n_1388), .B(n_1392), .Y(n_1385) );
OAI21xp5_ASAP7_75t_SL g1441 ( .A1(n_1386), .A2(n_1442), .B(n_1445), .Y(n_1441) );
INVxp67_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
AOI22xp5_ASAP7_75t_L g1797 ( .A1(n_1387), .A2(n_1448), .B1(n_1798), .B2(n_1802), .Y(n_1797) );
OAI21xp5_ASAP7_75t_L g1843 ( .A1(n_1387), .A2(n_1844), .B(n_1845), .Y(n_1843) );
INVx2_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
NAND2xp5_ASAP7_75t_L g1403 ( .A(n_1404), .B(n_1405), .Y(n_1403) );
NAND2xp5_ASAP7_75t_L g1432 ( .A(n_1405), .B(n_1433), .Y(n_1432) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1411), .Y(n_1410) );
AOI22xp5_ASAP7_75t_L g1411 ( .A1(n_1412), .A2(n_1454), .B1(n_1552), .B2(n_1553), .Y(n_1411) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1412), .Y(n_1552) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
XNOR2x1_ASAP7_75t_L g1413 ( .A(n_1414), .B(n_1453), .Y(n_1413) );
OR2x2_ASAP7_75t_L g1414 ( .A(n_1415), .B(n_1428), .Y(n_1414) );
NAND4xp25_ASAP7_75t_SL g1415 ( .A(n_1416), .B(n_1419), .C(n_1421), .D(n_1425), .Y(n_1415) );
NAND3xp33_ASAP7_75t_SL g1428 ( .A(n_1429), .B(n_1432), .C(n_1434), .Y(n_1428) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
INVx1_ASAP7_75t_L g1553 ( .A(n_1454), .Y(n_1553) );
AOI22xp33_ASAP7_75t_L g1454 ( .A1(n_1455), .A2(n_1456), .B1(n_1507), .B2(n_1551), .Y(n_1454) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
HB1xp67_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
AND3x1_ASAP7_75t_L g1458 ( .A(n_1459), .B(n_1490), .C(n_1498), .Y(n_1458) );
NOR2xp33_ASAP7_75t_L g1459 ( .A(n_1460), .B(n_1477), .Y(n_1459) );
INVx2_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1465), .Y(n_1464) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
INVx1_ASAP7_75t_L g1488 ( .A(n_1489), .Y(n_1488) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1503), .Y(n_1502) );
INVx2_ASAP7_75t_SL g1551 ( .A(n_1507), .Y(n_1551) );
NAND3xp33_ASAP7_75t_L g1508 ( .A(n_1509), .B(n_1533), .C(n_1542), .Y(n_1508) );
NOR2xp33_ASAP7_75t_L g1509 ( .A(n_1510), .B(n_1526), .Y(n_1509) );
OAI22xp5_ASAP7_75t_L g1521 ( .A1(n_1522), .A2(n_1523), .B1(n_1524), .B2(n_1525), .Y(n_1521) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
OAI221xp5_ASAP7_75t_SL g1554 ( .A1(n_1555), .A2(n_1780), .B1(n_1783), .B2(n_1827), .C(n_1833), .Y(n_1554) );
NOR5xp2_ASAP7_75t_L g1555 ( .A(n_1556), .B(n_1695), .C(n_1757), .D(n_1763), .E(n_1774), .Y(n_1555) );
AOI31xp33_ASAP7_75t_L g1556 ( .A1(n_1557), .A2(n_1639), .A3(n_1669), .B(n_1689), .Y(n_1556) );
AOI211xp5_ASAP7_75t_SL g1557 ( .A1(n_1558), .A2(n_1574), .B(n_1593), .C(n_1607), .Y(n_1557) );
A2O1A1Ixp33_ASAP7_75t_L g1696 ( .A1(n_1558), .A2(n_1697), .B(n_1699), .C(n_1711), .Y(n_1696) );
CKINVDCx6p67_ASAP7_75t_R g1558 ( .A(n_1559), .Y(n_1558) );
CKINVDCx6p67_ASAP7_75t_R g1559 ( .A(n_1560), .Y(n_1559) );
AND2x2_ASAP7_75t_L g1637 ( .A(n_1560), .B(n_1635), .Y(n_1637) );
INVx2_ASAP7_75t_L g1647 ( .A(n_1560), .Y(n_1647) );
NAND2xp5_ASAP7_75t_L g1706 ( .A(n_1560), .B(n_1707), .Y(n_1706) );
OAI22xp5_ASAP7_75t_L g1717 ( .A1(n_1560), .A2(n_1718), .B1(n_1720), .B2(n_1722), .Y(n_1717) );
AND2x4_ASAP7_75t_L g1560 ( .A(n_1561), .B(n_1568), .Y(n_1560) );
AND2x2_ASAP7_75t_L g1599 ( .A(n_1561), .B(n_1568), .Y(n_1599) );
INVx2_ASAP7_75t_L g1782 ( .A(n_1562), .Y(n_1782) );
AND2x6_ASAP7_75t_L g1562 ( .A(n_1563), .B(n_1564), .Y(n_1562) );
AND2x2_ASAP7_75t_L g1566 ( .A(n_1563), .B(n_1567), .Y(n_1566) );
AND2x4_ASAP7_75t_L g1569 ( .A(n_1563), .B(n_1570), .Y(n_1569) );
AND2x6_ASAP7_75t_L g1572 ( .A(n_1563), .B(n_1573), .Y(n_1572) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1563), .B(n_1567), .Y(n_1580) );
AND2x2_ASAP7_75t_L g1584 ( .A(n_1563), .B(n_1567), .Y(n_1584) );
OAI21xp5_ASAP7_75t_L g1887 ( .A1(n_1564), .A2(n_1888), .B(n_1889), .Y(n_1887) );
AND2x2_ASAP7_75t_L g1570 ( .A(n_1565), .B(n_1571), .Y(n_1570) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
NAND2xp5_ASAP7_75t_L g1575 ( .A(n_1576), .B(n_1581), .Y(n_1575) );
AND2x2_ASAP7_75t_L g1621 ( .A(n_1576), .B(n_1622), .Y(n_1621) );
NAND2xp5_ASAP7_75t_SL g1643 ( .A(n_1576), .B(n_1644), .Y(n_1643) );
OR2x2_ASAP7_75t_L g1722 ( .A(n_1576), .B(n_1723), .Y(n_1722) );
INVx2_ASAP7_75t_L g1726 ( .A(n_1576), .Y(n_1726) );
INVx2_ASAP7_75t_L g1576 ( .A(n_1577), .Y(n_1576) );
INVx3_ASAP7_75t_L g1601 ( .A(n_1577), .Y(n_1601) );
NOR2xp33_ASAP7_75t_L g1619 ( .A(n_1577), .B(n_1582), .Y(n_1619) );
NAND2xp5_ASAP7_75t_L g1651 ( .A(n_1577), .B(n_1652), .Y(n_1651) );
AND2x2_ASAP7_75t_L g1674 ( .A(n_1577), .B(n_1582), .Y(n_1674) );
AND2x2_ASAP7_75t_L g1678 ( .A(n_1577), .B(n_1616), .Y(n_1678) );
NAND2xp5_ASAP7_75t_L g1708 ( .A(n_1577), .B(n_1665), .Y(n_1708) );
NOR2xp33_ASAP7_75t_L g1716 ( .A(n_1577), .B(n_1627), .Y(n_1716) );
AND2x2_ASAP7_75t_L g1577 ( .A(n_1578), .B(n_1579), .Y(n_1577) );
NAND2xp5_ASAP7_75t_L g1761 ( .A(n_1581), .B(n_1611), .Y(n_1761) );
AND2x2_ASAP7_75t_L g1581 ( .A(n_1582), .B(n_1586), .Y(n_1581) );
CKINVDCx5p33_ASAP7_75t_R g1642 ( .A(n_1582), .Y(n_1642) );
NAND2xp5_ASAP7_75t_L g1653 ( .A(n_1582), .B(n_1654), .Y(n_1653) );
AND2x2_ASAP7_75t_L g1731 ( .A(n_1582), .B(n_1605), .Y(n_1731) );
OR2x2_ASAP7_75t_L g1743 ( .A(n_1582), .B(n_1618), .Y(n_1743) );
NAND2xp5_ASAP7_75t_L g1746 ( .A(n_1582), .B(n_1679), .Y(n_1746) );
AND2x2_ASAP7_75t_L g1582 ( .A(n_1583), .B(n_1585), .Y(n_1582) );
AND2x2_ASAP7_75t_L g1603 ( .A(n_1583), .B(n_1585), .Y(n_1603) );
INVx1_ASAP7_75t_L g1627 ( .A(n_1586), .Y(n_1627) );
AND2x2_ASAP7_75t_L g1684 ( .A(n_1586), .B(n_1674), .Y(n_1684) );
AND2x2_ASAP7_75t_L g1704 ( .A(n_1586), .B(n_1642), .Y(n_1704) );
AND2x2_ASAP7_75t_L g1586 ( .A(n_1587), .B(n_1590), .Y(n_1586) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1587), .Y(n_1606) );
INVx1_ASAP7_75t_L g1679 ( .A(n_1587), .Y(n_1679) );
NAND2xp5_ASAP7_75t_L g1587 ( .A(n_1588), .B(n_1589), .Y(n_1587) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1590), .Y(n_1605) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1590), .Y(n_1618) );
AND2x2_ASAP7_75t_L g1631 ( .A(n_1590), .B(n_1606), .Y(n_1631) );
OR2x2_ASAP7_75t_L g1645 ( .A(n_1590), .B(n_1606), .Y(n_1645) );
NAND2xp5_ASAP7_75t_L g1590 ( .A(n_1591), .B(n_1592), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1593 ( .A(n_1594), .B(n_1600), .Y(n_1593) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
OR2x2_ASAP7_75t_L g1595 ( .A(n_1596), .B(n_1599), .Y(n_1595) );
INVx3_ASAP7_75t_L g1616 ( .A(n_1596), .Y(n_1616) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1596), .B(n_1633), .Y(n_1632) );
AND2x2_ASAP7_75t_L g1646 ( .A(n_1596), .B(n_1647), .Y(n_1646) );
OR2x2_ASAP7_75t_L g1649 ( .A(n_1596), .B(n_1634), .Y(n_1649) );
NOR2xp33_ASAP7_75t_L g1657 ( .A(n_1596), .B(n_1610), .Y(n_1657) );
NAND2xp5_ASAP7_75t_L g1671 ( .A(n_1596), .B(n_1599), .Y(n_1671) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1596), .B(n_1610), .Y(n_1685) );
AND2x2_ASAP7_75t_L g1688 ( .A(n_1596), .B(n_1661), .Y(n_1688) );
AND2x2_ASAP7_75t_L g1721 ( .A(n_1596), .B(n_1665), .Y(n_1721) );
AND2x2_ASAP7_75t_L g1729 ( .A(n_1596), .B(n_1711), .Y(n_1729) );
INVx3_ASAP7_75t_L g1773 ( .A(n_1596), .Y(n_1773) );
AND2x4_ASAP7_75t_SL g1596 ( .A(n_1597), .B(n_1598), .Y(n_1596) );
AND2x2_ASAP7_75t_L g1615 ( .A(n_1599), .B(n_1616), .Y(n_1615) );
OR2x2_ASAP7_75t_L g1623 ( .A(n_1599), .B(n_1612), .Y(n_1623) );
OR2x2_ASAP7_75t_L g1634 ( .A(n_1599), .B(n_1635), .Y(n_1634) );
AND2x2_ASAP7_75t_L g1661 ( .A(n_1599), .B(n_1612), .Y(n_1661) );
NOR2xp33_ASAP7_75t_L g1744 ( .A(n_1599), .B(n_1692), .Y(n_1744) );
AND2x2_ASAP7_75t_L g1600 ( .A(n_1601), .B(n_1602), .Y(n_1600) );
INVx1_ASAP7_75t_L g1660 ( .A(n_1601), .Y(n_1660) );
AND2x2_ASAP7_75t_L g1698 ( .A(n_1601), .B(n_1631), .Y(n_1698) );
NOR2xp33_ASAP7_75t_L g1701 ( .A(n_1601), .B(n_1645), .Y(n_1701) );
O2A1O1Ixp33_ASAP7_75t_L g1703 ( .A1(n_1601), .A2(n_1661), .B(n_1704), .C(n_1705), .Y(n_1703) );
NAND2xp5_ASAP7_75t_L g1733 ( .A(n_1601), .B(n_1635), .Y(n_1733) );
NAND2xp5_ASAP7_75t_L g1736 ( .A(n_1601), .B(n_1737), .Y(n_1736) );
NOR2xp33_ASAP7_75t_L g1742 ( .A(n_1601), .B(n_1743), .Y(n_1742) );
NOR2xp33_ASAP7_75t_L g1745 ( .A(n_1601), .B(n_1746), .Y(n_1745) );
NAND3xp33_ASAP7_75t_L g1749 ( .A(n_1601), .B(n_1711), .C(n_1750), .Y(n_1749) );
NAND2xp5_ASAP7_75t_L g1766 ( .A(n_1601), .B(n_1633), .Y(n_1766) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1602), .Y(n_1662) );
AND2x2_ASAP7_75t_L g1602 ( .A(n_1603), .B(n_1604), .Y(n_1602) );
AOI32xp33_ASAP7_75t_L g1620 ( .A1(n_1603), .A2(n_1621), .A3(n_1624), .B1(n_1628), .B2(n_1632), .Y(n_1620) );
OR2x2_ASAP7_75t_L g1629 ( .A(n_1603), .B(n_1630), .Y(n_1629) );
OR2x2_ASAP7_75t_L g1667 ( .A(n_1603), .B(n_1668), .Y(n_1667) );
AND2x2_ASAP7_75t_L g1697 ( .A(n_1603), .B(n_1698), .Y(n_1697) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1604), .Y(n_1626) );
AND2x2_ASAP7_75t_L g1681 ( .A(n_1604), .B(n_1642), .Y(n_1681) );
AND2x2_ASAP7_75t_L g1683 ( .A(n_1604), .B(n_1619), .Y(n_1683) );
NAND2xp5_ASAP7_75t_L g1687 ( .A(n_1604), .B(n_1688), .Y(n_1687) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1605), .B(n_1606), .Y(n_1604) );
INVx1_ASAP7_75t_L g1654 ( .A(n_1606), .Y(n_1654) );
OAI211xp5_ASAP7_75t_L g1607 ( .A1(n_1608), .A2(n_1617), .B(n_1620), .C(n_1636), .Y(n_1607) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1609), .Y(n_1608) );
AND2x2_ASAP7_75t_L g1609 ( .A(n_1610), .B(n_1615), .Y(n_1609) );
AND2x2_ASAP7_75t_L g1719 ( .A(n_1610), .B(n_1673), .Y(n_1719) );
O2A1O1Ixp33_ASAP7_75t_L g1767 ( .A1(n_1610), .A2(n_1698), .B(n_1704), .C(n_1768), .Y(n_1767) );
INVx1_ASAP7_75t_L g1770 ( .A(n_1610), .Y(n_1770) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1611), .Y(n_1610) );
AND2x2_ASAP7_75t_L g1672 ( .A(n_1611), .B(n_1673), .Y(n_1672) );
AOI322xp5_ASAP7_75t_L g1741 ( .A1(n_1611), .A2(n_1657), .A3(n_1683), .B1(n_1729), .B2(n_1742), .C1(n_1744), .C2(n_1745), .Y(n_1741) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1612), .Y(n_1611) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1612), .Y(n_1635) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1612), .Y(n_1665) );
NAND2xp5_ASAP7_75t_L g1612 ( .A(n_1613), .B(n_1614), .Y(n_1612) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1615), .Y(n_1762) );
NAND2xp5_ASAP7_75t_L g1740 ( .A(n_1616), .B(n_1622), .Y(n_1740) );
OR2x2_ASAP7_75t_L g1752 ( .A(n_1616), .B(n_1623), .Y(n_1752) );
AOI32xp33_ASAP7_75t_L g1776 ( .A1(n_1616), .A2(n_1621), .A3(n_1710), .B1(n_1711), .B2(n_1777), .Y(n_1776) );
NAND2xp5_ASAP7_75t_L g1617 ( .A(n_1618), .B(n_1619), .Y(n_1617) );
INVx1_ASAP7_75t_L g1754 ( .A(n_1618), .Y(n_1754) );
AND2x2_ASAP7_75t_L g1638 ( .A(n_1619), .B(n_1631), .Y(n_1638) );
AOI311xp33_ASAP7_75t_L g1724 ( .A1(n_1622), .A2(n_1725), .A3(n_1726), .B(n_1727), .C(n_1738), .Y(n_1724) );
INVx1_ASAP7_75t_L g1622 ( .A(n_1623), .Y(n_1622) );
OAI321xp33_ASAP7_75t_L g1675 ( .A1(n_1623), .A2(n_1676), .A3(n_1677), .B1(n_1679), .B2(n_1680), .C(n_1682), .Y(n_1675) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
NAND2xp5_ASAP7_75t_L g1625 ( .A(n_1626), .B(n_1627), .Y(n_1625) );
INVx1_ASAP7_75t_L g1628 ( .A(n_1629), .Y(n_1628) );
OR2x2_ASAP7_75t_L g1779 ( .A(n_1630), .B(n_1642), .Y(n_1779) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
NAND2xp5_ASAP7_75t_L g1668 ( .A(n_1631), .B(n_1660), .Y(n_1668) );
AND2x2_ASAP7_75t_L g1673 ( .A(n_1631), .B(n_1674), .Y(n_1673) );
AND2x2_ASAP7_75t_L g1756 ( .A(n_1633), .B(n_1660), .Y(n_1756) );
INVx2_ASAP7_75t_SL g1633 ( .A(n_1634), .Y(n_1633) );
NAND2xp5_ASAP7_75t_L g1636 ( .A(n_1637), .B(n_1638), .Y(n_1636) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1637), .Y(n_1676) );
AOI221xp5_ASAP7_75t_L g1639 ( .A1(n_1640), .A2(n_1646), .B1(n_1648), .B2(n_1650), .C(n_1655), .Y(n_1639) );
INVx1_ASAP7_75t_L g1640 ( .A(n_1641), .Y(n_1640) );
OR2x2_ASAP7_75t_L g1641 ( .A(n_1642), .B(n_1643), .Y(n_1641) );
AND2x2_ASAP7_75t_L g1710 ( .A(n_1642), .B(n_1679), .Y(n_1710) );
AND2x2_ASAP7_75t_L g1713 ( .A(n_1642), .B(n_1701), .Y(n_1713) );
AND2x2_ASAP7_75t_L g1737 ( .A(n_1642), .B(n_1654), .Y(n_1737) );
NAND2xp5_ASAP7_75t_L g1739 ( .A(n_1644), .B(n_1674), .Y(n_1739) );
INVx1_ASAP7_75t_L g1644 ( .A(n_1645), .Y(n_1644) );
INVx1_ASAP7_75t_L g1702 ( .A(n_1646), .Y(n_1702) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1649), .Y(n_1648) );
INVxp67_ASAP7_75t_SL g1650 ( .A(n_1651), .Y(n_1650) );
INVx1_ASAP7_75t_L g1652 ( .A(n_1653), .Y(n_1652) );
A2O1A1Ixp33_ASAP7_75t_L g1655 ( .A1(n_1656), .A2(n_1658), .B(n_1662), .C(n_1663), .Y(n_1655) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1657), .Y(n_1656) );
INVx1_ASAP7_75t_L g1658 ( .A(n_1659), .Y(n_1658) );
AND2x2_ASAP7_75t_L g1659 ( .A(n_1660), .B(n_1661), .Y(n_1659) );
CKINVDCx14_ASAP7_75t_R g1775 ( .A(n_1661), .Y(n_1775) );
NAND2xp5_ASAP7_75t_L g1725 ( .A(n_1662), .B(n_1723), .Y(n_1725) );
NAND2xp5_ASAP7_75t_L g1663 ( .A(n_1664), .B(n_1666), .Y(n_1663) );
NAND2xp5_ASAP7_75t_L g1758 ( .A(n_1664), .B(n_1759), .Y(n_1758) );
INVx1_ASAP7_75t_L g1664 ( .A(n_1665), .Y(n_1664) );
INVx1_ASAP7_75t_L g1666 ( .A(n_1667), .Y(n_1666) );
NAND2xp5_ASAP7_75t_L g1714 ( .A(n_1667), .B(n_1715), .Y(n_1714) );
AOI211xp5_ASAP7_75t_L g1669 ( .A1(n_1670), .A2(n_1672), .B(n_1675), .C(n_1686), .Y(n_1669) );
NAND3xp33_ASAP7_75t_L g1734 ( .A(n_1670), .B(n_1691), .C(n_1735), .Y(n_1734) );
INVx1_ASAP7_75t_L g1670 ( .A(n_1671), .Y(n_1670) );
A2O1A1Ixp33_ASAP7_75t_L g1727 ( .A1(n_1671), .A2(n_1728), .B(n_1730), .C(n_1734), .Y(n_1727) );
NOR2xp33_ASAP7_75t_L g1705 ( .A(n_1676), .B(n_1680), .Y(n_1705) );
OAI221xp5_ASAP7_75t_SL g1738 ( .A1(n_1676), .A2(n_1680), .B1(n_1739), .B2(n_1740), .C(n_1741), .Y(n_1738) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1678), .Y(n_1677) );
INVx1_ASAP7_75t_L g1750 ( .A(n_1679), .Y(n_1750) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
OAI21xp5_ASAP7_75t_L g1682 ( .A1(n_1683), .A2(n_1684), .B(n_1685), .Y(n_1682) );
NAND2xp5_ASAP7_75t_L g1769 ( .A(n_1684), .B(n_1770), .Y(n_1769) );
AOI221xp5_ASAP7_75t_L g1712 ( .A1(n_1685), .A2(n_1688), .B1(n_1713), .B2(n_1714), .C(n_1717), .Y(n_1712) );
INVx1_ASAP7_75t_L g1778 ( .A(n_1685), .Y(n_1778) );
INVxp67_ASAP7_75t_SL g1686 ( .A(n_1687), .Y(n_1686) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1690), .Y(n_1689) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1691), .Y(n_1690) );
AND2x2_ASAP7_75t_L g1772 ( .A(n_1691), .B(n_1773), .Y(n_1772) );
INVx1_ASAP7_75t_L g1691 ( .A(n_1692), .Y(n_1691) );
INVx1_ASAP7_75t_L g1711 ( .A(n_1692), .Y(n_1711) );
AND2x2_ASAP7_75t_L g1692 ( .A(n_1693), .B(n_1694), .Y(n_1692) );
NAND4xp25_ASAP7_75t_L g1695 ( .A(n_1696), .B(n_1712), .C(n_1724), .D(n_1747), .Y(n_1695) );
CKINVDCx14_ASAP7_75t_R g1760 ( .A(n_1697), .Y(n_1760) );
OAI211xp5_ASAP7_75t_SL g1699 ( .A1(n_1700), .A2(n_1702), .B(n_1703), .C(n_1706), .Y(n_1699) );
INVx1_ASAP7_75t_L g1700 ( .A(n_1701), .Y(n_1700) );
INVx1_ASAP7_75t_L g1723 ( .A(n_1704), .Y(n_1723) );
O2A1O1Ixp33_ASAP7_75t_L g1747 ( .A1(n_1704), .A2(n_1748), .B(n_1751), .C(n_1753), .Y(n_1747) );
NOR2xp33_ASAP7_75t_L g1707 ( .A(n_1708), .B(n_1709), .Y(n_1707) );
INVx1_ASAP7_75t_L g1709 ( .A(n_1710), .Y(n_1709) );
INVx1_ASAP7_75t_L g1715 ( .A(n_1716), .Y(n_1715) );
INVx1_ASAP7_75t_L g1718 ( .A(n_1719), .Y(n_1718) );
INVx1_ASAP7_75t_L g1720 ( .A(n_1721), .Y(n_1720) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1722), .Y(n_1759) );
O2A1O1Ixp33_ASAP7_75t_L g1753 ( .A1(n_1728), .A2(n_1739), .B(n_1754), .C(n_1755), .Y(n_1753) );
INVx1_ASAP7_75t_L g1728 ( .A(n_1729), .Y(n_1728) );
NAND2xp5_ASAP7_75t_L g1730 ( .A(n_1731), .B(n_1732), .Y(n_1730) );
O2A1O1Ixp33_ASAP7_75t_L g1763 ( .A1(n_1731), .A2(n_1764), .B(n_1767), .C(n_1771), .Y(n_1763) );
INVx1_ASAP7_75t_L g1732 ( .A(n_1733), .Y(n_1732) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1736), .Y(n_1735) );
INVxp67_ASAP7_75t_SL g1748 ( .A(n_1749), .Y(n_1748) );
INVx1_ASAP7_75t_L g1751 ( .A(n_1752), .Y(n_1751) );
A2O1A1Ixp33_ASAP7_75t_L g1774 ( .A1(n_1752), .A2(n_1760), .B(n_1775), .C(n_1776), .Y(n_1774) );
INVxp67_ASAP7_75t_L g1755 ( .A(n_1756), .Y(n_1755) );
AOI31xp33_ASAP7_75t_L g1757 ( .A1(n_1758), .A2(n_1760), .A3(n_1761), .B(n_1762), .Y(n_1757) );
INVxp67_ASAP7_75t_L g1764 ( .A(n_1765), .Y(n_1764) );
INVx1_ASAP7_75t_L g1765 ( .A(n_1766), .Y(n_1765) );
INVx1_ASAP7_75t_L g1768 ( .A(n_1769), .Y(n_1768) );
INVx1_ASAP7_75t_L g1771 ( .A(n_1772), .Y(n_1771) );
NOR2xp33_ASAP7_75t_L g1777 ( .A(n_1778), .B(n_1779), .Y(n_1777) );
CKINVDCx20_ASAP7_75t_R g1780 ( .A(n_1781), .Y(n_1780) );
CKINVDCx20_ASAP7_75t_R g1781 ( .A(n_1782), .Y(n_1781) );
CKINVDCx6p67_ASAP7_75t_R g1783 ( .A(n_1784), .Y(n_1783) );
HB1xp67_ASAP7_75t_L g1784 ( .A(n_1785), .Y(n_1784) );
HB1xp67_ASAP7_75t_L g1785 ( .A(n_1786), .Y(n_1785) );
INVx1_ASAP7_75t_L g1786 ( .A(n_1787), .Y(n_1786) );
NAND3xp33_ASAP7_75t_L g1787 ( .A(n_1788), .B(n_1820), .C(n_1824), .Y(n_1787) );
INVx1_ASAP7_75t_L g1821 ( .A(n_1789), .Y(n_1821) );
AOI22xp5_ASAP7_75t_L g1791 ( .A1(n_1792), .A2(n_1793), .B1(n_1794), .B2(n_1796), .Y(n_1791) );
INVx1_ASAP7_75t_L g1822 ( .A(n_1804), .Y(n_1822) );
AND2x2_ASAP7_75t_L g1804 ( .A(n_1805), .B(n_1813), .Y(n_1804) );
INVx1_ASAP7_75t_L g1826 ( .A(n_1815), .Y(n_1826) );
INVx1_ASAP7_75t_L g1825 ( .A(n_1817), .Y(n_1825) );
OAI21xp5_ASAP7_75t_L g1820 ( .A1(n_1821), .A2(n_1822), .B(n_1823), .Y(n_1820) );
OAI21xp33_ASAP7_75t_L g1824 ( .A1(n_1823), .A2(n_1825), .B(n_1826), .Y(n_1824) );
CKINVDCx20_ASAP7_75t_R g1827 ( .A(n_1828), .Y(n_1827) );
CKINVDCx20_ASAP7_75t_R g1828 ( .A(n_1829), .Y(n_1828) );
INVx3_ASAP7_75t_L g1829 ( .A(n_1830), .Y(n_1829) );
BUFx3_ASAP7_75t_L g1830 ( .A(n_1831), .Y(n_1830) );
HB1xp67_ASAP7_75t_SL g1834 ( .A(n_1835), .Y(n_1834) );
BUFx3_ASAP7_75t_L g1835 ( .A(n_1836), .Y(n_1835) );
INVxp33_ASAP7_75t_SL g1837 ( .A(n_1838), .Y(n_1837) );
INVx1_ASAP7_75t_L g1885 ( .A(n_1839), .Y(n_1885) );
AND2x2_ASAP7_75t_L g1839 ( .A(n_1840), .B(n_1872), .Y(n_1839) );
AOI21xp5_ASAP7_75t_L g1840 ( .A1(n_1841), .A2(n_1842), .B(n_1862), .Y(n_1840) );
NAND4xp25_ASAP7_75t_L g1842 ( .A(n_1843), .B(n_1846), .C(n_1850), .D(n_1856), .Y(n_1842) );
HB1xp67_ASAP7_75t_L g1886 ( .A(n_1887), .Y(n_1886) );
INVx1_ASAP7_75t_L g1889 ( .A(n_1890), .Y(n_1889) );
endmodule