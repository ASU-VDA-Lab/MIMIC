module fake_jpeg_8156_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx8_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx2_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx11_ASAP7_75t_SL g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_19),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_21),
.Y(n_27)
);

HAxp5_ASAP7_75t_SL g21 ( 
.A(n_9),
.B(n_1),
.CON(n_21),
.SN(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_19),
.A2(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_9),
.B1(n_17),
.B2(n_11),
.Y(n_34)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_34),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_27),
.A2(n_14),
.B1(n_12),
.B2(n_16),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

AOI32xp33_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_8),
.A3(n_18),
.B1(n_25),
.B2(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_28),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_28),
.B1(n_26),
.B2(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_13),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_22),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_47),
.C(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_46),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_33),
.C(n_35),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_40),
.B1(n_31),
.B2(n_17),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g49 ( 
.A(n_47),
.B(n_40),
.Y(n_49)
);

AO221x1_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_32),
.B1(n_11),
.B2(n_37),
.C(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_52),
.Y(n_54)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_53),
.B(n_50),
.Y(n_55)
);

AO21x1_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_54),
.B(n_26),
.Y(n_56)
);

AOI322xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_2),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_1),
.Y(n_57)
);

AOI221xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_5),
.B1(n_7),
.B2(n_22),
.C(n_40),
.Y(n_58)
);


endmodule