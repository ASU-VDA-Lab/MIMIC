module fake_jpeg_32056_n_547 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_547);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_547;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx8_ASAP7_75t_SL g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_57),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_58),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_59),
.Y(n_135)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_63),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_64),
.Y(n_160)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_22),
.B1(n_50),
.B2(n_49),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_69),
.A2(n_21),
.B1(n_49),
.B2(n_47),
.Y(n_125)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_72),
.Y(n_155)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_73),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_29),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_77),
.Y(n_105)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_75),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_78),
.Y(n_166)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_79),
.Y(n_167)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_36),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_90),
.Y(n_111)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_87),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_37),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_92),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

BUFx4f_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_103),
.Y(n_132)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_44),
.Y(n_108)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_104),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_108),
.B(n_139),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_55),
.A2(n_44),
.B1(n_42),
.B2(n_39),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_118),
.A2(n_150),
.B1(n_165),
.B2(n_26),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_99),
.B(n_22),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_123),
.B(n_148),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_125),
.A2(n_145),
.B1(n_27),
.B2(n_28),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_81),
.A2(n_21),
.B1(n_47),
.B2(n_43),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_98),
.A2(n_46),
.B1(n_24),
.B2(n_44),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_53),
.B(n_50),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_64),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_151),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_52),
.A2(n_72),
.B1(n_78),
.B2(n_58),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_77),
.B(n_34),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_L g154 ( 
.A1(n_103),
.A2(n_24),
.B(n_26),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g194 ( 
.A1(n_154),
.A2(n_38),
.B(n_39),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_76),
.B(n_34),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_156),
.B(n_159),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_73),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_71),
.B(n_31),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_162),
.B(n_164),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_63),
.B(n_31),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_59),
.A2(n_25),
.B1(n_43),
.B2(n_27),
.Y(n_165)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_169),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_75),
.B1(n_89),
.B2(n_93),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_170),
.A2(n_172),
.B1(n_183),
.B2(n_185),
.Y(n_272)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_110),
.Y(n_171)
);

INVx13_ASAP7_75t_L g251 ( 
.A(n_171),
.Y(n_251)
);

OA22x2_ASAP7_75t_L g172 ( 
.A1(n_111),
.A2(n_83),
.B1(n_94),
.B2(n_97),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_173),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_174),
.Y(n_247)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_176),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_178),
.A2(n_189),
.B1(n_193),
.B2(n_202),
.Y(n_244)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_126),
.Y(n_179)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_179),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_118),
.B(n_26),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_181),
.B(n_186),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_182),
.Y(n_246)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_184),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_117),
.A2(n_84),
.B1(n_92),
.B2(n_91),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_132),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_129),
.Y(n_188)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_188),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_145),
.A2(n_66),
.B1(n_86),
.B2(n_88),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_190),
.Y(n_267)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_130),
.Y(n_191)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_191),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_119),
.Y(n_192)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_192),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_166),
.A2(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_193)
);

A2O1A1O1Ixp25_ASAP7_75t_L g266 ( 
.A1(n_194),
.A2(n_115),
.B(n_10),
.C(n_11),
.D(n_12),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_107),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_195),
.Y(n_238)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_144),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_196),
.B(n_205),
.Y(n_237)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_114),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_105),
.B(n_30),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_198),
.B(n_201),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_199),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_134),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_200),
.Y(n_258)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_128),
.A2(n_42),
.B(n_39),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_158),
.A2(n_96),
.B1(n_67),
.B2(n_38),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_166),
.A2(n_41),
.B1(n_38),
.B2(n_42),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_203),
.A2(n_206),
.B1(n_210),
.B2(n_211),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_124),
.B(n_41),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_204),
.B(n_216),
.Y(n_269)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_121),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_133),
.A2(n_90),
.B1(n_82),
.B2(n_87),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_130),
.Y(n_207)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_207),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_152),
.A2(n_87),
.B1(n_76),
.B2(n_46),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_153),
.Y(n_209)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_134),
.A2(n_46),
.B1(n_1),
.B2(n_2),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_109),
.A2(n_46),
.B1(n_1),
.B2(n_2),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_213),
.Y(n_240)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_119),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_129),
.A2(n_0),
.B(n_1),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_214),
.Y(n_260)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_138),
.Y(n_215)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_215),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_109),
.B(n_146),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_157),
.B(n_0),
.C(n_3),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_217),
.B(n_9),
.Y(n_276)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_131),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_218),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_135),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_219),
.A2(n_228),
.B1(n_7),
.B2(n_9),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_167),
.B(n_4),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_221),
.Y(n_253)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_114),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_135),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_222),
.A2(n_136),
.B1(n_106),
.B2(n_152),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_146),
.B(n_4),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_223),
.B(n_9),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_122),
.A2(n_5),
.B(n_7),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_225),
.A2(n_122),
.B(n_8),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_160),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_229),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_160),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_227),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_131),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_137),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_241),
.A2(n_225),
.B(n_214),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_248),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_172),
.A2(n_106),
.B1(n_136),
.B2(n_116),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_250),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_L g252 ( 
.A1(n_181),
.A2(n_168),
.B1(n_161),
.B2(n_137),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_252),
.A2(n_188),
.B1(n_190),
.B2(n_207),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_180),
.B(n_224),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_259),
.B(n_263),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_172),
.A2(n_116),
.B1(n_161),
.B2(n_147),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_261),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_187),
.B(n_157),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_264),
.A2(n_268),
.B1(n_185),
.B2(n_206),
.Y(n_303)
);

OR2x6_ASAP7_75t_L g305 ( 
.A(n_266),
.B(n_279),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_230),
.A2(n_168),
.B1(n_147),
.B2(n_155),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_204),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_270),
.B(n_273),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_209),
.Y(n_273)
);

AND2x2_ASAP7_75t_SL g274 ( 
.A(n_186),
.B(n_155),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_216),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_227),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_280),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_276),
.B(n_9),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_172),
.A2(n_141),
.B1(n_10),
.B2(n_11),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_177),
.B(n_141),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_217),
.Y(n_296)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_239),
.Y(n_283)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_283),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_284),
.B(n_298),
.Y(n_343)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_239),
.Y(n_285)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_285),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_183),
.B1(n_169),
.B2(n_171),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_287),
.A2(n_262),
.B1(n_231),
.B2(n_234),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_288),
.A2(n_308),
.B(n_326),
.Y(n_360)
);

OAI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_260),
.A2(n_230),
.B1(n_215),
.B2(n_218),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_289),
.A2(n_290),
.B1(n_303),
.B2(n_234),
.Y(n_335)
);

OAI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_260),
.A2(n_230),
.B1(n_184),
.B2(n_191),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_235),
.Y(n_291)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_291),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_242),
.A2(n_228),
.B(n_199),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_292),
.A2(n_264),
.B(n_232),
.Y(n_332)
);

AND2x2_ASAP7_75t_SL g293 ( 
.A(n_269),
.B(n_223),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_293),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_253),
.B(n_249),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_294),
.Y(n_334)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_235),
.Y(n_295)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_295),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_296),
.B(n_299),
.Y(n_349)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_236),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_297),
.B(n_304),
.Y(n_362)
);

AND2x2_ASAP7_75t_SL g298 ( 
.A(n_269),
.B(n_176),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_233),
.B(n_211),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_247),
.Y(n_300)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_300),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_233),
.B(n_270),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_302),
.B(n_306),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_221),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_237),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_307),
.Y(n_336)
);

O2A1O1Ixp33_ASAP7_75t_L g308 ( 
.A1(n_241),
.A2(n_197),
.B(n_182),
.C(n_174),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_274),
.B(n_173),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_309),
.B(n_318),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_274),
.B(n_222),
.C(n_200),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_310),
.B(n_325),
.C(n_255),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_257),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_312),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_240),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_313),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_316),
.B(n_320),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_236),
.B(n_182),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_317),
.Y(n_352)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_245),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_272),
.A2(n_195),
.B1(n_13),
.B2(n_14),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_319),
.A2(n_322),
.B1(n_323),
.B2(n_258),
.Y(n_340)
);

MAJx2_ASAP7_75t_L g320 ( 
.A(n_276),
.B(n_12),
.C(n_13),
.Y(n_320)
);

INVx3_ASAP7_75t_SL g321 ( 
.A(n_238),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_258),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_252),
.A2(n_244),
.B1(n_242),
.B2(n_256),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_244),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_268),
.B(n_15),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_324),
.B(n_271),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_278),
.B(n_17),
.C(n_18),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_266),
.A2(n_17),
.B(n_18),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_256),
.B(n_17),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_327),
.B(n_328),
.Y(n_371)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_245),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_267),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_330),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_332),
.A2(n_367),
.B(n_300),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_333),
.A2(n_337),
.B1(n_355),
.B2(n_366),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_335),
.B(n_363),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_329),
.A2(n_315),
.B1(n_292),
.B2(n_303),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_322),
.A2(n_231),
.B1(n_273),
.B2(n_238),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_338),
.A2(n_340),
.B1(n_359),
.B2(n_321),
.Y(n_376)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_339),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_307),
.B(n_275),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_341),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_312),
.B(n_255),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_344),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_345),
.B(n_310),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_284),
.B(n_278),
.C(n_271),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_347),
.B(n_354),
.C(n_365),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_353),
.B(n_370),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_302),
.B(n_254),
.C(n_265),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_315),
.A2(n_262),
.B1(n_254),
.B2(n_265),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_301),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_357),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_327),
.A2(n_267),
.B1(n_282),
.B2(n_243),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_301),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_296),
.B(n_251),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_305),
.A2(n_232),
.B1(n_282),
.B2(n_243),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_314),
.A2(n_247),
.B(n_277),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_313),
.B(n_251),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_332),
.A2(n_305),
.B1(n_319),
.B2(n_323),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_373),
.A2(n_388),
.B1(n_399),
.B2(n_403),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_376),
.A2(n_379),
.B1(n_385),
.B2(n_396),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_351),
.B(n_301),
.Y(n_377)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_377),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_342),
.B(n_286),
.Y(n_378)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_378),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_340),
.A2(n_305),
.B1(n_298),
.B2(n_314),
.Y(n_379)
);

NAND3xp33_ASAP7_75t_L g381 ( 
.A(n_336),
.B(n_311),
.C(n_305),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_381),
.B(n_368),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_351),
.B(n_363),
.Y(n_382)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_382),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_357),
.A2(n_288),
.B(n_308),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_384),
.A2(n_390),
.B(n_391),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_338),
.A2(n_305),
.B1(n_298),
.B2(n_324),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_386),
.B(n_365),
.Y(n_411)
);

OAI21xp33_ASAP7_75t_L g387 ( 
.A1(n_342),
.A2(n_305),
.B(n_309),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_387),
.A2(n_393),
.B(n_362),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_337),
.A2(n_299),
.B1(n_306),
.B2(n_304),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_360),
.A2(n_326),
.B(n_283),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_371),
.B(n_293),
.Y(n_392)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_392),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_367),
.A2(n_277),
.B(n_297),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_358),
.Y(n_394)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_394),
.Y(n_429)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_358),
.Y(n_395)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_395),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_362),
.A2(n_293),
.B1(n_285),
.B2(n_318),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_343),
.B(n_316),
.C(n_320),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_398),
.B(n_401),
.Y(n_424)
);

OAI22xp33_ASAP7_75t_SL g399 ( 
.A1(n_353),
.A2(n_335),
.B1(n_366),
.B2(n_356),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_371),
.B(n_291),
.Y(n_400)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_400),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_349),
.B(n_295),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_334),
.A2(n_328),
.B1(n_321),
.B2(n_330),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_402),
.A2(n_331),
.B(n_368),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_349),
.A2(n_246),
.B1(n_325),
.B2(n_356),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_360),
.A2(n_246),
.B1(n_345),
.B2(n_361),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_405),
.A2(n_403),
.B1(n_388),
.B2(n_373),
.Y(n_423)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_406),
.Y(n_437)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_383),
.Y(n_408)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_408),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_383),
.B(n_336),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_410),
.B(n_413),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_411),
.B(n_398),
.C(n_402),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_397),
.B(n_346),
.Y(n_413)
);

NAND2x1_ASAP7_75t_L g451 ( 
.A(n_414),
.B(n_385),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_380),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_415),
.B(n_430),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_397),
.B(n_346),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_416),
.B(n_421),
.Y(n_457)
);

A2O1A1Ixp33_ASAP7_75t_L g417 ( 
.A1(n_377),
.A2(n_361),
.B(n_343),
.C(n_348),
.Y(n_417)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_417),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_386),
.B(n_347),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_420),
.B(n_374),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_378),
.B(n_352),
.Y(n_421)
);

OAI22x1_ASAP7_75t_L g422 ( 
.A1(n_391),
.A2(n_362),
.B1(n_355),
.B2(n_359),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_422),
.A2(n_423),
.B1(n_433),
.B2(n_435),
.Y(n_452)
);

AOI211xp5_ASAP7_75t_L g426 ( 
.A1(n_404),
.A2(n_348),
.B(n_350),
.C(n_354),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_426),
.A2(n_389),
.B1(n_393),
.B2(n_396),
.Y(n_446)
);

A2O1A1O1Ixp25_ASAP7_75t_L g442 ( 
.A1(n_427),
.A2(n_390),
.B(n_384),
.C(n_389),
.D(n_392),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_380),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_382),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_431),
.B(n_400),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_375),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_432),
.B(n_375),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_372),
.A2(n_350),
.B1(n_369),
.B2(n_364),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_425),
.B(n_404),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_438),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_426),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_439),
.B(n_462),
.Y(n_467)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_441),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_442),
.B(n_456),
.Y(n_473)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_443),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_412),
.A2(n_405),
.B1(n_372),
.B2(n_379),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_445),
.A2(n_446),
.B1(n_419),
.B2(n_435),
.Y(n_465)
);

BUFx12_ASAP7_75t_L g447 ( 
.A(n_422),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_447),
.Y(n_466)
);

BUFx12f_ASAP7_75t_SL g448 ( 
.A(n_408),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_448),
.B(n_459),
.Y(n_479)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_451),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_374),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_453),
.B(n_458),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_409),
.B(n_401),
.Y(n_454)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_454),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_409),
.B(n_395),
.Y(n_455)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_455),
.Y(n_477)
);

BUFx5_ASAP7_75t_L g459 ( 
.A(n_414),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_420),
.B(n_394),
.C(n_406),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_460),
.B(n_461),
.C(n_424),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_411),
.B(n_376),
.C(n_331),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_407),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_419),
.A2(n_423),
.B1(n_428),
.B2(n_433),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_463),
.B(n_464),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_418),
.B(n_415),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_465),
.B(n_446),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_468),
.B(n_461),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_438),
.B(n_418),
.Y(n_472)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_472),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_440),
.B(n_436),
.Y(n_474)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_474),
.Y(n_498)
);

XOR2x2_ASAP7_75t_SL g478 ( 
.A(n_451),
.B(n_407),
.Y(n_478)
);

FAx1_ASAP7_75t_SL g493 ( 
.A(n_478),
.B(n_451),
.CI(n_462),
.CON(n_493),
.SN(n_493)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_456),
.B(n_417),
.C(n_430),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_483),
.C(n_484),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_460),
.B(n_428),
.C(n_436),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_453),
.B(n_429),
.C(n_434),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_452),
.A2(n_429),
.B1(n_434),
.B2(n_437),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_485),
.A2(n_445),
.B1(n_464),
.B2(n_455),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_440),
.B(n_437),
.Y(n_486)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_486),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_487),
.B(n_465),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_488),
.A2(n_496),
.B1(n_497),
.B2(n_477),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_470),
.A2(n_439),
.B1(n_457),
.B2(n_449),
.Y(n_489)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_489),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_491),
.B(n_492),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_450),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_493),
.B(n_494),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_467),
.B(n_449),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_472),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_495),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_467),
.A2(n_448),
.B1(n_443),
.B2(n_447),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_466),
.A2(n_447),
.B1(n_444),
.B2(n_442),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_468),
.B(n_458),
.C(n_444),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_500),
.B(n_501),
.C(n_483),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_484),
.B(n_454),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_478),
.A2(n_459),
.B(n_471),
.Y(n_503)
);

FAx1_ASAP7_75t_L g505 ( 
.A(n_503),
.B(n_479),
.CI(n_480),
.CON(n_505),
.SN(n_505)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_504),
.B(n_506),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_505),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_496),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_490),
.A2(n_485),
.B1(n_469),
.B2(n_471),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_507),
.A2(n_513),
.B1(n_488),
.B2(n_477),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_508),
.B(n_509),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_503),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_510),
.A2(n_482),
.B1(n_475),
.B2(n_474),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_491),
.B(n_473),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_514),
.C(n_499),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_495),
.A2(n_498),
.B1(n_502),
.B2(n_469),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_501),
.B(n_473),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_518),
.B(n_514),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_511),
.A2(n_499),
.B(n_500),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_519),
.B(n_520),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_521),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_504),
.B(n_487),
.C(n_476),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_522),
.B(n_526),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_476),
.C(n_497),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_511),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_527),
.B(n_517),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_528),
.B(n_531),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_522),
.B(n_505),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_532),
.B(n_518),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_530),
.A2(n_525),
.B1(n_516),
.B2(n_523),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_534),
.B(n_535),
.C(n_525),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_529),
.B(n_510),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_537),
.A2(n_533),
.B(n_524),
.Y(n_538)
);

AO21x1_ASAP7_75t_L g540 ( 
.A1(n_538),
.A2(n_539),
.B(n_536),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_540),
.A2(n_541),
.B(n_505),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_SL g541 ( 
.A1(n_538),
.A2(n_535),
.B(n_530),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_542),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_543),
.B(n_513),
.C(n_508),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_544),
.B(n_486),
.C(n_507),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_545),
.B(n_475),
.C(n_512),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_546),
.B(n_493),
.Y(n_547)
);


endmodule