module fake_jpeg_9920_n_341 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx10_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_44),
.Y(n_64)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_19),
.B(n_9),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_53),
.B(n_69),
.Y(n_74)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_24),
.B1(n_17),
.B2(n_20),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_57),
.A2(n_20),
.B1(n_17),
.B2(n_24),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_59),
.B(n_46),
.Y(n_96)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_34),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_33),
.Y(n_69)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_52),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_75),
.A2(n_84),
.B1(n_87),
.B2(n_93),
.Y(n_116)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_56),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_53),
.B(n_28),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_85),
.B(n_90),
.Y(n_102)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_94),
.B1(n_61),
.B2(n_49),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_33),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_33),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_97),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_43),
.B(n_61),
.C(n_55),
.Y(n_121)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

NAND2xp33_ASAP7_75t_SL g125 ( 
.A(n_98),
.B(n_46),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_66),
.A2(n_17),
.B1(n_24),
.B2(n_46),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_45),
.B1(n_69),
.B2(n_18),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_60),
.B(n_64),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_105),
.A2(n_117),
.B(n_118),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_64),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_127),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_99),
.A2(n_22),
.B1(n_18),
.B2(n_45),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_109),
.A2(n_119),
.B(n_121),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_67),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_114),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_112),
.A2(n_122),
.B1(n_88),
.B2(n_79),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_60),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_1),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_1),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_92),
.A2(n_41),
.B(n_35),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_61),
.B1(n_43),
.B2(n_49),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_120),
.A2(n_84),
.B1(n_94),
.B2(n_75),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_1),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_124),
.B(n_18),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_1),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g138 ( 
.A(n_125),
.B(n_121),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_41),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_129),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_130),
.B(n_137),
.Y(n_183)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_139),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_106),
.B1(n_126),
.B2(n_115),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_104),
.Y(n_134)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_101),
.A2(n_43),
.B1(n_87),
.B2(n_88),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_135),
.A2(n_144),
.B1(n_131),
.B2(n_146),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_40),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_136),
.B(n_143),
.Y(n_185)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_138),
.A2(n_150),
.B(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_113),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_141),
.A2(n_145),
.B1(n_156),
.B2(n_126),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_108),
.B(n_38),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_101),
.A2(n_112),
.B1(n_105),
.B2(n_125),
.Y(n_144)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_146),
.A2(n_147),
.B1(n_152),
.B2(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_102),
.B(n_40),
.Y(n_148)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_102),
.B(n_98),
.Y(n_151)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

NAND2xp33_ASAP7_75t_SL g153 ( 
.A(n_109),
.B(n_98),
.Y(n_153)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_38),
.C(n_40),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_106),
.C(n_124),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_103),
.B(n_79),
.Y(n_155)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_118),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_117),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_161),
.C(n_163),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_135),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_160),
.B(n_167),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_65),
.B1(n_52),
.B2(n_22),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_117),
.Y(n_163)
);

AND2x4_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_123),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_166),
.B(n_169),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_165),
.A2(n_156),
.B1(n_48),
.B2(n_65),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_149),
.B(n_130),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_133),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_139),
.A2(n_123),
.B1(n_124),
.B2(n_104),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_129),
.C(n_142),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_178),
.C(n_184),
.Y(n_203)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_110),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_132),
.B(n_141),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_173),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_40),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_115),
.B1(n_100),
.B2(n_116),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_179),
.A2(n_154),
.B1(n_150),
.B2(n_148),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_138),
.A2(n_22),
.B1(n_32),
.B2(n_19),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_187),
.B(n_188),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_39),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_136),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_189),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_140),
.A2(n_100),
.B(n_34),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_140),
.A2(n_35),
.B(n_23),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_151),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_39),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_47),
.C(n_35),
.Y(n_212)
);

AND2x6_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_140),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_191),
.A2(n_194),
.B(n_211),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_192),
.A2(n_193),
.B(n_200),
.Y(n_227)
);

AND2x6_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_2),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_198),
.B(n_202),
.Y(n_236)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_205),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_156),
.B(n_145),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_204),
.A2(n_52),
.B(n_72),
.Y(n_239)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_209),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_48),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_212),
.C(n_161),
.Y(n_229)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_210),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

FAx1_ASAP7_75t_SL g216 ( 
.A(n_182),
.B(n_164),
.CI(n_170),
.CON(n_216),
.SN(n_216)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_216),
.B(n_188),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_158),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_218),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_176),
.Y(n_219)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_165),
.Y(n_220)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_163),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_221),
.B(n_223),
.C(n_229),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_184),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_180),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_226),
.Y(n_249)
);

NOR4xp25_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_182),
.C(n_169),
.D(n_187),
.Y(n_225)
);

NAND3xp33_ASAP7_75t_L g264 ( 
.A(n_225),
.B(n_237),
.C(n_247),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_195),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_178),
.C(n_159),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_241),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_232),
.B(n_237),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_234),
.A2(n_202),
.B1(n_196),
.B2(n_218),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_196),
.A2(n_174),
.B(n_181),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_239),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_203),
.B(n_47),
.C(n_71),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_200),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_242),
.B(n_244),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_215),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_197),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_2),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_247),
.A2(n_211),
.B(n_193),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_250),
.B(n_252),
.Y(n_271)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_240),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_253),
.Y(n_284)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_227),
.A2(n_191),
.B(n_216),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_254),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_217),
.Y(n_255)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_194),
.B1(n_216),
.B2(n_212),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_256),
.A2(n_259),
.B1(n_260),
.B2(n_263),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_228),
.A2(n_32),
.B1(n_31),
.B2(n_28),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_246),
.A2(n_31),
.B1(n_26),
.B2(n_21),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_262),
.B(n_267),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_228),
.A2(n_26),
.B1(n_21),
.B2(n_23),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_264),
.B(n_268),
.Y(n_276)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_227),
.A2(n_27),
.B(n_47),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_230),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_269),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_241),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_278),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_231),
.C(n_221),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_277),
.C(n_279),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_229),
.C(n_234),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_223),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_243),
.C(n_233),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_232),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_269),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_266),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_3),
.Y(n_301)
);

A2O1A1Ixp33_ASAP7_75t_L g282 ( 
.A1(n_252),
.A2(n_242),
.B(n_224),
.C(n_238),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_282),
.A2(n_285),
.B1(n_268),
.B2(n_276),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_235),
.C(n_247),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_248),
.C(n_27),
.Y(n_299)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_284),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_290),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_257),
.B1(n_250),
.B2(n_249),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_288),
.A2(n_299),
.B1(n_300),
.B2(n_294),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_271),
.B(n_259),
.CI(n_263),
.CON(n_289),
.SN(n_289)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_289),
.B(n_297),
.Y(n_310)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_286),
.Y(n_290)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_295),
.Y(n_314)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_270),
.Y(n_296)
);

INVxp33_ASAP7_75t_SL g312 ( 
.A(n_296),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_273),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_299),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_29),
.C(n_25),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_25),
.C(n_29),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_5),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_275),
.B1(n_270),
.B2(n_289),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_311),
.C(n_8),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_5),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_304),
.B(n_307),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_308),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_29),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_313),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_294),
.A2(n_25),
.B1(n_6),
.B2(n_7),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_292),
.C(n_25),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_317),
.C(n_324),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_303),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_318),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_7),
.C(n_8),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_319),
.A2(n_310),
.B1(n_311),
.B2(n_16),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_304),
.A2(n_9),
.B1(n_13),
.B2(n_14),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_322),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_13),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_13),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_305),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_328),
.A2(n_331),
.B(n_15),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_15),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_315),
.A2(n_323),
.B(n_324),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_330),
.B(n_14),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_14),
.C(n_15),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_332),
.B(n_333),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_334),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_336),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_327),
.C(n_326),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_327),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_325),
.C(n_331),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_16),
.Y(n_341)
);


endmodule