module real_jpeg_33063_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_455;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_0),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_0),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_1),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_1),
.B(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_1),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_1),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_1),
.B(n_235),
.Y(n_234)
);

AND2x2_ASAP7_75t_SL g275 ( 
.A(n_1),
.B(n_276),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_2),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_2),
.B(n_117),
.Y(n_116)
);

AND2x4_ASAP7_75t_SL g123 ( 
.A(n_2),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_2),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_2),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_2),
.B(n_113),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_2),
.B(n_375),
.Y(n_374)
);

AND2x2_ASAP7_75t_SL g447 ( 
.A(n_2),
.B(n_127),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_3),
.A2(n_19),
.B(n_454),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_3),
.B(n_455),
.Y(n_454)
);

NAND2xp33_ASAP7_75t_R g136 ( 
.A(n_4),
.B(n_137),
.Y(n_136)
);

AND2x4_ASAP7_75t_L g184 ( 
.A(n_4),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_4),
.B(n_154),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_4),
.B(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_4),
.B(n_436),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_5),
.Y(n_455)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

NAND2x1_ASAP7_75t_SL g86 ( 
.A(n_6),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_6),
.B(n_139),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_6),
.A2(n_139),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_6),
.B(n_43),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g258 ( 
.A(n_6),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_6),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_6),
.B(n_127),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_7),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_7),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_7),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_9),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_9),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_10),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_10),
.B(n_131),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_10),
.B(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_10),
.B(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g343 ( 
.A(n_10),
.B(n_344),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_10),
.B(n_95),
.Y(n_398)
);

AND2x4_ASAP7_75t_SL g432 ( 
.A(n_10),
.B(n_433),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_11),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_11),
.Y(n_237)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_11),
.Y(n_283)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_12),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_12),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_12),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_12),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_12),
.B(n_212),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_12),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_12),
.B(n_106),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_12),
.B(n_401),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_14),
.Y(n_132)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_14),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_15),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_15),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_15),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_15),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_15),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_15),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_15),
.B(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_16),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_16),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_17),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_17),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_17),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_17),
.B(n_341),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_17),
.B(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_17),
.B(n_150),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_415),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_358),
.B(n_412),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_314),
.B(n_354),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_191),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_144),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_24),
.B(n_144),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_74),
.C(n_98),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_26),
.A2(n_27),
.B1(n_100),
.B2(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_45),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_28),
.B(n_46),
.C(n_72),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_29),
.B(n_35),
.C(n_39),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_32),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_32),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_38),
.Y(n_203)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_38),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_38),
.Y(n_288)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_44),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_44),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_63),
.B1(n_72),
.B2(n_73),
.Y(n_45)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

MAJx2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_53),
.C(n_58),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_58),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_51),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_52),
.B(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_58),
.A2(n_78),
.B1(n_428),
.B2(n_429),
.Y(n_427)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_62),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_62),
.Y(n_209)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_67),
.B1(n_68),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_64),
.B(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_64),
.A2(n_80),
.B1(n_352),
.B2(n_353),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_64),
.B(n_116),
.Y(n_378)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_71),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_74),
.B(n_194),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_74),
.B(n_194),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.C(n_81),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_75),
.B(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_79),
.B(n_82),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.C(n_92),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_83),
.B(n_86),
.Y(n_245)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_92),
.B(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_119),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_101),
.B(n_134),
.C(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.C(n_114),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_102),
.A2(n_103),
.B1(n_107),
.B2(n_108),
.Y(n_218)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_109),
.B(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_114),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_115),
.A2(n_352),
.B(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_116),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_116),
.A2(n_211),
.B1(n_215),
.B2(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_116),
.B(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_116),
.A2(n_215),
.B1(n_371),
.B2(n_372),
.Y(n_370)
);

MAJx2_ASAP7_75t_L g443 ( 
.A(n_116),
.B(n_374),
.C(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_118),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_134),
.B2(n_143),
.Y(n_119)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_126),
.C(n_129),
.Y(n_157)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_129),
.B1(n_130),
.B2(n_133),
.Y(n_125)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_129),
.B(n_386),
.C(n_387),
.Y(n_437)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2x1_ASAP7_75t_L g379 ( 
.A(n_130),
.B(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

NOR2xp67_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_141),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_141),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_172),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_145),
.B(n_173),
.C(n_175),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_171),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_158),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_147),
.B(n_158),
.C(n_171),
.Y(n_318)
);

XOR2x2_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_156),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_149),
.B(n_152),
.C(n_324),
.Y(n_323)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_155),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_157),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_162),
.B1(n_169),
.B2(n_170),
.Y(n_158)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_159),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_159),
.B(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_161),
.Y(n_385)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_168),
.Y(n_162)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_163),
.B(n_164),
.C(n_169),
.Y(n_349)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

XNOR2x1_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_187),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_176),
.B(n_188),
.C(n_189),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

XOR2x2_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_177),
.B(n_180),
.C(n_184),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_178),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_184),
.Y(n_179)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_188),
.Y(n_190)
);

OAI21x1_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_219),
.B(n_313),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_196),
.B(n_197),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_L g313 ( 
.A(n_193),
.B(n_196),
.C(n_197),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.C(n_216),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_198),
.B(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_200),
.B(n_217),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.C(n_210),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_204),
.B1(n_205),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_202),
.B(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_202),
.B(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_202),
.Y(n_444)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.Y(n_210)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_211),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_248),
.B(n_312),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_246),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_221),
.B(n_246),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.C(n_243),
.Y(n_221)
);

INVxp33_ASAP7_75t_SL g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_223),
.B(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_226),
.A2(n_227),
.B1(n_244),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_233),
.C(n_238),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_229),
.B1(n_233),
.B2(n_234),
.Y(n_253)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_241),
.Y(n_295)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

OAI21x1_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_268),
.B(n_311),
.Y(n_248)
);

NOR2xp67_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_265),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_250),
.B(n_265),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.C(n_257),
.Y(n_250)
);

XNOR2x2_ASAP7_75t_L g307 ( 
.A(n_251),
.B(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_254),
.A2(n_255),
.B1(n_257),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_257),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_262),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_262),
.Y(n_272)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI21x1_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_305),
.B(n_310),
.Y(n_268)
);

OAI21x1_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_291),
.B(n_304),
.Y(n_269)
);

NOR2x1_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_284),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_271),
.B(n_284),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_272),
.B(n_275),
.C(n_277),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_277),
.B2(n_278),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_282),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_289),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_289),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_285),
.B(n_298),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_297),
.B(n_303),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_296),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_296),
.Y(n_303)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp67_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_307),
.Y(n_310)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_315),
.A2(n_356),
.B(n_357),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_316),
.B(n_317),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_318),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_335),
.B2(n_336),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_320),
.Y(n_409)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_334),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_325),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_323),
.Y(n_364)
);

INVxp33_ASAP7_75t_L g365 ( 
.A(n_325),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_331),
.B1(n_332),
.B2(n_333),
.Y(n_325)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_326),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_329),
.B2(n_330),
.Y(n_326)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_327),
.Y(n_330)
);

MAJx2_ASAP7_75t_L g393 ( 
.A(n_328),
.B(n_330),
.C(n_331),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_334),
.Y(n_363)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_336),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_348),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_338),
.B(n_349),
.C(n_350),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_342),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_340),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_340),
.B(n_345),
.C(n_346),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_343),
.A2(n_345),
.B1(n_346),
.B2(n_347),
.Y(n_342)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_343),
.Y(n_346)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_344),
.Y(n_383)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_345),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_406),
.B(n_407),
.Y(n_360)
);

NAND3xp33_ASAP7_75t_L g414 ( 
.A(n_361),
.B(n_406),
.C(n_407),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_366),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_362),
.B(n_366),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_362),
.B(n_419),
.C(n_420),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.C(n_365),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_368),
.B1(n_388),
.B2(n_389),
.Y(n_366)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_367),
.Y(n_420)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_376),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_370),
.B(n_377),
.C(n_379),
.Y(n_439)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_374),
.Y(n_373)
);

XOR2x1_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_379),
.Y(n_376)
);

OAI22x1_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_384),
.B1(n_386),
.B2(n_387),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_381),
.Y(n_386)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_383),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_384),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_389),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_391),
.B1(n_392),
.B2(n_405),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_390),
.Y(n_405)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_394),
.B1(n_403),
.B2(n_404),
.Y(n_392)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_393),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_393),
.B(n_405),
.C(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_394),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_395),
.B(n_397),
.C(n_400),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_398),
.B1(n_399),
.B2(n_400),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_397),
.A2(n_398),
.B1(n_446),
.B2(n_447),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_404),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_410),
.C(n_411),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_R g415 ( 
.A(n_416),
.B(n_450),
.Y(n_415)
);

INVxp33_ASAP7_75t_SL g416 ( 
.A(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_421),
.Y(n_417)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_418),
.Y(n_453)
);

INVxp33_ASAP7_75t_L g452 ( 
.A(n_421),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_424),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_438),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_430),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_428),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_437),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_434),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_441),
.A2(n_442),
.B1(n_448),
.B2(n_449),
.Y(n_440)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_441),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_442),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_445),
.Y(n_442)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVxp33_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);


endmodule