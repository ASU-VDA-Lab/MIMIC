module fake_jpeg_5938_n_180 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx11_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_31),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_0),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_18),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_37),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_27),
.B1(n_18),
.B2(n_26),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_42),
.B1(n_45),
.B2(n_50),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_27),
.B1(n_24),
.B2(n_26),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_29),
.A2(n_24),
.B1(n_15),
.B2(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_31),
.A2(n_23),
.B1(n_21),
.B2(n_17),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_48),
.A2(n_52),
.B1(n_53),
.B2(n_31),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_25),
.B1(n_19),
.B2(n_22),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_22),
.B1(n_28),
.B2(n_21),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_51),
.B(n_0),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_33),
.A2(n_23),
.B1(n_22),
.B2(n_21),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_31),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_56),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_68),
.Y(n_72)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_66),
.Y(n_73)
);

AOI22x1_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_53),
.B1(n_51),
.B2(n_44),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_59),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_30),
.Y(n_62)
);

NOR3xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_43),
.C(n_40),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_58),
.B1(n_62),
.B2(n_44),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_39),
.B(n_32),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_1),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_1),
.Y(n_67)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_70),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_43),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_86),
.B1(n_58),
.B2(n_59),
.Y(n_98)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_52),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_34),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_80),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_41),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_52),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_60),
.C(n_63),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_80),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_40),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_88),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_55),
.B(n_44),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_88),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_96),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_101),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_94),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_72),
.Y(n_113)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_99),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_100),
.B1(n_74),
.B2(n_82),
.Y(n_108)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_89),
.A2(n_56),
.B1(n_47),
.B2(n_65),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_65),
.C(n_38),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_75),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_103),
.B(n_79),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_102),
.C(n_91),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_100),
.B1(n_38),
.B2(n_34),
.Y(n_134)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_93),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_72),
.B(n_77),
.Y(n_114)
);

NOR3xp33_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_122),
.C(n_106),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_94),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_115),
.A2(n_120),
.B1(n_81),
.B2(n_112),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_101),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_119),
.B1(n_81),
.B2(n_85),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_79),
.Y(n_118)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_77),
.B1(n_73),
.B2(n_80),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_99),
.B(n_73),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_130),
.C(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_134),
.B1(n_116),
.B2(n_111),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_106),
.C(n_98),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_111),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_104),
.C(n_92),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_135),
.B(n_2),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_117),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_142),
.C(n_144),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_108),
.B(n_116),
.C(n_120),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_141),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_129),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_81),
.C(n_61),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_146),
.C(n_126),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_10),
.C(n_3),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_154),
.C(n_155),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_141),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_2),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_146),
.Y(n_156)
);

AOI21xp33_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_123),
.B(n_124),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_144),
.C(n_145),
.Y(n_155)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_138),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_155),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_139),
.C(n_4),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_157),
.C(n_158),
.Y(n_167)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_161),
.B(n_4),
.Y(n_165)
);

OAI221xp5_ASAP7_75t_L g168 ( 
.A1(n_162),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_7),
.C(n_8),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_159),
.A2(n_152),
.B1(n_147),
.B2(n_150),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_156),
.B1(n_6),
.B2(n_7),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_168),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_167),
.B(n_5),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_164),
.B1(n_9),
.B2(n_10),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_8),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_172),
.B(n_166),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_173),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_174),
.B(n_175),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_172),
.B(n_170),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_177),
.C(n_8),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_9),
.Y(n_180)
);


endmodule