module fake_jpeg_3830_n_298 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_273;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVxp67_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_9),
.B(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_37),
.B(n_38),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_39),
.B(n_42),
.Y(n_84)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_44),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_7),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_7),
.Y(n_45)
);

NAND2xp33_ASAP7_75t_SL g98 ( 
.A(n_45),
.B(n_47),
.Y(n_98)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_7),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_50),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_52),
.B(n_59),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_38),
.Y(n_53)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_54),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_29),
.B1(n_22),
.B2(n_16),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_55),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_115)
);

CKINVDCx6p67_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_34),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_61),
.B(n_64),
.Y(n_124)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_69),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_34),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_16),
.B1(n_29),
.B2(n_24),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_16),
.B1(n_29),
.B2(n_24),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_24),
.B1(n_23),
.B2(n_22),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_37),
.A2(n_23),
.B1(n_22),
.B2(n_15),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_70),
.A2(n_80),
.B1(n_86),
.B2(n_89),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_25),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_74),
.Y(n_118)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_36),
.B(n_25),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_78),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_36),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_15),
.B1(n_26),
.B2(n_20),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_33),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_88),
.Y(n_126)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_83),
.Y(n_121)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

CKINVDCx12_ASAP7_75t_R g85 ( 
.A(n_41),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_91),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_48),
.A2(n_17),
.B1(n_20),
.B2(n_26),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_39),
.A2(n_17),
.B1(n_33),
.B2(n_14),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_48),
.A2(n_15),
.B1(n_31),
.B2(n_18),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_42),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_28),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_48),
.A2(n_31),
.B1(n_18),
.B2(n_28),
.Y(n_97)
);

XNOR2x1_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

AO22x1_ASAP7_75t_SL g100 ( 
.A1(n_49),
.A2(n_28),
.B1(n_32),
.B2(n_19),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_56),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_57),
.B(n_32),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_125),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_58),
.B(n_84),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_32),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_68),
.Y(n_136)
);

AND2x4_ASAP7_75t_SL g129 ( 
.A(n_100),
.B(n_98),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_128),
.B(n_105),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_130),
.B(n_151),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_124),
.B(n_93),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_131),
.B(n_137),
.Y(n_183)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_134),
.Y(n_182)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_136),
.B(n_146),
.Y(n_190)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_56),
.C(n_70),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_138),
.B(n_147),
.C(n_160),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_129),
.A2(n_72),
.B1(n_79),
.B2(n_87),
.Y(n_139)
);

OAI22x1_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_102),
.B1(n_123),
.B2(n_111),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_72),
.B1(n_87),
.B2(n_79),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_145),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_51),
.B1(n_63),
.B2(n_65),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_142),
.A2(n_151),
.B(n_159),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_117),
.A2(n_80),
.B1(n_67),
.B2(n_89),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_144),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_97),
.B1(n_51),
.B2(n_52),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_28),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_129),
.A2(n_32),
.B1(n_19),
.B2(n_74),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_19),
.B1(n_32),
.B2(n_74),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_148),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_94),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_154),
.Y(n_193)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_150),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_19),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

BUFx24_ASAP7_75t_SL g184 ( 
.A(n_152),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_108),
.B(n_9),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_153),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_94),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

INVxp67_ASAP7_75t_SL g177 ( 
.A(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_62),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_0),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_107),
.A2(n_60),
.B1(n_1),
.B2(n_2),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_110),
.C(n_104),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_162),
.A2(n_101),
.B(n_103),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_163),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_141),
.A2(n_127),
.B1(n_124),
.B2(n_123),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_164),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_168),
.A2(n_176),
.B1(n_174),
.B2(n_194),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_122),
.B(n_118),
.Y(n_169)
);

AOI221xp5_ASAP7_75t_L g204 ( 
.A1(n_169),
.A2(n_154),
.B1(n_151),
.B2(n_160),
.C(n_143),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_118),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_178),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_176),
.A2(n_0),
.B(n_2),
.Y(n_219)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_187),
.Y(n_213)
);

NOR2x1_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_141),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_181),
.B(n_112),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_120),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_142),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_159),
.B(n_103),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_188),
.B(n_10),
.Y(n_217)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_112),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_130),
.B(n_104),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_130),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_147),
.C(n_162),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_138),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_198),
.C(n_199),
.Y(n_229)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_181),
.C(n_190),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_216),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_201),
.Y(n_235)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_205),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_137),
.Y(n_203)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_144),
.Y(n_206)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_140),
.C(n_145),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_210),
.C(n_215),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_209),
.A2(n_170),
.B1(n_175),
.B2(n_173),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_101),
.C(n_163),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_212),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_161),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_190),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_220),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_218),
.B(n_173),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_219),
.B(n_164),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_116),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_214),
.A2(n_165),
.B1(n_191),
.B2(n_174),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_223),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_166),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_226),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_228),
.B(n_213),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_218),
.A2(n_165),
.B1(n_168),
.B2(n_180),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_230),
.A2(n_232),
.B1(n_207),
.B2(n_202),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_214),
.A2(n_192),
.B1(n_187),
.B2(n_190),
.Y(n_232)
);

OAI322xp33_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_172),
.A3(n_195),
.B1(n_188),
.B2(n_183),
.C1(n_167),
.C2(n_184),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_213),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_170),
.Y(n_236)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_236),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_237),
.A2(n_238),
.B(n_200),
.Y(n_250)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_240),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_197),
.C(n_199),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_243),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_209),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_244),
.A2(n_238),
.B(n_222),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_252),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_246),
.Y(n_257)
);

AO221x1_ASAP7_75t_L g248 ( 
.A1(n_239),
.A2(n_177),
.B1(n_179),
.B2(n_186),
.C(n_171),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_248),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_250),
.B(n_255),
.Y(n_259)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_198),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_256),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_254),
.A2(n_230),
.B1(n_223),
.B2(n_232),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_205),
.C(n_208),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_231),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_266),
.Y(n_274)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_222),
.B(n_208),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_267),
.B(n_256),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_242),
.B(n_224),
.Y(n_261)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

XOR2x1_ASAP7_75t_SL g265 ( 
.A(n_250),
.B(n_234),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_265),
.A2(n_225),
.B1(n_198),
.B2(n_245),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_242),
.B(n_239),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_268),
.B(n_167),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_269),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_259),
.A2(n_249),
.B1(n_225),
.B2(n_252),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_270),
.A2(n_273),
.B(n_275),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_265),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_276),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_241),
.C(n_243),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_267),
.B(n_175),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_253),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_240),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_278),
.B(n_237),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_280),
.A2(n_282),
.B(n_227),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_270),
.B(n_251),
.Y(n_282)
);

AOI322xp5_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_260),
.A3(n_258),
.B1(n_262),
.B2(n_228),
.C1(n_255),
.C2(n_264),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_285),
.C(n_275),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_289),
.C(n_277),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_287),
.B(n_288),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_246),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_279),
.A2(n_271),
.B(n_273),
.Y(n_289)
);

AOI21x1_ASAP7_75t_SL g290 ( 
.A1(n_281),
.A2(n_240),
.B(n_227),
.Y(n_290)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_219),
.C(n_240),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_283),
.B1(n_257),
.B2(n_251),
.Y(n_291)
);

AO21x1_ASAP7_75t_L g296 ( 
.A1(n_291),
.A2(n_292),
.B(n_221),
.Y(n_296)
);

OAI322xp33_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_217),
.A3(n_263),
.B1(n_216),
.B2(n_221),
.C1(n_5),
.C2(n_8),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_296),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_293),
.Y(n_298)
);


endmodule