module fake_jpeg_27178_n_225 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_36),
.Y(n_45)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_38),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_1),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_18),
.B1(n_31),
.B2(n_26),
.Y(n_47)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_27),
.B1(n_31),
.B2(n_26),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_40),
.B1(n_36),
.B2(n_18),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_27),
.B1(n_42),
.B2(n_35),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_56),
.B1(n_58),
.B2(n_40),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_16),
.Y(n_75)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_17),
.B1(n_25),
.B2(n_33),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_17),
.B1(n_25),
.B2(n_33),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_59),
.A2(n_73),
.B1(n_41),
.B2(n_20),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_64),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_44),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_63),
.B(n_65),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_34),
.B(n_38),
.C(n_39),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_57),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_39),
.B(n_38),
.C(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_67),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_30),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_22),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_72),
.B(n_74),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_16),
.B1(n_21),
.B2(n_22),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_38),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_75),
.B(n_77),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_29),
.Y(n_100)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_19),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_34),
.B1(n_36),
.B2(n_19),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_79),
.A2(n_80),
.B1(n_53),
.B2(n_50),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_24),
.B1(n_23),
.B2(n_29),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_82),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_52),
.B(n_20),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_20),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_50),
.Y(n_105)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_54),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_86),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_105),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_78),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_52),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_77),
.Y(n_121)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_97),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_106),
.B1(n_79),
.B2(n_75),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_64),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_101),
.Y(n_125)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_15),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_107),
.Y(n_124)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

CKINVDCx10_ASAP7_75t_R g108 ( 
.A(n_67),
.Y(n_108)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_41),
.B(n_24),
.C(n_23),
.Y(n_133)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_111),
.B(n_54),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_120),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_63),
.B(n_65),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_115),
.A2(n_131),
.B(n_117),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_69),
.Y(n_116)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

AO21x1_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_75),
.B(n_76),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_4),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_118),
.A2(n_133),
.B1(n_98),
.B2(n_97),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_74),
.C(n_65),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_126),
.C(n_91),
.Y(n_144)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_92),
.B1(n_99),
.B2(n_95),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_132),
.B1(n_98),
.B2(n_108),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_89),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_123),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_86),
.C(n_60),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_89),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_130),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_60),
.Y(n_129)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_24),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_83),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_135),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_80),
.B1(n_71),
.B2(n_81),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_134),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_96),
.B(n_23),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_104),
.B1(n_93),
.B2(n_103),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_136),
.A2(n_152),
.B1(n_155),
.B2(n_127),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_147),
.B1(n_151),
.B2(n_114),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_111),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_143),
.B(n_127),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_156),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_107),
.C(n_91),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_149),
.C(n_133),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_71),
.C(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_121),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_150),
.B(n_5),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_118),
.A2(n_110),
.B1(n_29),
.B2(n_41),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_157),
.B(n_133),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_3),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_154),
.A2(n_122),
.A3(n_112),
.B1(n_125),
.B2(n_132),
.C1(n_133),
.C2(n_114),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_152),
.Y(n_186)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_120),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_161),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_164),
.B1(n_165),
.B2(n_170),
.Y(n_179)
);

BUFx12_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_163),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_141),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_166),
.A2(n_173),
.B1(n_148),
.B2(n_127),
.Y(n_183)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_6),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_138),
.Y(n_172)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_155),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_156),
.C(n_136),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_165),
.A2(n_147),
.B1(n_145),
.B2(n_150),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_180),
.B1(n_175),
.B2(n_170),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_166),
.A2(n_145),
.B1(n_151),
.B2(n_144),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_159),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_162),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_187),
.B(n_171),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_179),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_193),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_191),
.A2(n_198),
.B1(n_182),
.B2(n_178),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_186),
.Y(n_205)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_159),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_177),
.B(n_160),
.Y(n_195)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_196),
.A2(n_197),
.B1(n_181),
.B2(n_188),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_173),
.B1(n_169),
.B2(n_163),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_198),
.Y(n_199)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_180),
.C(n_185),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_201),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_203),
.A2(n_189),
.B1(n_193),
.B2(n_182),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_206),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_212),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_204),
.A2(n_189),
.B1(n_184),
.B2(n_163),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_199),
.Y(n_214)
);

BUFx24_ASAP7_75t_SL g212 ( 
.A(n_206),
.Y(n_212)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_214),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_202),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_216),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_200),
.C(n_209),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_6),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_7),
.C(n_8),
.Y(n_220)
);

AOI322xp5_ASAP7_75t_L g222 ( 
.A1(n_220),
.A2(n_221),
.A3(n_218),
.B1(n_15),
.B2(n_219),
.C1(n_8),
.C2(n_9),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_217),
.A2(n_10),
.B(n_12),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_222),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_8),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_9),
.Y(n_225)
);


endmodule