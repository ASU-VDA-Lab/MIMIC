module real_jpeg_11891_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx10_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_3),
.A2(n_30),
.B1(n_32),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_3),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_4),
.A2(n_20),
.B1(n_23),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_4),
.A2(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_7),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_7),
.A2(n_22),
.B1(n_56),
.B2(n_57),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_7),
.A2(n_22),
.B1(n_30),
.B2(n_32),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_8),
.B(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_8),
.B(n_56),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_SL g75 ( 
.A1(n_8),
.A2(n_55),
.B(n_56),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_8),
.B(n_26),
.C(n_32),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_8),
.A2(n_20),
.B1(n_23),
.B2(n_86),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_8),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_9),
.A2(n_30),
.B1(n_32),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_10),
.A2(n_30),
.B1(n_32),
.B2(n_47),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_10),
.A2(n_20),
.B1(n_23),
.B2(n_47),
.Y(n_70)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_78),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_77),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_51),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_16),
.B(n_51),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_36),
.C(n_42),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_17),
.A2(n_18),
.B1(n_36),
.B2(n_37),
.Y(n_105)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_24),
.B1(n_33),
.B2(n_34),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_19),
.A2(n_24),
.B1(n_33),
.B2(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_SL g23 ( 
.A(n_20),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g39 ( 
.A1(n_20),
.A2(n_23),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_20),
.A2(n_41),
.B(n_54),
.C(n_59),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_20),
.B(n_83),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND3xp33_ASAP7_75t_SL g59 ( 
.A(n_23),
.B(n_40),
.C(n_57),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_24),
.A2(n_33),
.B1(n_34),
.B2(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_29),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_27),
.B1(n_30),
.B2(n_32),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_29),
.B(n_86),
.Y(n_99)
);

INVx5_ASAP7_75t_SL g32 ( 
.A(n_30),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_30),
.B(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_39),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_40),
.A2(n_41),
.B1(n_56),
.B2(n_57),
.Y(n_74)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_42),
.B(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B(n_48),
.Y(n_42)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_43),
.A2(n_44),
.B1(n_89),
.B2(n_96),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_44),
.B(n_86),
.Y(n_94)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_45),
.A2(n_61),
.B1(n_88),
.B2(n_90),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_46),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_61),
.B(n_62),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_67),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_52)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_102),
.B(n_106),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_91),
.B(n_101),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_87),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_87),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_84),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_97),
.B(n_100),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_99),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_104),
.Y(n_106)
);


endmodule