module fake_netlist_1_8109_n_38 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
BUFx2_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_3), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_10), .Y(n_13) );
INVx4_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
NOR2xp33_ASAP7_75t_R g15 ( .A(n_1), .B(n_9), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_6), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_1), .Y(n_17) );
AOI22xp5_ASAP7_75t_L g18 ( .A1(n_11), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_18) );
OAI22xp5_ASAP7_75t_L g19 ( .A1(n_11), .A2(n_0), .B1(n_2), .B2(n_4), .Y(n_19) );
AOI22xp5_ASAP7_75t_L g20 ( .A1(n_11), .A2(n_5), .B1(n_7), .B2(n_8), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_14), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_17), .B(n_5), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
CKINVDCx16_ASAP7_75t_R g24 ( .A(n_22), .Y(n_24) );
AOI22xp33_ASAP7_75t_L g25 ( .A1(n_19), .A2(n_17), .B1(n_14), .B2(n_12), .Y(n_25) );
AO21x1_ASAP7_75t_L g26 ( .A1(n_18), .A2(n_14), .B(n_13), .Y(n_26) );
NOR2xp33_ASAP7_75t_R g27 ( .A(n_24), .B(n_12), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_23), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_24), .B(n_14), .Y(n_29) );
NAND4xp75_ASAP7_75t_L g30 ( .A(n_29), .B(n_26), .C(n_20), .D(n_13), .Y(n_30) );
OAI221xp5_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_25), .B1(n_16), .B2(n_23), .C(n_14), .Y(n_31) );
OAI22xp33_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_27), .B1(n_28), .B2(n_26), .Y(n_32) );
NOR2xp33_ASAP7_75t_SL g33 ( .A(n_30), .B(n_15), .Y(n_33) );
INVx1_ASAP7_75t_SL g34 ( .A(n_33), .Y(n_34) );
HB1xp67_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
BUFx6f_ASAP7_75t_L g36 ( .A(n_33), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_34), .Y(n_37) );
AOI22xp33_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_36), .B1(n_35), .B2(n_7), .Y(n_38) );
endmodule