module fake_jpeg_5864_n_217 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_217);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_217;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_SL g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_32),
.B(n_35),
.Y(n_71)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_36),
.B(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_37),
.B(n_38),
.Y(n_76)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_39),
.A2(n_47),
.B1(n_27),
.B2(n_21),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_40),
.B(n_42),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_5),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_46),
.B(n_31),
.Y(n_49)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_49),
.B(n_62),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_36),
.C(n_41),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_53),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_31),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_51),
.B(n_55),
.Y(n_104)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_20),
.C(n_29),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_30),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_56),
.Y(n_89)
);

AO22x1_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_18),
.B1(n_19),
.B2(n_23),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_57),
.A2(n_60),
.B1(n_81),
.B2(n_25),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_58),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_27),
.B1(n_19),
.B2(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_67),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_38),
.A2(n_27),
.B1(n_29),
.B2(n_24),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_28),
.B1(n_6),
.B2(n_8),
.Y(n_101)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_70),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_32),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_78),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_33),
.B(n_30),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_39),
.A2(n_24),
.B1(n_16),
.B2(n_26),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_39),
.B(n_16),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_3),
.Y(n_113)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_86),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_41),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_41),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_88),
.B(n_8),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_28),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_80),
.C(n_58),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_25),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_84),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_48),
.B1(n_75),
.B2(n_87),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_101),
.A2(n_11),
.B1(n_13),
.B2(n_103),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_63),
.A2(n_5),
.B(n_13),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_102),
.A2(n_110),
.B(n_10),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_63),
.A2(n_28),
.B1(n_1),
.B2(n_2),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_103),
.A2(n_4),
.B1(n_10),
.B2(n_11),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_113),
.B(n_76),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_117),
.B(n_120),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_119),
.B(n_131),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_79),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_71),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_124),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_79),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_122),
.B(n_125),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_91),
.A2(n_48),
.B1(n_54),
.B2(n_75),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_58),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_73),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_56),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_143),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_133),
.C(n_141),
.Y(n_144)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_143),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_100),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_130),
.B(n_132),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_0),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_64),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_93),
.A2(n_56),
.B(n_69),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_80),
.B1(n_59),
.B2(n_69),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_1),
.Y(n_137)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_4),
.Y(n_138)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

NOR3xp33_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_142),
.C(n_102),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_112),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_140),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_94),
.A2(n_11),
.B1(n_13),
.B2(n_96),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_94),
.A2(n_96),
.B1(n_112),
.B2(n_92),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_147),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_140),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_163),
.B(n_117),
.Y(n_170)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_156),
.B(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_116),
.Y(n_159)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_116),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_160),
.Y(n_171)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_161),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_105),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_131),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_121),
.C(n_128),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_168),
.C(n_169),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_120),
.B(n_133),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_167),
.A2(n_170),
.B(n_174),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_152),
.B(n_130),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_126),
.C(n_134),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_119),
.C(n_132),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_148),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_155),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_118),
.B1(n_142),
.B2(n_136),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_175),
.A2(n_179),
.B1(n_157),
.B2(n_153),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_153),
.A2(n_92),
.B1(n_138),
.B2(n_111),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_177),
.A2(n_145),
.B1(n_164),
.B2(n_148),
.Y(n_189)
);

FAx1_ASAP7_75t_SL g178 ( 
.A(n_163),
.B(n_135),
.CI(n_106),
.CON(n_178),
.SN(n_178)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_178),
.B(n_161),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_151),
.A2(n_111),
.B1(n_97),
.B2(n_99),
.Y(n_179)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

AOI221xp5_ASAP7_75t_L g183 ( 
.A1(n_167),
.A2(n_162),
.B1(n_165),
.B2(n_154),
.C(n_150),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_180),
.Y(n_198)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_185),
.A2(n_188),
.B(n_191),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_175),
.A2(n_151),
.B1(n_158),
.B2(n_149),
.Y(n_187)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_189),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_166),
.C(n_168),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

AOI321xp33_ASAP7_75t_L g202 ( 
.A1(n_196),
.A2(n_198),
.A3(n_185),
.B1(n_191),
.B2(n_186),
.C(n_184),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_190),
.C(n_172),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_169),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_193),
.B(n_188),
.Y(n_201)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_202),
.A2(n_206),
.B1(n_171),
.B2(n_178),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_200),
.B(n_197),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_204),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_194),
.A2(n_192),
.B(n_176),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

AO22x1_ASAP7_75t_L g208 ( 
.A1(n_205),
.A2(n_200),
.B1(n_197),
.B2(n_195),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_198),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_199),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_212),
.C(n_213),
.Y(n_214)
);

MAJx2_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_208),
.C(n_196),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_214),
.Y(n_215)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_213),
.B(n_181),
.Y(n_216)
);

BUFx24_ASAP7_75t_SL g217 ( 
.A(n_216),
.Y(n_217)
);


endmodule