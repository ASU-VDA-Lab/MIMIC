module fake_jpeg_22097_n_345 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx8_ASAP7_75t_SL g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_9),
.B(n_14),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_38),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_40),
.B(n_44),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_15),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_30),
.B1(n_17),
.B2(n_35),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_50),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_18),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_20),
.B1(n_28),
.B2(n_26),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_53),
.A2(n_59),
.B1(n_21),
.B2(n_34),
.Y(n_97)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_55),
.B(n_66),
.Y(n_119)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_20),
.B1(n_28),
.B2(n_26),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_28),
.B1(n_21),
.B2(n_34),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_61),
.A2(n_27),
.B1(n_31),
.B2(n_23),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_64),
.Y(n_111)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_74),
.B(n_35),
.Y(n_95)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_45),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_83),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_37),
.B1(n_47),
.B2(n_21),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_86),
.A2(n_97),
.B1(n_104),
.B2(n_68),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_67),
.B(n_50),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_87),
.B(n_92),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_37),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_89),
.B(n_90),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_37),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_46),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_47),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_94),
.B(n_100),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_95),
.A2(n_15),
.B(n_13),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_47),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_109),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_41),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_60),
.A2(n_17),
.B1(n_31),
.B2(n_27),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_101),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_54),
.B(n_25),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_103),
.B(n_110),
.Y(n_149)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_53),
.B(n_14),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_41),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_65),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_60),
.A2(n_51),
.B1(n_48),
.B2(n_44),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_114),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_59),
.B(n_41),
.Y(n_115)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_71),
.A2(n_82),
.B(n_79),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_116),
.A2(n_57),
.B(n_78),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_55),
.A2(n_32),
.B1(n_24),
.B2(n_29),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_122),
.B1(n_78),
.B2(n_70),
.Y(n_135)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_121),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_57),
.A2(n_43),
.B1(n_39),
.B2(n_41),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_94),
.C(n_108),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_127),
.C(n_138),
.Y(n_162)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_139),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_41),
.C(n_40),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_90),
.B(n_43),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_128),
.B(n_137),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_129),
.B(n_12),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_131),
.A2(n_105),
.B(n_85),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_102),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_132),
.Y(n_173)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_140),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_117),
.B1(n_120),
.B2(n_84),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_43),
.C(n_69),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_148),
.Y(n_166)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_150),
.Y(n_172)
);

NAND2xp33_ASAP7_75t_SL g144 ( 
.A(n_96),
.B(n_1),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_152),
.B(n_91),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_93),
.B(n_70),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_151),
.A2(n_122),
.B1(n_23),
.B2(n_24),
.Y(n_170)
);

NOR2x1_ASAP7_75t_L g152 ( 
.A(n_95),
.B(n_1),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_110),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_155),
.B(n_156),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_88),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_158),
.B(n_159),
.Y(n_210)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_88),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_161),
.B(n_163),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_143),
.B(n_97),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_131),
.A2(n_68),
.B1(n_99),
.B2(n_120),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_174),
.B1(n_181),
.B2(n_183),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_SL g218 ( 
.A(n_165),
.B(n_171),
.C(n_8),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_102),
.Y(n_167)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_168),
.A2(n_170),
.B1(n_147),
.B2(n_106),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_169),
.Y(n_192)
);

A2O1A1O1Ixp25_ASAP7_75t_L g171 ( 
.A1(n_128),
.A2(n_23),
.B(n_24),
.C(n_32),
.D(n_29),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_138),
.A2(n_99),
.B1(n_84),
.B2(n_109),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_175),
.B(n_186),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_111),
.Y(n_176)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_123),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_177),
.B(n_179),
.Y(n_198)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_127),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_141),
.A2(n_118),
.B1(n_85),
.B2(n_105),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g183 ( 
.A1(n_141),
.A2(n_18),
.B1(n_29),
.B2(n_32),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_184),
.A2(n_185),
.B(n_2),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_136),
.A2(n_18),
.B(n_106),
.C(n_98),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_111),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_125),
.B(n_98),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_140),
.B(n_145),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_137),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_189),
.B(n_196),
.C(n_209),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_190),
.A2(n_191),
.B1(n_218),
.B2(n_183),
.Y(n_246)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_152),
.B1(n_144),
.B2(n_125),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_160),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_194),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_159),
.A2(n_152),
.B1(n_136),
.B2(n_149),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_195),
.A2(n_199),
.B(n_203),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_187),
.B(n_162),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_197),
.A2(n_200),
.B(n_205),
.Y(n_228)
);

O2A1O1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_124),
.B(n_107),
.C(n_4),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_184),
.A2(n_2),
.B(n_3),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_179),
.A2(n_139),
.B1(n_12),
.B2(n_11),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_163),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_206),
.A2(n_168),
.B1(n_175),
.B2(n_178),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_156),
.A2(n_4),
.B(n_5),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_207),
.A2(n_172),
.B(n_154),
.C(n_185),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_11),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_11),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_217),
.C(n_181),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_188),
.A2(n_4),
.B(n_6),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_213),
.A2(n_215),
.B1(n_178),
.B2(n_157),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_177),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_215)
);

MAJx2_ASAP7_75t_L g216 ( 
.A(n_165),
.B(n_7),
.C(n_8),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_216),
.B(n_220),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_8),
.C(n_9),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_155),
.B(n_9),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_172),
.Y(n_222)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_224),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_225),
.B(n_191),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_154),
.Y(n_227)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_227),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_173),
.Y(n_232)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_197),
.B(n_219),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_233),
.A2(n_237),
.B(n_238),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_234),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_213),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_235),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_207),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_171),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_192),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_206),
.B(n_158),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_244),
.B(n_211),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_200),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_245),
.B1(n_246),
.B2(n_215),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_10),
.C(n_237),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_166),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_193),
.A2(n_205),
.B1(n_195),
.B2(n_190),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_248),
.B1(n_199),
.B2(n_191),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_204),
.A2(n_221),
.B1(n_202),
.B2(n_217),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_251),
.A2(n_253),
.B1(n_265),
.B2(n_266),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_196),
.C(n_189),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_263),
.C(n_271),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_247),
.A2(n_201),
.B1(n_202),
.B2(n_216),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_259),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_261),
.A2(n_240),
.B(n_222),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_209),
.C(n_157),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_264),
.B(n_228),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_242),
.A2(n_214),
.B1(n_191),
.B2(n_182),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_233),
.A2(n_183),
.B1(n_180),
.B2(n_169),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_180),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_229),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_169),
.B1(n_9),
.B2(n_10),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_269),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_245),
.Y(n_276)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_281),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_250),
.A2(n_223),
.B1(n_234),
.B2(n_235),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_278),
.A2(n_287),
.B1(n_265),
.B2(n_225),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_251),
.A2(n_241),
.B1(n_225),
.B2(n_228),
.Y(n_279)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_279),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_255),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_257),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_229),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_243),
.C(n_229),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_263),
.C(n_271),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_227),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_286),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_266),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_270),
.A2(n_232),
.B1(n_241),
.B2(n_231),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_253),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_289),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_259),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_290),
.B(n_261),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_293),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_295),
.C(n_304),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_268),
.C(n_267),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_279),
.B(n_255),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_302),
.Y(n_314)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_280),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_239),
.Y(n_303)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_303),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_231),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_313),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_275),
.C(n_272),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_315),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_300),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_309),
.A2(n_311),
.B(n_290),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_298),
.A2(n_276),
.B(n_288),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_274),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_305),
.A2(n_287),
.B1(n_278),
.B2(n_277),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_283),
.C(n_285),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_317),
.A2(n_292),
.B(n_262),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_302),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_243),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_304),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_320),
.C(n_307),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_326),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_296),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_325),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_310),
.A2(n_291),
.B(n_249),
.Y(n_325)
);

NOR2x1_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_249),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_327),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_328),
.B(n_332),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_316),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_308),
.C(n_307),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_333),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_327),
.C(n_312),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_334),
.A2(n_314),
.B1(n_254),
.B2(n_312),
.Y(n_336)
);

AND3x1_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_324),
.C(n_325),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_336),
.C(n_293),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_337),
.A2(n_330),
.B(n_329),
.Y(n_339)
);

AOI321xp33_ASAP7_75t_L g341 ( 
.A1(n_339),
.A2(n_340),
.A3(n_338),
.B1(n_337),
.B2(n_273),
.C(n_244),
.Y(n_341)
);

OAI321xp33_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_273),
.A3(n_245),
.B1(n_282),
.B2(n_260),
.C(n_238),
.Y(n_342)
);

AOI21x1_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_260),
.B(n_238),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_10),
.B(n_331),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_344),
.Y(n_345)
);


endmodule