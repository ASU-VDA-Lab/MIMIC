module real_aes_16916_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_1034;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_1499;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_286;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1403;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_0), .A2(n_209), .B1(n_449), .B2(n_795), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_0), .A2(n_71), .B1(n_353), .B2(n_815), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_1), .A2(n_3), .B1(n_1158), .B2(n_1161), .Y(n_1171) );
INVx1_ASAP7_75t_L g706 ( .A(n_2), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_2), .A2(n_101), .B1(n_449), .B2(n_726), .Y(n_725) );
XNOR2xp5_ASAP7_75t_L g1362 ( .A(n_3), .B(n_1363), .Y(n_1362) );
AOI22xp33_ASAP7_75t_L g1458 ( .A1(n_3), .A2(n_1459), .B1(n_1494), .B2(n_1499), .Y(n_1458) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_4), .A2(n_121), .B1(n_356), .B2(n_361), .Y(n_355) );
AOI22xp33_ASAP7_75t_SL g445 ( .A1(n_4), .A2(n_127), .B1(n_446), .B2(n_448), .Y(n_445) );
INVx1_ASAP7_75t_L g1020 ( .A(n_5), .Y(n_1020) );
XNOR2x2_ASAP7_75t_L g570 ( .A(n_6), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g804 ( .A(n_7), .Y(n_804) );
OAI22xp33_ASAP7_75t_L g823 ( .A1(n_7), .A2(n_72), .B1(n_376), .B2(n_824), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_8), .A2(n_221), .B1(n_449), .B2(n_795), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_8), .A2(n_267), .B1(n_353), .B2(n_636), .Y(n_856) );
INVx1_ASAP7_75t_L g295 ( .A(n_9), .Y(n_295) );
AND2x2_ASAP7_75t_L g402 ( .A(n_9), .B(n_232), .Y(n_402) );
AND2x2_ASAP7_75t_L g428 ( .A(n_9), .B(n_429), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g894 ( .A(n_9), .B(n_305), .Y(n_894) );
AOI22xp33_ASAP7_75t_SL g344 ( .A1(n_10), .A2(n_165), .B1(n_345), .B2(n_352), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_10), .A2(n_17), .B1(n_432), .B2(n_436), .C(n_443), .Y(n_431) );
OAI22xp33_ASAP7_75t_L g589 ( .A1(n_11), .A2(n_48), .B1(n_387), .B2(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g610 ( .A(n_11), .Y(n_610) );
AOI22xp33_ASAP7_75t_SL g1067 ( .A1(n_12), .A2(n_194), .B1(n_514), .B2(n_708), .Y(n_1067) );
INVxp67_ASAP7_75t_SL g1072 ( .A(n_12), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g1474 ( .A1(n_13), .A2(n_79), .B1(n_449), .B2(n_736), .Y(n_1474) );
AOI22xp33_ASAP7_75t_L g1489 ( .A1(n_13), .A2(n_137), .B1(n_353), .B2(n_514), .Y(n_1489) );
INVx2_ASAP7_75t_L g1154 ( .A(n_14), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_14), .B(n_102), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_14), .B(n_1160), .Y(n_1162) );
CKINVDCx5p33_ASAP7_75t_R g645 ( .A(n_15), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_16), .A2(n_91), .B1(n_418), .B2(n_694), .Y(n_850) );
AOI22xp33_ASAP7_75t_SL g372 ( .A1(n_17), .A2(n_33), .B1(n_373), .B2(n_374), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_18), .A2(n_250), .B1(n_584), .B2(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1086 ( .A(n_18), .Y(n_1086) );
INVx1_ASAP7_75t_L g330 ( .A(n_19), .Y(n_330) );
OAI22xp33_ASAP7_75t_L g375 ( .A1(n_20), .A2(n_214), .B1(n_376), .B2(n_387), .Y(n_375) );
INVx1_ASAP7_75t_L g456 ( .A(n_20), .Y(n_456) );
XNOR2xp5_ASAP7_75t_L g739 ( .A(n_21), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g651 ( .A(n_22), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_23), .A2(n_51), .B1(n_356), .B2(n_1030), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_23), .A2(n_279), .B1(n_601), .B2(n_673), .Y(n_1040) );
AOI22xp5_ASAP7_75t_L g1187 ( .A1(n_24), .A2(n_237), .B1(n_1158), .B2(n_1161), .Y(n_1187) );
INVx1_ASAP7_75t_L g730 ( .A(n_25), .Y(n_730) );
AOI22xp33_ASAP7_75t_SL g707 ( .A1(n_26), .A2(n_77), .B1(n_514), .B2(n_708), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_26), .A2(n_277), .B1(n_433), .B2(n_443), .C(n_657), .Y(n_724) );
INVx1_ASAP7_75t_L g729 ( .A(n_27), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_28), .A2(n_163), .B1(n_1106), .B2(n_1108), .Y(n_1105) );
AOI221xp5_ASAP7_75t_L g1128 ( .A1(n_28), .A2(n_230), .B1(n_436), .B2(n_759), .C(n_1129), .Y(n_1128) );
XNOR2xp5_ASAP7_75t_L g1460 ( .A(n_29), .B(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1018 ( .A(n_30), .Y(n_1018) );
OAI221xp5_ASAP7_75t_L g1042 ( .A1(n_30), .A2(n_145), .B1(n_613), .B2(n_614), .C(n_1043), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_31), .A2(n_96), .B1(n_418), .B2(n_694), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_32), .A2(n_277), .B1(n_514), .B2(n_708), .Y(n_717) );
AOI22xp33_ASAP7_75t_SL g735 ( .A1(n_32), .A2(n_77), .B1(n_673), .B2(n_736), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_33), .A2(n_461), .B(n_465), .C(n_477), .Y(n_460) );
AOI22xp33_ASAP7_75t_SL g578 ( .A1(n_34), .A2(n_160), .B1(n_514), .B2(n_579), .Y(n_578) );
INVxp67_ASAP7_75t_SL g616 ( .A(n_34), .Y(n_616) );
AOI22xp33_ASAP7_75t_SL g1027 ( .A1(n_35), .A2(n_279), .B1(n_361), .B2(n_1028), .Y(n_1027) );
AOI221xp5_ASAP7_75t_L g1046 ( .A1(n_35), .A2(n_51), .B1(n_523), .B2(n_838), .C(n_1047), .Y(n_1046) );
AOI22xp5_ASAP7_75t_L g1176 ( .A1(n_36), .A2(n_270), .B1(n_1151), .B2(n_1177), .Y(n_1176) );
XNOR2xp5_ASAP7_75t_L g828 ( .A(n_37), .B(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g1120 ( .A(n_38), .Y(n_1120) );
INVx1_ASAP7_75t_L g789 ( .A(n_39), .Y(n_789) );
INVx1_ASAP7_75t_L g1381 ( .A(n_40), .Y(n_1381) );
INVx1_ASAP7_75t_L g1095 ( .A(n_41), .Y(n_1095) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_42), .A2(n_64), .B1(n_408), .B2(n_418), .Y(n_407) );
OAI211xp5_ASAP7_75t_L g422 ( .A1(n_42), .A2(n_423), .B(n_430), .C(n_451), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g1180 ( .A1(n_43), .A2(n_248), .B1(n_1158), .B2(n_1161), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_44), .A2(n_170), .B1(n_449), .B2(n_801), .Y(n_844) );
AOI22xp33_ASAP7_75t_SL g858 ( .A1(n_44), .A2(n_122), .B1(n_390), .B2(n_505), .Y(n_858) );
INVx1_ASAP7_75t_L g954 ( .A(n_45), .Y(n_954) );
AO22x1_ASAP7_75t_L g1184 ( .A1(n_45), .A2(n_62), .B1(n_1151), .B2(n_1166), .Y(n_1184) );
OAI22xp33_ASAP7_75t_L g1421 ( .A1(n_46), .A2(n_168), .B1(n_1422), .B2(n_1423), .Y(n_1421) );
OAI22xp5_ASAP7_75t_L g1429 ( .A1(n_46), .A2(n_117), .B1(n_1430), .B2(n_1431), .Y(n_1429) );
XNOR2x2_ASAP7_75t_L g311 ( .A(n_47), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g609 ( .A(n_48), .Y(n_609) );
AOI21xp33_ASAP7_75t_L g758 ( .A1(n_49), .A2(n_657), .B(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g767 ( .A(n_49), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_50), .A2(n_230), .B1(n_1030), .B2(n_1106), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_50), .A2(n_163), .B1(n_446), .B2(n_448), .Y(n_1124) );
INVx1_ASAP7_75t_L g1372 ( .A(n_52), .Y(n_1372) );
INVx1_ASAP7_75t_L g337 ( .A(n_53), .Y(n_337) );
INVx1_ASAP7_75t_L g351 ( .A(n_53), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_54), .A2(n_126), .B1(n_514), .B2(n_579), .Y(n_1111) );
AOI221xp5_ASAP7_75t_L g1122 ( .A1(n_54), .A2(n_75), .B1(n_443), .B2(n_604), .C(n_1123), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_55), .A2(n_80), .B1(n_509), .B2(n_513), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g521 ( .A1(n_55), .A2(n_255), .B1(n_522), .B2(n_523), .C(n_524), .Y(n_521) );
INVx1_ASAP7_75t_L g692 ( .A(n_56), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_57), .A2(n_204), .B1(n_446), .B2(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g768 ( .A(n_57), .Y(n_768) );
INVx1_ASAP7_75t_L g1410 ( .A(n_58), .Y(n_1410) );
OAI211xp5_ASAP7_75t_L g1434 ( .A1(n_58), .A2(n_1435), .B(n_1436), .C(n_1438), .Y(n_1434) );
AOI221xp5_ASAP7_75t_L g1472 ( .A1(n_59), .A2(n_133), .B1(n_657), .B2(n_838), .C(n_1473), .Y(n_1472) );
AOI22xp33_ASAP7_75t_SL g1490 ( .A1(n_59), .A2(n_200), .B1(n_390), .B2(n_505), .Y(n_1490) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_60), .A2(n_127), .B1(n_361), .B2(n_364), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g466 ( .A1(n_60), .A2(n_121), .B1(n_467), .B2(n_470), .C(n_473), .Y(n_466) );
INVx1_ASAP7_75t_L g1022 ( .A(n_61), .Y(n_1022) );
INVx1_ASAP7_75t_L g288 ( .A(n_63), .Y(n_288) );
INVx2_ASAP7_75t_L g327 ( .A(n_65), .Y(n_327) );
AOI221xp5_ASAP7_75t_L g744 ( .A1(n_66), .A2(n_239), .B1(n_443), .B2(n_745), .C(n_746), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_66), .A2(n_276), .B1(n_353), .B2(n_514), .Y(n_769) );
INVx1_ASAP7_75t_L g1385 ( .A(n_67), .Y(n_1385) );
CKINVDCx5p33_ASAP7_75t_R g1013 ( .A(n_68), .Y(n_1013) );
INVx1_ASAP7_75t_L g1057 ( .A(n_69), .Y(n_1057) );
OAI222xp33_ASAP7_75t_L g1082 ( .A1(n_69), .A2(n_247), .B1(n_536), .B2(n_558), .C1(n_1083), .C2(n_1087), .Y(n_1082) );
AOI22xp5_ASAP7_75t_L g1181 ( .A1(n_70), .A2(n_185), .B1(n_1151), .B2(n_1166), .Y(n_1181) );
AOI221xp5_ASAP7_75t_L g798 ( .A1(n_71), .A2(n_202), .B1(n_433), .B2(n_443), .C(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g803 ( .A(n_72), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_73), .A2(n_142), .B1(n_505), .B2(n_507), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_73), .A2(n_144), .B1(n_526), .B2(n_529), .Y(n_525) );
AO221x2_ASAP7_75t_L g1223 ( .A1(n_74), .A2(n_219), .B1(n_1158), .B2(n_1161), .C(n_1224), .Y(n_1223) );
AOI22xp33_ASAP7_75t_SL g1104 ( .A1(n_75), .A2(n_224), .B1(n_374), .B2(n_514), .Y(n_1104) );
AOI22xp33_ASAP7_75t_SL g635 ( .A1(n_76), .A2(n_190), .B1(n_579), .B2(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_76), .A2(n_241), .B1(n_446), .B2(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g1094 ( .A(n_78), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g1492 ( .A1(n_79), .A2(n_275), .B1(n_514), .B2(n_1493), .Y(n_1492) );
INVx1_ASAP7_75t_L g556 ( .A(n_80), .Y(n_556) );
INVx1_ASAP7_75t_L g980 ( .A(n_81), .Y(n_980) );
AOI221xp5_ASAP7_75t_L g993 ( .A1(n_81), .A2(n_130), .B1(n_657), .B2(n_745), .C(n_994), .Y(n_993) );
AOI21xp33_ASAP7_75t_L g793 ( .A1(n_82), .A2(n_746), .B(n_759), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_82), .A2(n_179), .B1(n_505), .B2(n_817), .Y(n_816) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_83), .A2(n_217), .B1(n_408), .B2(n_596), .Y(n_1014) );
OAI211xp5_ASAP7_75t_L g1033 ( .A1(n_83), .A2(n_519), .B(n_1034), .C(n_1041), .Y(n_1033) );
OAI211xp5_ASAP7_75t_L g785 ( .A1(n_84), .A2(n_613), .B(n_786), .C(n_790), .Y(n_785) );
INVx1_ASAP7_75t_L g812 ( .A(n_84), .Y(n_812) );
INVx1_ASAP7_75t_L g500 ( .A(n_85), .Y(n_500) );
OAI211xp5_ASAP7_75t_L g518 ( .A1(n_85), .A2(n_519), .B(n_520), .C(n_531), .Y(n_518) );
INVx1_ASAP7_75t_L g1100 ( .A(n_86), .Y(n_1100) );
CKINVDCx5p33_ASAP7_75t_R g1407 ( .A(n_87), .Y(n_1407) );
INVx1_ASAP7_75t_L g833 ( .A(n_88), .Y(n_833) );
INVx1_ASAP7_75t_L g1059 ( .A(n_89), .Y(n_1059) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_90), .A2(n_132), .B1(n_408), .B2(n_596), .Y(n_595) );
OAI211xp5_ASAP7_75t_L g840 ( .A1(n_91), .A2(n_519), .B(n_841), .C(n_845), .Y(n_840) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_92), .Y(n_565) );
INVx1_ASAP7_75t_L g892 ( .A(n_93), .Y(n_892) );
AOI221xp5_ASAP7_75t_L g919 ( .A1(n_93), .A2(n_222), .B1(n_774), .B2(n_920), .C(n_922), .Y(n_919) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_94), .Y(n_290) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_94), .B(n_288), .Y(n_1152) );
AOI22xp33_ASAP7_75t_SL g638 ( .A1(n_95), .A2(n_280), .B1(n_639), .B2(n_641), .Y(n_638) );
AOI21xp33_ASAP7_75t_L g669 ( .A1(n_95), .A2(n_548), .B(n_670), .Y(n_669) );
OAI211xp5_ASAP7_75t_SL g796 ( .A1(n_96), .A2(n_423), .B(n_797), .C(n_802), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_97), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_98), .A2(n_266), .B1(n_387), .B2(n_590), .Y(n_652) );
INVx1_ASAP7_75t_L g660 ( .A(n_98), .Y(n_660) );
CKINVDCx5p33_ASAP7_75t_R g713 ( .A(n_99), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_100), .A2(n_128), .B1(n_505), .B2(n_581), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_100), .A2(n_176), .B1(n_548), .B2(n_621), .C(n_623), .Y(n_620) );
INVx1_ASAP7_75t_L g716 ( .A(n_101), .Y(n_716) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_102), .B(n_1154), .Y(n_1153) );
INVx1_ASAP7_75t_L g1160 ( .A(n_102), .Y(n_1160) );
OAI22xp33_ASAP7_75t_L g944 ( .A1(n_103), .A2(n_238), .B1(n_945), .B2(n_948), .Y(n_944) );
INVxp67_ASAP7_75t_SL g951 ( .A(n_103), .Y(n_951) );
INVx1_ASAP7_75t_L g1380 ( .A(n_104), .Y(n_1380) );
AOI22xp5_ASAP7_75t_L g1479 ( .A1(n_105), .A2(n_200), .B1(n_736), .B2(n_749), .Y(n_1479) );
AOI22xp5_ASAP7_75t_L g1491 ( .A1(n_105), .A2(n_133), .B1(n_505), .B2(n_1064), .Y(n_1491) );
OAI21xp33_ASAP7_75t_L g560 ( .A1(n_106), .A2(n_561), .B(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g1477 ( .A(n_107), .Y(n_1477) );
INVx1_ASAP7_75t_L g1482 ( .A(n_108), .Y(n_1482) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_109), .A2(n_255), .B1(n_507), .B2(n_509), .Y(n_506) );
INVx1_ASAP7_75t_L g546 ( .A(n_109), .Y(n_546) );
INVx1_ASAP7_75t_L g701 ( .A(n_110), .Y(n_701) );
AOI21xp33_ASAP7_75t_L g734 ( .A1(n_110), .A2(n_548), .B(n_657), .Y(n_734) );
INVx2_ASAP7_75t_L g329 ( .A(n_111), .Y(n_329) );
INVx1_ASAP7_75t_L g371 ( .A(n_111), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_111), .B(n_327), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_112), .A2(n_158), .B1(n_362), .B2(n_925), .Y(n_984) );
INVx1_ASAP7_75t_L g995 ( .A(n_112), .Y(n_995) );
AOI21xp33_ASAP7_75t_L g836 ( .A1(n_113), .A2(n_837), .B(n_838), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_113), .A2(n_170), .B1(n_505), .B2(n_817), .Y(n_857) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_114), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g1170 ( .A1(n_115), .A2(n_216), .B1(n_1151), .B2(n_1166), .Y(n_1170) );
INVx1_ASAP7_75t_L g576 ( .A(n_116), .Y(n_576) );
OAI221xp5_ASAP7_75t_L g612 ( .A1(n_116), .A2(n_196), .B1(n_613), .B2(n_614), .C(n_615), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g1414 ( .A1(n_117), .A2(n_125), .B1(n_1415), .B2(n_1418), .Y(n_1414) );
INVx1_ASAP7_75t_L g904 ( .A(n_118), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g868 ( .A1(n_119), .A2(n_150), .B1(n_869), .B2(n_870), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_119), .A2(n_208), .B1(n_505), .B2(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g1079 ( .A(n_120), .Y(n_1079) );
INVxp67_ASAP7_75t_SL g835 ( .A(n_122), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_123), .A2(n_233), .B1(n_596), .B2(n_694), .Y(n_693) );
OAI211xp5_ASAP7_75t_L g722 ( .A1(n_123), .A2(n_519), .B(n_723), .C(n_728), .Y(n_722) );
INVx1_ASAP7_75t_L g849 ( .A(n_124), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g1445 ( .A1(n_125), .A2(n_168), .B1(n_1446), .B2(n_1448), .Y(n_1445) );
AOI22xp33_ASAP7_75t_L g1127 ( .A1(n_126), .A2(n_224), .B1(n_448), .B2(n_736), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_128), .A2(n_180), .B1(n_601), .B2(n_602), .Y(n_600) );
XNOR2xp5_ASAP7_75t_L g955 ( .A(n_129), .B(n_956), .Y(n_955) );
AOI221xp5_ASAP7_75t_L g973 ( .A1(n_130), .A2(n_252), .B1(n_354), .B2(n_974), .C(n_975), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_131), .A2(n_162), .B1(n_583), .B2(n_1066), .Y(n_1065) );
INVx1_ASAP7_75t_L g1085 ( .A(n_131), .Y(n_1085) );
OAI211xp5_ASAP7_75t_L g598 ( .A1(n_132), .A2(n_423), .B(n_599), .C(n_608), .Y(n_598) );
AOI22xp33_ASAP7_75t_SL g1061 ( .A1(n_134), .A2(n_210), .B1(n_514), .B2(n_1062), .Y(n_1061) );
INVxp67_ASAP7_75t_SL g1088 ( .A(n_134), .Y(n_1088) );
INVx1_ASAP7_75t_L g847 ( .A(n_135), .Y(n_847) );
OAI22xp33_ASAP7_75t_L g860 ( .A1(n_135), .A2(n_186), .B1(n_590), .B2(n_824), .Y(n_860) );
AOI22xp33_ASAP7_75t_SL g1031 ( .A1(n_136), .A2(n_153), .B1(n_374), .B2(n_815), .Y(n_1031) );
AOI221xp5_ASAP7_75t_L g1035 ( .A1(n_136), .A2(n_184), .B1(n_524), .B2(n_1036), .C(n_1038), .Y(n_1035) );
AOI221xp5_ASAP7_75t_L g1478 ( .A1(n_137), .A2(n_275), .B1(n_438), .B2(n_607), .C(n_745), .Y(n_1478) );
INVx1_ASAP7_75t_L g1481 ( .A(n_138), .Y(n_1481) );
INVx1_ASAP7_75t_L g752 ( .A(n_139), .Y(n_752) );
INVxp67_ASAP7_75t_SL g633 ( .A(n_140), .Y(n_633) );
OAI211xp5_ASAP7_75t_L g654 ( .A1(n_140), .A2(n_519), .B(n_655), .C(n_659), .Y(n_654) );
AOI22xp33_ASAP7_75t_SL g642 ( .A1(n_141), .A2(n_260), .B1(n_639), .B2(n_641), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_141), .A2(n_280), .B1(n_449), .B2(n_527), .Y(n_658) );
INVx1_ASAP7_75t_L g541 ( .A(n_142), .Y(n_541) );
OAI21xp5_ASAP7_75t_L g1483 ( .A1(n_143), .A2(n_694), .B(n_1484), .Y(n_1483) );
AOI22xp33_ASAP7_75t_SL g503 ( .A1(n_144), .A2(n_147), .B1(n_504), .B2(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g1017 ( .A(n_145), .Y(n_1017) );
OAI22xp33_ASAP7_75t_L g963 ( .A1(n_146), .A2(n_273), .B1(n_945), .B2(n_948), .Y(n_963) );
INVxp33_ASAP7_75t_SL g1004 ( .A(n_146), .Y(n_1004) );
INVx1_ASAP7_75t_L g550 ( .A(n_147), .Y(n_550) );
AOI22xp33_ASAP7_75t_SL g760 ( .A1(n_148), .A2(n_276), .B1(n_425), .B2(n_736), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_148), .A2(n_239), .B1(n_514), .B2(n_774), .Y(n_773) );
OAI21xp5_ASAP7_75t_L g1091 ( .A1(n_149), .A2(n_694), .B(n_1092), .Y(n_1091) );
AOI22xp33_ASAP7_75t_SL g916 ( .A1(n_150), .A2(n_263), .B1(n_641), .B2(n_917), .Y(n_916) );
AO22x1_ASAP7_75t_L g1185 ( .A1(n_151), .A2(n_235), .B1(n_1158), .B2(n_1161), .Y(n_1185) );
INVx1_ASAP7_75t_L g751 ( .A(n_152), .Y(n_751) );
INVxp67_ASAP7_75t_SL g1045 ( .A(n_153), .Y(n_1045) );
INVx1_ASAP7_75t_L g1078 ( .A(n_154), .Y(n_1078) );
INVx1_ASAP7_75t_L g630 ( .A(n_155), .Y(n_630) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_155), .A2(n_157), .B1(n_536), .B2(n_558), .C(n_664), .Y(n_663) );
BUFx3_ASAP7_75t_L g321 ( .A(n_156), .Y(n_321) );
INVx1_ASAP7_75t_L g631 ( .A(n_157), .Y(n_631) );
INVx1_ASAP7_75t_L g989 ( .A(n_158), .Y(n_989) );
CKINVDCx5p33_ASAP7_75t_R g966 ( .A(n_159), .Y(n_966) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_160), .A2(n_244), .B1(n_604), .B2(n_605), .C(n_607), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_161), .A2(n_241), .B1(n_504), .B2(n_579), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_161), .A2(n_190), .B1(n_433), .B2(n_443), .C(n_657), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g1075 ( .A1(n_162), .A2(n_250), .B1(n_449), .B2(n_1076), .Y(n_1075) );
INVx1_ASAP7_75t_L g970 ( .A(n_164), .Y(n_970) );
AOI221xp5_ASAP7_75t_L g987 ( .A1(n_164), .A2(n_203), .B1(n_657), .B2(n_745), .C(n_988), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_165), .B(n_476), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g842 ( .A1(n_166), .A2(n_267), .B1(n_433), .B2(n_524), .C(n_843), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_166), .A2(n_221), .B1(n_374), .B2(n_504), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g1167 ( .A1(n_167), .A2(n_181), .B1(n_1158), .B2(n_1161), .Y(n_1167) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_169), .Y(n_302) );
INVx1_ASAP7_75t_L g958 ( .A(n_171), .Y(n_958) );
INVx1_ASAP7_75t_L g1384 ( .A(n_172), .Y(n_1384) );
CKINVDCx20_ASAP7_75t_R g1113 ( .A(n_173), .Y(n_1113) );
CKINVDCx5p33_ASAP7_75t_R g967 ( .A(n_174), .Y(n_967) );
AOI221xp5_ASAP7_75t_L g887 ( .A1(n_175), .A2(n_208), .B1(n_870), .B2(n_888), .C(n_890), .Y(n_887) );
AOI221xp5_ASAP7_75t_L g918 ( .A1(n_175), .A2(n_215), .B1(n_514), .B2(n_579), .C(n_821), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_176), .A2(n_180), .B1(n_581), .B2(n_584), .Y(n_580) );
OAI211xp5_ASAP7_75t_L g1402 ( .A1(n_177), .A2(n_1084), .B(n_1403), .C(n_1406), .Y(n_1402) );
INVx1_ASAP7_75t_L g1442 ( .A(n_177), .Y(n_1442) );
AOI22xp33_ASAP7_75t_SL g1024 ( .A1(n_178), .A2(n_184), .B1(n_514), .B2(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g1044 ( .A(n_178), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_179), .A2(n_257), .B1(n_449), .B2(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g978 ( .A(n_182), .Y(n_978) );
INVx1_ASAP7_75t_L g1465 ( .A(n_183), .Y(n_1465) );
INVx1_ASAP7_75t_L g846 ( .A(n_186), .Y(n_846) );
AOI22xp5_ASAP7_75t_L g1188 ( .A1(n_187), .A2(n_249), .B1(n_1151), .B2(n_1166), .Y(n_1188) );
INVx1_ASAP7_75t_L g1374 ( .A(n_188), .Y(n_1374) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_189), .Y(n_594) );
OAI221xp5_ASAP7_75t_L g753 ( .A1(n_191), .A2(n_242), .B1(n_536), .B2(n_558), .C(n_754), .Y(n_753) );
OAI22xp33_ASAP7_75t_L g775 ( .A1(n_191), .A2(n_242), .B1(n_496), .B2(n_719), .Y(n_775) );
INVx1_ASAP7_75t_L g497 ( .A(n_192), .Y(n_497) );
OAI222xp33_ASAP7_75t_L g535 ( .A1(n_192), .A2(n_274), .B1(n_536), .B2(n_537), .C1(n_549), .C2(n_557), .Y(n_535) );
INVx1_ASAP7_75t_L g566 ( .A(n_193), .Y(n_566) );
INVxp67_ASAP7_75t_SL g1090 ( .A(n_194), .Y(n_1090) );
CKINVDCx5p33_ASAP7_75t_R g1101 ( .A(n_195), .Y(n_1101) );
INVx1_ASAP7_75t_L g575 ( .A(n_196), .Y(n_575) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_197), .Y(n_534) );
INVx1_ASAP7_75t_L g1118 ( .A(n_198), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1165 ( .A1(n_199), .A2(n_245), .B1(n_1151), .B2(n_1166), .Y(n_1165) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_201), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_202), .A2(n_209), .B1(n_374), .B2(n_815), .Y(n_818) );
AOI21xp33_ASAP7_75t_L g983 ( .A1(n_203), .A2(n_366), .B(n_922), .Y(n_983) );
INVx1_ASAP7_75t_L g772 ( .A(n_204), .Y(n_772) );
INVx1_ASAP7_75t_L g1114 ( .A(n_205), .Y(n_1114) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_206), .Y(n_406) );
INVxp67_ASAP7_75t_SL g791 ( .A(n_207), .Y(n_791) );
AOI22xp33_ASAP7_75t_SL g822 ( .A1(n_207), .A2(n_257), .B1(n_361), .B2(n_390), .Y(n_822) );
AOI21xp33_ASAP7_75t_L g1074 ( .A1(n_210), .A2(n_607), .B(n_837), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_211), .B(n_626), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_211), .A2(n_647), .B1(n_648), .B2(n_679), .Y(n_646) );
INVx1_ASAP7_75t_L g681 ( .A(n_211), .Y(n_681) );
AO22x1_ASAP7_75t_L g1150 ( .A1(n_212), .A2(n_236), .B1(n_1151), .B2(n_1155), .Y(n_1150) );
OA22x2_ASAP7_75t_L g782 ( .A1(n_213), .A2(n_783), .B1(n_826), .B2(n_827), .Y(n_782) );
CKINVDCx16_ASAP7_75t_R g826 ( .A(n_213), .Y(n_826) );
INVx1_ASAP7_75t_L g452 ( .A(n_214), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g871 ( .A1(n_215), .A2(n_222), .B1(n_872), .B2(n_874), .C(n_876), .Y(n_871) );
INVx1_ASAP7_75t_L g316 ( .A(n_218), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_220), .A2(n_278), .B1(n_596), .B2(n_694), .Y(n_778) );
INVxp67_ASAP7_75t_SL g907 ( .A(n_223), .Y(n_907) );
OAI221xp5_ASAP7_75t_L g936 ( .A1(n_223), .A2(n_227), .B1(n_937), .B2(n_939), .C(n_941), .Y(n_936) );
INVx1_ASAP7_75t_L g777 ( .A(n_225), .Y(n_777) );
OAI211xp5_ASAP7_75t_SL g964 ( .A1(n_226), .A2(n_934), .B(n_941), .C(n_965), .Y(n_964) );
INVx1_ASAP7_75t_L g1000 ( .A(n_226), .Y(n_1000) );
OAI221xp5_ASAP7_75t_L g878 ( .A1(n_227), .A2(n_240), .B1(n_879), .B2(n_884), .C(n_885), .Y(n_878) );
OAI211xp5_ASAP7_75t_L g831 ( .A1(n_228), .A2(n_613), .B(n_832), .C(n_834), .Y(n_831) );
INVx1_ASAP7_75t_L g854 ( .A(n_228), .Y(n_854) );
AOI22xp5_ASAP7_75t_L g1175 ( .A1(n_229), .A2(n_256), .B1(n_1158), .B2(n_1161), .Y(n_1175) );
INVx1_ASAP7_75t_L g1470 ( .A(n_231), .Y(n_1470) );
BUFx3_ASAP7_75t_L g305 ( .A(n_232), .Y(n_305) );
INVx1_ASAP7_75t_L g429 ( .A(n_232), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g1226 ( .A(n_234), .Y(n_1226) );
XOR2x2_ASAP7_75t_L g1010 ( .A(n_236), .B(n_1011), .Y(n_1010) );
INVxp67_ASAP7_75t_SL g899 ( .A(n_238), .Y(n_899) );
OAI22xp5_ASAP7_75t_L g926 ( .A1(n_240), .A2(n_243), .B1(n_927), .B2(n_930), .Y(n_926) );
INVxp67_ASAP7_75t_SL g909 ( .A(n_243), .Y(n_909) );
AOI22xp33_ASAP7_75t_SL g587 ( .A1(n_244), .A2(n_262), .B1(n_514), .B2(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g324 ( .A(n_246), .Y(n_324) );
INVx2_ASAP7_75t_L g343 ( .A(n_246), .Y(n_343) );
INVx1_ASAP7_75t_L g385 ( .A(n_246), .Y(n_385) );
INVx1_ASAP7_75t_L g1056 ( .A(n_247), .Y(n_1056) );
INVx1_ASAP7_75t_L g1368 ( .A(n_251), .Y(n_1368) );
INVx1_ASAP7_75t_L g990 ( .A(n_252), .Y(n_990) );
INVx1_ASAP7_75t_L g1471 ( .A(n_253), .Y(n_1471) );
AO22x1_ASAP7_75t_L g1157 ( .A1(n_254), .A2(n_271), .B1(n_1158), .B2(n_1161), .Y(n_1157) );
INVx1_ASAP7_75t_L g806 ( .A(n_258), .Y(n_806) );
INVx1_ASAP7_75t_L g1136 ( .A(n_259), .Y(n_1136) );
INVx1_ASAP7_75t_L g665 ( .A(n_260), .Y(n_665) );
OAI21xp5_ASAP7_75t_L g1134 ( .A1(n_261), .A2(n_408), .B(n_1135), .Y(n_1134) );
INVxp67_ASAP7_75t_SL g619 ( .A(n_262), .Y(n_619) );
INVx1_ASAP7_75t_L g891 ( .A(n_263), .Y(n_891) );
INVx1_ASAP7_75t_L g1375 ( .A(n_264), .Y(n_1375) );
OAI22xp33_ASAP7_75t_SL g718 ( .A1(n_265), .A2(n_272), .B1(n_496), .B2(n_719), .Y(n_718) );
OAI221xp5_ASAP7_75t_L g731 ( .A1(n_265), .A2(n_272), .B1(n_558), .B2(n_613), .C(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g662 ( .A(n_266), .Y(n_662) );
XNOR2xp5_ASAP7_75t_L g689 ( .A(n_268), .B(n_690), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g972 ( .A(n_269), .Y(n_972) );
INVxp67_ASAP7_75t_SL g961 ( .A(n_273), .Y(n_961) );
INVx1_ASAP7_75t_L g494 ( .A(n_274), .Y(n_494) );
OAI211xp5_ASAP7_75t_L g742 ( .A1(n_278), .A2(n_519), .B(n_743), .C(n_750), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_306), .B(n_1143), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_291), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g1457 ( .A(n_285), .B(n_294), .Y(n_1457) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g1498 ( .A(n_287), .B(n_290), .Y(n_1498) );
INVx1_ASAP7_75t_L g1501 ( .A(n_287), .Y(n_1501) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g1504 ( .A(n_290), .B(n_1501), .Y(n_1504) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_296), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g1426 ( .A(n_294), .B(n_1427), .Y(n_1426) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_L g444 ( .A(n_295), .B(n_305), .Y(n_444) );
AND2x4_ASAP7_75t_L g474 ( .A(n_295), .B(n_304), .Y(n_474) );
AND2x4_ASAP7_75t_SL g1456 ( .A(n_296), .B(n_1457), .Y(n_1456) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x6_ASAP7_75t_L g297 ( .A(n_298), .B(n_303), .Y(n_297) );
INVxp67_ASAP7_75t_L g476 ( .A(n_298), .Y(n_476) );
OR2x6_ASAP7_75t_L g1416 ( .A(n_298), .B(n_1417), .Y(n_1416) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx3_ASAP7_75t_L g552 ( .A(n_299), .Y(n_552) );
BUFx4f_ASAP7_75t_L g1371 ( .A(n_299), .Y(n_1371) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx2_ASAP7_75t_L g404 ( .A(n_301), .Y(n_404) );
INVx1_ASAP7_75t_L g412 ( .A(n_301), .Y(n_412) );
INVx2_ASAP7_75t_L g427 ( .A(n_301), .Y(n_427) );
AND2x2_ASAP7_75t_L g435 ( .A(n_301), .B(n_302), .Y(n_435) );
AND2x2_ASAP7_75t_L g441 ( .A(n_301), .B(n_442), .Y(n_441) );
NAND2x1_ASAP7_75t_L g540 ( .A(n_301), .B(n_302), .Y(n_540) );
INVx1_ASAP7_75t_L g405 ( .A(n_302), .Y(n_405) );
AND2x2_ASAP7_75t_L g426 ( .A(n_302), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g442 ( .A(n_302), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_302), .B(n_427), .Y(n_464) );
BUFx2_ASAP7_75t_L g480 ( .A(n_302), .Y(n_480) );
OR2x2_ASAP7_75t_L g545 ( .A(n_302), .B(n_404), .Y(n_545) );
OR2x6_ASAP7_75t_L g1422 ( .A(n_303), .B(n_552), .Y(n_1422) );
INVxp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g1405 ( .A(n_304), .Y(n_1405) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx2_ASAP7_75t_L g1409 ( .A(n_305), .Y(n_1409) );
AND2x4_ASAP7_75t_L g1413 ( .A(n_305), .B(n_411), .Y(n_1413) );
OAI22xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_1008), .B1(n_1141), .B2(n_1142), .Y(n_306) );
INVx1_ASAP7_75t_L g1141 ( .A(n_307), .Y(n_1141) );
XNOR2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_684), .Y(n_307) );
XOR2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_489), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND3xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_393), .C(n_421), .Y(n_312) );
NOR3xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_375), .C(n_391), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_338), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B1(n_330), .B2(n_331), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_316), .A2(n_330), .B1(n_478), .B2(n_482), .Y(n_477) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_322), .Y(n_317) );
NAND2x1_ASAP7_75t_L g496 ( .A(n_318), .B(n_322), .Y(n_496) );
AND2x4_ASAP7_75t_SL g811 ( .A(n_318), .B(n_322), .Y(n_811) );
AND2x6_ASAP7_75t_L g938 ( .A(n_318), .B(n_325), .Y(n_938) );
INVx3_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x4_ASAP7_75t_L g362 ( .A(n_320), .B(n_335), .Y(n_362) );
NAND2x1p5_ASAP7_75t_L g416 ( .A(n_320), .B(n_417), .Y(n_416) );
BUFx2_ASAP7_75t_L g1441 ( .A(n_320), .Y(n_1441) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g348 ( .A(n_321), .Y(n_348) );
AND2x4_ASAP7_75t_L g354 ( .A(n_321), .B(n_336), .Y(n_354) );
OR2x2_ASAP7_75t_L g379 ( .A(n_321), .B(n_350), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_321), .B(n_337), .Y(n_399) );
AND2x4_ASAP7_75t_L g331 ( .A(n_322), .B(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g392 ( .A(n_322), .B(n_353), .Y(n_392) );
AND2x4_ASAP7_75t_SL g720 ( .A(n_322), .B(n_332), .Y(n_720) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
OR2x2_ASAP7_75t_L g400 ( .A(n_323), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g897 ( .A(n_323), .Y(n_897) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g370 ( .A(n_324), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_324), .B(n_428), .Y(n_902) );
NAND2x1p5_ASAP7_75t_L g419 ( .A(n_325), .B(n_347), .Y(n_419) );
AND2x2_ASAP7_75t_L g940 ( .A(n_325), .B(n_334), .Y(n_940) );
INVx1_ASAP7_75t_L g943 ( .A(n_325), .Y(n_943) );
AND2x4_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
NAND3x1_ASAP7_75t_L g369 ( .A(n_326), .B(n_370), .C(n_371), .Y(n_369) );
NAND2x1p5_ASAP7_75t_L g821 ( .A(n_326), .B(n_371), .Y(n_821) );
OR2x4_ASAP7_75t_L g1430 ( .A(n_326), .B(n_379), .Y(n_1430) );
INVx1_ASAP7_75t_L g1433 ( .A(n_326), .Y(n_1433) );
AND2x4_ASAP7_75t_L g1437 ( .A(n_326), .B(n_354), .Y(n_1437) );
OR2x6_ASAP7_75t_L g1449 ( .A(n_326), .B(n_705), .Y(n_1449) );
INVx3_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx3_ASAP7_75t_L g341 ( .A(n_327), .Y(n_341) );
NAND2xp33_ASAP7_75t_SL g699 ( .A(n_327), .B(n_329), .Y(n_699) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND3x4_ASAP7_75t_L g340 ( .A(n_329), .B(n_341), .C(n_342), .Y(n_340) );
HB1xp67_ASAP7_75t_L g1452 ( .A(n_329), .Y(n_1452) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_331), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_331), .A2(n_495), .B1(n_575), .B2(n_576), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_331), .A2(n_495), .B1(n_630), .B2(n_631), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_331), .A2(n_495), .B1(n_1017), .B2(n_1018), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_331), .A2(n_495), .B1(n_1113), .B2(n_1114), .Y(n_1112) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g417 ( .A(n_337), .Y(n_417) );
AOI33xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_344), .A3(n_355), .B1(n_363), .B2(n_367), .B3(n_372), .Y(n_338) );
AOI33xp33_ASAP7_75t_L g502 ( .A1(n_339), .A2(n_503), .A3(n_506), .B1(n_511), .B2(n_512), .B3(n_515), .Y(n_502) );
AOI33xp33_ASAP7_75t_L g1023 ( .A1(n_339), .A2(n_515), .A3(n_1024), .B1(n_1027), .B2(n_1029), .B3(n_1031), .Y(n_1023) );
AOI33xp33_ASAP7_75t_L g1103 ( .A1(n_339), .A2(n_1104), .A3(n_1105), .B1(n_1109), .B2(n_1110), .B3(n_1111), .Y(n_1103) );
BUFx3_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI33xp33_ASAP7_75t_L g577 ( .A1(n_340), .A2(n_367), .A3(n_578), .B1(n_580), .B2(n_586), .B3(n_587), .Y(n_577) );
AOI33xp33_ASAP7_75t_L g634 ( .A1(n_340), .A2(n_515), .A3(n_635), .B1(n_638), .B2(n_642), .B3(n_643), .Y(n_634) );
AOI33xp33_ASAP7_75t_L g813 ( .A1(n_340), .A2(n_814), .A3(n_816), .B1(n_818), .B2(n_819), .B3(n_822), .Y(n_813) );
AOI33xp33_ASAP7_75t_L g855 ( .A1(n_340), .A2(n_819), .A3(n_856), .B1(n_857), .B2(n_858), .B3(n_859), .Y(n_855) );
AOI33xp33_ASAP7_75t_L g1060 ( .A1(n_340), .A2(n_1061), .A3(n_1063), .B1(n_1065), .B2(n_1067), .B3(n_1068), .Y(n_1060) );
AOI33xp33_ASAP7_75t_L g1488 ( .A1(n_340), .A2(n_819), .A3(n_1489), .B1(n_1490), .B2(n_1491), .B3(n_1492), .Y(n_1488) );
INVx3_ASAP7_75t_L g1440 ( .A(n_341), .Y(n_1440) );
INVx1_ASAP7_75t_L g488 ( .A(n_342), .Y(n_488) );
INVx2_ASAP7_75t_SL g559 ( .A(n_342), .Y(n_559) );
OAI31xp33_ASAP7_75t_SL g962 ( .A1(n_342), .A2(n_963), .A3(n_964), .B(n_968), .Y(n_962) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx2_ASAP7_75t_L g678 ( .A(n_343), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_343), .B(n_402), .Y(n_881) );
AND2x4_ASAP7_75t_L g563 ( .A(n_345), .B(n_389), .Y(n_563) );
AND2x4_ASAP7_75t_L g1021 ( .A(n_345), .B(n_389), .Y(n_1021) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx3_ASAP7_75t_L g504 ( .A(n_346), .Y(n_504) );
INVx8_ASAP7_75t_L g514 ( .A(n_346), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g974 ( .A(n_346), .Y(n_974) );
INVx8_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx3_ASAP7_75t_L g373 ( .A(n_347), .Y(n_373) );
BUFx3_ASAP7_75t_L g925 ( .A(n_347), .Y(n_925) );
AND2x2_ASAP7_75t_L g928 ( .A(n_347), .B(n_929), .Y(n_928) );
AND2x4_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
AND2x4_ASAP7_75t_L g359 ( .A(n_348), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVxp67_ASAP7_75t_L g360 ( .A(n_351), .Y(n_360) );
BUFx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx2_ASAP7_75t_L g374 ( .A(n_354), .Y(n_374) );
INVx2_ASAP7_75t_L g510 ( .A(n_354), .Y(n_510) );
BUFx3_ASAP7_75t_L g579 ( .A(n_354), .Y(n_579) );
BUFx2_ASAP7_75t_L g588 ( .A(n_354), .Y(n_588) );
BUFx2_ASAP7_75t_L g708 ( .A(n_354), .Y(n_708) );
AND2x2_ASAP7_75t_L g931 ( .A(n_354), .B(n_929), .Y(n_931) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI221xp5_ASAP7_75t_L g700 ( .A1(n_358), .A2(n_701), .B1(n_702), .B2(n_706), .C(n_707), .Y(n_700) );
INVx3_ASAP7_75t_L g817 ( .A(n_358), .Y(n_817) );
INVx1_ASAP7_75t_L g917 ( .A(n_358), .Y(n_917) );
OR2x6_ASAP7_75t_SL g945 ( .A(n_358), .B(n_946), .Y(n_945) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_359), .Y(n_366) );
BUFx8_ASAP7_75t_L g390 ( .A(n_359), .Y(n_390) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_359), .Y(n_583) );
BUFx3_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx12f_ASAP7_75t_L g505 ( .A(n_362), .Y(n_505) );
INVx5_ASAP7_75t_L g585 ( .A(n_362), .Y(n_585) );
BUFx2_ASAP7_75t_L g641 ( .A(n_362), .Y(n_641) );
AND2x4_ASAP7_75t_L g949 ( .A(n_362), .B(n_947), .Y(n_949) );
BUFx3_ASAP7_75t_L g1030 ( .A(n_362), .Y(n_1030) );
INVx8_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx3_ASAP7_75t_L g508 ( .A(n_365), .Y(n_508) );
INVx5_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_SL g640 ( .A(n_366), .Y(n_640) );
INVx3_ASAP7_75t_L g921 ( .A(n_366), .Y(n_921) );
BUFx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx2_ASAP7_75t_L g515 ( .A(n_368), .Y(n_515) );
INVx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx3_ASAP7_75t_L g710 ( .A(n_369), .Y(n_710) );
INVx2_ASAP7_75t_SL g637 ( .A(n_373), .Y(n_637) );
BUFx3_ASAP7_75t_L g815 ( .A(n_373), .Y(n_815) );
INVx1_ASAP7_75t_L g1026 ( .A(n_374), .Y(n_1026) );
OR2x6_ASAP7_75t_L g376 ( .A(n_377), .B(n_380), .Y(n_376) );
OR2x2_ASAP7_75t_L g590 ( .A(n_377), .B(n_380), .Y(n_590) );
INVx2_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx3_ASAP7_75t_L g1391 ( .A(n_379), .Y(n_1391) );
OR2x4_ASAP7_75t_L g1432 ( .A(n_379), .B(n_1433), .Y(n_1432) );
INVxp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g825 ( .A(n_381), .B(n_817), .Y(n_825) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g389 ( .A(n_382), .Y(n_389) );
OR2x2_ASAP7_75t_L g396 ( .A(n_382), .B(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g414 ( .A(n_382), .B(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_386), .Y(n_382) );
OR2x2_ASAP7_75t_L g698 ( .A(n_383), .B(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_SL g877 ( .A(n_383), .B(n_444), .Y(n_877) );
INVx1_ASAP7_75t_L g998 ( .A(n_383), .Y(n_998) );
HB1xp67_ASAP7_75t_L g1454 ( .A(n_383), .Y(n_1454) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx2_ASAP7_75t_L g413 ( .A(n_384), .Y(n_413) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g929 ( .A(n_386), .Y(n_929) );
INVx1_ASAP7_75t_L g947 ( .A(n_386), .Y(n_947) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_388), .A2(n_532), .B1(n_534), .B2(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_388), .A2(n_563), .B1(n_729), .B2(n_730), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_388), .A2(n_563), .B1(n_751), .B2(n_752), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_388), .A2(n_1020), .B1(n_1021), .B2(n_1022), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_388), .A2(n_563), .B1(n_1118), .B2(n_1120), .Y(n_1135) );
AND2x4_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx2_ASAP7_75t_SL g766 ( .A(n_390), .Y(n_766) );
HB1xp67_ASAP7_75t_L g1028 ( .A(n_390), .Y(n_1028) );
INVx2_ASAP7_75t_SL g1107 ( .A(n_390), .Y(n_1107) );
NOR3xp33_ASAP7_75t_L g695 ( .A(n_391), .B(n_696), .C(n_718), .Y(n_695) );
NOR3xp33_ASAP7_75t_L g851 ( .A(n_391), .B(n_852), .C(n_860), .Y(n_851) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx3_ASAP7_75t_L g516 ( .A(n_392), .Y(n_516) );
INVx3_ASAP7_75t_L g592 ( .A(n_392), .Y(n_592) );
NOR3xp33_ASAP7_75t_L g762 ( .A(n_392), .B(n_763), .C(n_775), .Y(n_762) );
NOR3xp33_ASAP7_75t_L g808 ( .A(n_392), .B(n_809), .C(n_823), .Y(n_808) );
AOI211xp5_ASAP7_75t_L g1485 ( .A1(n_392), .A2(n_1099), .B(n_1477), .C(n_1486), .Y(n_1485) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_406), .B(n_407), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_394), .B(n_565), .Y(n_564) );
AOI21xp33_ASAP7_75t_SL g593 ( .A1(n_394), .A2(n_594), .B(n_595), .Y(n_593) );
NAND2xp33_ASAP7_75t_L g644 ( .A(n_394), .B(n_645), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_394), .A2(n_692), .B(n_693), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g776 ( .A1(n_394), .A2(n_777), .B(n_778), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_394), .A2(n_806), .B(n_807), .Y(n_805) );
AOI21xp33_ASAP7_75t_L g848 ( .A1(n_394), .A2(n_849), .B(n_850), .Y(n_848) );
AOI21xp5_ASAP7_75t_L g1012 ( .A1(n_394), .A2(n_1013), .B(n_1014), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_394), .B(n_1094), .Y(n_1093) );
AOI221xp5_ASAP7_75t_L g1098 ( .A1(n_394), .A2(n_1099), .B1(n_1100), .B2(n_1101), .C(n_1102), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1464 ( .A(n_394), .B(n_1465), .Y(n_1464) );
INVx8_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_396), .B(n_400), .Y(n_395) );
BUFx3_ASAP7_75t_L g971 ( .A(n_397), .Y(n_971) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx6f_ASAP7_75t_L g715 ( .A(n_398), .Y(n_715) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx2_ASAP7_75t_L g705 ( .A(n_399), .Y(n_705) );
INVx1_ASAP7_75t_L g898 ( .A(n_401), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_402), .B(n_411), .Y(n_410) );
AND2x6_ASAP7_75t_L g450 ( .A(n_402), .B(n_434), .Y(n_450) );
INVx1_ASAP7_75t_L g481 ( .A(n_402), .Y(n_481) );
AND2x2_ASAP7_75t_L g787 ( .A(n_402), .B(n_788), .Y(n_787) );
INVx3_ASAP7_75t_L g447 ( .A(n_403), .Y(n_447) );
AND2x2_ASAP7_75t_L g455 ( .A(n_403), .B(n_428), .Y(n_455) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_403), .Y(n_528) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_408), .Y(n_561) );
INVx2_ASAP7_75t_L g650 ( .A(n_408), .Y(n_650) );
AND2x4_ASAP7_75t_L g408 ( .A(n_409), .B(n_414), .Y(n_408) );
AND2x4_ASAP7_75t_L g694 ( .A(n_409), .B(n_414), .Y(n_694) );
INVx2_ASAP7_75t_SL g1002 ( .A(n_409), .Y(n_1002) );
OR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_413), .Y(n_409) );
OR2x2_ASAP7_75t_L g884 ( .A(n_410), .B(n_413), .Y(n_884) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVxp67_ASAP7_75t_L g420 ( .A(n_413), .Y(n_420) );
INVx1_ASAP7_75t_L g913 ( .A(n_413), .Y(n_913) );
INVx1_ASAP7_75t_L g1427 ( .A(n_413), .Y(n_1427) );
INVx3_ASAP7_75t_L g982 ( .A(n_415), .Y(n_982) );
INVx4_ASAP7_75t_L g1393 ( .A(n_415), .Y(n_1393) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx2_ASAP7_75t_L g942 ( .A(n_416), .Y(n_942) );
BUFx2_ASAP7_75t_L g1444 ( .A(n_417), .Y(n_1444) );
INVx5_ASAP7_75t_L g501 ( .A(n_418), .Y(n_501) );
INVx3_ASAP7_75t_L g1099 ( .A(n_418), .Y(n_1099) );
OR2x6_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
OR2x2_ASAP7_75t_L g596 ( .A(n_419), .B(n_420), .Y(n_596) );
INVx2_ASAP7_75t_L g935 ( .A(n_419), .Y(n_935) );
OAI21xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_460), .B(n_485), .Y(n_421) );
INVx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_SL g519 ( .A(n_424), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_424), .B(n_1059), .Y(n_1080) );
AOI221xp5_ASAP7_75t_L g1121 ( .A1(n_424), .A2(n_450), .B1(n_1100), .B2(n_1122), .C(n_1124), .Y(n_1121) );
AND2x4_ASAP7_75t_L g424 ( .A(n_425), .B(n_428), .Y(n_424) );
INVx1_ASAP7_75t_L g530 ( .A(n_425), .Y(n_530) );
BUFx2_ASAP7_75t_L g602 ( .A(n_425), .Y(n_602) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx3_ASAP7_75t_L g449 ( .A(n_426), .Y(n_449) );
INVx2_ASAP7_75t_L g674 ( .A(n_426), .Y(n_674) );
BUFx3_ASAP7_75t_L g749 ( .A(n_426), .Y(n_749) );
AND2x4_ASAP7_75t_L g459 ( .A(n_428), .B(n_440), .Y(n_459) );
AND2x4_ASAP7_75t_SL g484 ( .A(n_428), .B(n_434), .Y(n_484) );
AND2x2_ASAP7_75t_L g953 ( .A(n_428), .B(n_440), .Y(n_953) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_428), .B(n_903), .Y(n_1476) );
HB1xp67_ASAP7_75t_L g1417 ( .A(n_429), .Y(n_1417) );
AOI21xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_445), .B(n_450), .Y(n_430) );
BUFx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx3_ASAP7_75t_L g522 ( .A(n_434), .Y(n_522) );
BUFx3_ASAP7_75t_L g604 ( .A(n_434), .Y(n_604) );
BUFx3_ASAP7_75t_L g623 ( .A(n_434), .Y(n_623) );
BUFx3_ASAP7_75t_L g745 ( .A(n_434), .Y(n_745) );
INVx1_ASAP7_75t_L g1037 ( .A(n_434), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_434), .B(n_1405), .Y(n_1404) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g469 ( .A(n_435), .Y(n_469) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g606 ( .A(n_439), .Y(n_606) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g747 ( .A(n_440), .Y(n_747) );
BUFx6f_ASAP7_75t_L g837 ( .A(n_440), .Y(n_837) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g472 ( .A(n_441), .Y(n_472) );
BUFx3_ASAP7_75t_L g657 ( .A(n_441), .Y(n_657) );
AND2x4_ASAP7_75t_L g1424 ( .A(n_441), .B(n_1417), .Y(n_1424) );
INVx4_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g524 ( .A(n_444), .Y(n_524) );
INVx4_ASAP7_75t_L g607 ( .A(n_444), .Y(n_607) );
AND2x4_ASAP7_75t_L g996 ( .A(n_444), .B(n_997), .Y(n_996) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g601 ( .A(n_447), .Y(n_601) );
INVx2_ASAP7_75t_SL g736 ( .A(n_447), .Y(n_736) );
INVx1_ASAP7_75t_L g795 ( .A(n_447), .Y(n_795) );
INVx1_ASAP7_75t_L g1076 ( .A(n_447), .Y(n_1076) );
BUFx3_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_450), .A2(n_521), .B(n_525), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_450), .A2(n_600), .B(n_603), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_450), .A2(n_656), .B(n_658), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_450), .A2(n_724), .B(n_725), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_450), .A2(n_744), .B(n_748), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g797 ( .A1(n_450), .A2(n_798), .B(n_800), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g841 ( .A1(n_450), .A2(n_842), .B(n_844), .Y(n_841) );
AOI21xp5_ASAP7_75t_SL g1034 ( .A1(n_450), .A2(n_1035), .B(n_1040), .Y(n_1034) );
INVx1_ASAP7_75t_L g1081 ( .A(n_450), .Y(n_1081) );
AOI221xp5_ASAP7_75t_L g1475 ( .A1(n_450), .A2(n_1476), .B1(n_1477), .B2(n_1478), .C(n_1479), .Y(n_1475) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B1(n_456), .B2(n_457), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_453), .A2(n_532), .B1(n_533), .B2(n_534), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_453), .A2(n_609), .B1(n_610), .B2(n_611), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_453), .A2(n_611), .B1(n_803), .B2(n_804), .Y(n_802) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx6f_ASAP7_75t_L g661 ( .A(n_455), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_455), .A2(n_459), .B1(n_751), .B2(n_752), .Y(n_750) );
AND2x4_ASAP7_75t_L g912 ( .A(n_455), .B(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_459), .Y(n_533) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_459), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_459), .A2(n_660), .B1(n_661), .B2(n_662), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_459), .A2(n_661), .B1(n_729), .B2(n_730), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_459), .A2(n_661), .B1(n_1020), .B2(n_1022), .Y(n_1041) );
AOI22xp5_ASAP7_75t_L g1077 ( .A1(n_459), .A2(n_661), .B1(n_1078), .B2(n_1079), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g1480 ( .A1(n_459), .A2(n_661), .B1(n_1481), .B2(n_1482), .Y(n_1480) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g555 ( .A(n_462), .Y(n_555) );
INVx2_ASAP7_75t_SL g618 ( .A(n_462), .Y(n_618) );
INVx2_ASAP7_75t_L g991 ( .A(n_462), .Y(n_991) );
INVx8_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx2_ASAP7_75t_L g889 ( .A(n_463), .Y(n_889) );
OR2x2_ASAP7_75t_L g1420 ( .A(n_463), .B(n_1409), .Y(n_1420) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_475), .Y(n_465) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g1473 ( .A(n_468), .Y(n_1473) );
BUFx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g1131 ( .A(n_469), .Y(n_1131) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g622 ( .A(n_471), .Y(n_622) );
INVx2_ASAP7_75t_L g1039 ( .A(n_471), .Y(n_1039) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g523 ( .A(n_472), .Y(n_523) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g548 ( .A(n_474), .Y(n_548) );
INVx1_ASAP7_75t_L g759 ( .A(n_474), .Y(n_759) );
INVx3_ASAP7_75t_L g838 ( .A(n_474), .Y(n_838) );
INVx1_ASAP7_75t_L g1089 ( .A(n_476), .Y(n_1089) );
INVx2_ASAP7_75t_L g558 ( .A(n_478), .Y(n_558) );
INVx2_ASAP7_75t_L g614 ( .A(n_478), .Y(n_614) );
NOR2x1_ASAP7_75t_L g478 ( .A(n_479), .B(n_481), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx2_ASAP7_75t_L g788 ( .A(n_480), .Y(n_788) );
INVx1_ASAP7_75t_L g883 ( .A(n_480), .Y(n_883) );
AND2x4_ASAP7_75t_L g1408 ( .A(n_480), .B(n_1409), .Y(n_1408) );
INVx2_ASAP7_75t_L g536 ( .A(n_482), .Y(n_536) );
INVx2_ASAP7_75t_L g613 ( .A(n_482), .Y(n_613) );
INVx4_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx3_ASAP7_75t_L g1126 ( .A(n_484), .Y(n_1126) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g914 ( .A1(n_487), .A2(n_915), .B(n_932), .C(n_950), .Y(n_914) );
BUFx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g761 ( .A(n_488), .Y(n_761) );
HB1xp67_ASAP7_75t_L g1048 ( .A(n_488), .Y(n_1048) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_567), .B1(n_568), .B2(n_683), .Y(n_489) );
INVx1_ASAP7_75t_L g683 ( .A(n_490), .Y(n_683) );
XOR2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_566), .Y(n_490) );
NAND3x1_ASAP7_75t_SL g491 ( .A(n_492), .B(n_517), .C(n_564), .Y(n_491) );
AND4x1_ASAP7_75t_L g492 ( .A(n_493), .B(n_499), .C(n_502), .D(n_516), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B1(n_497), .B2(n_498), .Y(n_493) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_501), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_501), .B(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g774 ( .A(n_510), .Y(n_774) );
INVx1_ASAP7_75t_L g1062 ( .A(n_510), .Y(n_1062) );
INVx2_ASAP7_75t_L g1493 ( .A(n_510), .Y(n_1493) );
BUFx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NAND4xp75_ASAP7_75t_L g1011 ( .A(n_516), .B(n_1012), .C(n_1015), .D(n_1032), .Y(n_1011) );
NAND3xp33_ASAP7_75t_SL g1102 ( .A(n_516), .B(n_1103), .C(n_1112), .Y(n_1102) );
O2A1O1Ixp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_535), .B(n_559), .C(n_560), .Y(n_517) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx3_ASAP7_75t_L g727 ( .A(n_528), .Y(n_727) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OAI221xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_541), .B1(n_542), .B2(n_546), .C(n_547), .Y(n_537) );
BUFx2_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_SL g757 ( .A(n_539), .Y(n_757) );
OR2x2_ASAP7_75t_L g906 ( .A(n_539), .B(n_902), .Y(n_906) );
BUFx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx6f_ASAP7_75t_L g668 ( .A(n_540), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g1373 ( .A1(n_542), .A2(n_1374), .B1(n_1375), .B2(n_1376), .Y(n_1373) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx4_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx3_ASAP7_75t_L g873 ( .A(n_545), .Y(n_873) );
INVx1_ASAP7_75t_L g1379 ( .A(n_545), .Y(n_1379) );
OAI221xp5_ASAP7_75t_L g1083 ( .A1(n_547), .A2(n_873), .B1(n_1084), .B2(n_1085), .C(n_1086), .Y(n_1083) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_551), .B1(n_553), .B2(n_556), .Y(n_549) );
OAI221xp5_ASAP7_75t_L g615 ( .A1(n_551), .A2(n_616), .B1(n_617), .B2(n_619), .C(n_620), .Y(n_615) );
INVx1_ASAP7_75t_L g870 ( .A(n_551), .Y(n_870) );
OAI221xp5_ASAP7_75t_L g1043 ( .A1(n_551), .A2(n_554), .B1(n_1044), .B2(n_1045), .C(n_1046), .Y(n_1043) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g988 ( .A1(n_552), .A2(n_989), .B1(n_990), .B2(n_991), .Y(n_988) );
OAI22x1_ASAP7_75t_SL g994 ( .A1(n_552), .A2(n_972), .B1(n_991), .B2(n_995), .Y(n_994) );
BUFx3_ASAP7_75t_L g1383 ( .A(n_552), .Y(n_1383) );
BUFx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g869 ( .A(n_554), .Y(n_869) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OAI21xp5_ASAP7_75t_L g597 ( .A1(n_559), .A2(n_598), .B(n_612), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g1484 ( .A1(n_563), .A2(n_825), .B1(n_1481), .B2(n_1482), .Y(n_1484) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B1(n_624), .B2(n_682), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND3xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_593), .C(n_597), .Y(n_571) );
NOR3xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_589), .C(n_591), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_577), .Y(n_573) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g712 ( .A(n_583), .Y(n_712) );
AND2x4_ASAP7_75t_L g1447 ( .A(n_583), .B(n_1433), .Y(n_1447) );
INVx2_ASAP7_75t_R g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g1066 ( .A(n_585), .Y(n_1066) );
INVx1_ASAP7_75t_L g1108 ( .A(n_585), .Y(n_1108) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND4xp25_ASAP7_75t_SL g628 ( .A(n_592), .B(n_629), .C(n_632), .D(n_634), .Y(n_628) );
AND4x1_ASAP7_75t_L g1054 ( .A(n_592), .B(n_1055), .C(n_1058), .D(n_1060), .Y(n_1054) );
BUFx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_611), .A2(n_661), .B1(n_846), .B2(n_847), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_611), .A2(n_1118), .B1(n_1119), .B2(n_1120), .Y(n_1117) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI22xp33_ASAP7_75t_L g1367 ( .A1(n_618), .A2(n_1368), .B1(n_1369), .B2(n_1372), .Y(n_1367) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g682 ( .A(n_624), .Y(n_682) );
NAND2x1p5_ASAP7_75t_L g624 ( .A(n_625), .B(n_646), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_644), .Y(n_626) );
INVxp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NOR2xp33_ASAP7_75t_SL g679 ( .A(n_628), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_644), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_653), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .B(n_652), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_663), .B(n_675), .Y(n_653) );
INVx1_ASAP7_75t_L g671 ( .A(n_657), .Y(n_671) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_657), .Y(n_799) );
BUFx2_ASAP7_75t_L g1123 ( .A(n_657), .Y(n_1123) );
HB1xp67_ASAP7_75t_L g1119 ( .A(n_661), .Y(n_1119) );
OAI211xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B(n_669), .C(n_672), .Y(n_664) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g733 ( .A(n_667), .Y(n_733) );
INVx2_ASAP7_75t_L g1084 ( .A(n_667), .Y(n_1084) );
INVx4_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
BUFx4f_ASAP7_75t_L g792 ( .A(n_668), .Y(n_792) );
BUFx4f_ASAP7_75t_L g875 ( .A(n_668), .Y(n_875) );
OR2x6_ASAP7_75t_L g885 ( .A(n_668), .B(n_886), .Y(n_885) );
BUFx4f_ASAP7_75t_L g1073 ( .A(n_668), .Y(n_1073) );
BUFx4f_ASAP7_75t_L g1376 ( .A(n_668), .Y(n_1376) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g843 ( .A(n_671), .Y(n_843) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx3_ASAP7_75t_L g903 ( .A(n_674), .Y(n_903) );
OAI21xp5_ASAP7_75t_L g721 ( .A1(n_675), .A2(n_722), .B(n_731), .Y(n_721) );
OAI21xp5_ASAP7_75t_SL g784 ( .A1(n_675), .A2(n_785), .B(n_796), .Y(n_784) );
OAI21xp5_ASAP7_75t_SL g830 ( .A1(n_675), .A2(n_831), .B(n_840), .Y(n_830) );
AOI21xp5_ASAP7_75t_L g1115 ( .A1(n_675), .A2(n_1116), .B(n_1134), .Y(n_1115) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g1467 ( .A(n_676), .Y(n_1467) );
BUFx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OR2x6_ASAP7_75t_L g820 ( .A(n_678), .B(n_821), .Y(n_820) );
AND2x4_ASAP7_75t_L g893 ( .A(n_678), .B(n_894), .Y(n_893) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_862), .B1(n_1006), .B2(n_1007), .Y(n_684) );
INVx2_ASAP7_75t_L g1007 ( .A(n_685), .Y(n_1007) );
AOI22x1_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .B1(n_781), .B2(n_861), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
BUFx3_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AO22x2_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_738), .B1(n_739), .B2(n_780), .Y(n_688) );
INVx1_ASAP7_75t_L g780 ( .A(n_689), .Y(n_780) );
AND4x1_ASAP7_75t_L g690 ( .A(n_691), .B(n_695), .C(n_721), .D(n_737), .Y(n_690) );
OAI22xp5_ASAP7_75t_SL g696 ( .A1(n_697), .A2(n_700), .B1(n_709), .B2(n_711), .Y(n_696) );
BUFx4f_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
BUFx8_ASAP7_75t_L g764 ( .A(n_698), .Y(n_764) );
BUFx2_ASAP7_75t_L g922 ( .A(n_699), .Y(n_922) );
OAI221xp5_ASAP7_75t_L g765 ( .A1(n_702), .A2(n_766), .B1(n_767), .B2(n_768), .C(n_769), .Y(n_765) );
INVx3_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
BUFx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
BUFx3_ASAP7_75t_L g1396 ( .A(n_705), .Y(n_1396) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
CKINVDCx5p33_ASAP7_75t_R g770 ( .A(n_710), .Y(n_770) );
INVx2_ASAP7_75t_L g1398 ( .A(n_710), .Y(n_1398) );
OAI221xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_713), .B1(n_714), .B2(n_716), .C(n_717), .Y(n_711) );
INVx1_ASAP7_75t_L g1064 ( .A(n_712), .Y(n_1064) );
OAI22xp33_ASAP7_75t_SL g1397 ( .A1(n_712), .A2(n_714), .B1(n_1375), .B2(n_1385), .Y(n_1397) );
OAI211xp5_ASAP7_75t_L g732 ( .A1(n_713), .A2(n_733), .B(n_734), .C(n_735), .Y(n_732) );
OAI221xp5_ASAP7_75t_L g771 ( .A1(n_714), .A2(n_755), .B1(n_766), .B2(n_772), .C(n_773), .Y(n_771) );
CKINVDCx8_ASAP7_75t_R g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_720), .A2(n_789), .B1(n_811), .B2(n_812), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_720), .A2(n_811), .B1(n_833), .B2(n_854), .Y(n_853) );
AOI22xp5_ASAP7_75t_L g1055 ( .A1(n_720), .A2(n_811), .B1(n_1056), .B2(n_1057), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1487 ( .A1(n_720), .A2(n_811), .B1(n_1470), .B2(n_1471), .Y(n_1487) );
INVx2_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g801 ( .A(n_727), .Y(n_801) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AND4x1_ASAP7_75t_L g740 ( .A(n_741), .B(n_762), .C(n_776), .D(n_779), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_753), .B(n_761), .Y(n_741) );
INVx2_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
OAI211xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_756), .B(n_758), .C(n_760), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g1377 ( .A1(n_756), .A2(n_1378), .B1(n_1380), .B2(n_1381), .Y(n_1377) );
INVx5_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
O2A1O1Ixp5_ASAP7_75t_SL g1069 ( .A1(n_761), .A2(n_1070), .B(n_1082), .C(n_1091), .Y(n_1069) );
OAI22xp5_ASAP7_75t_SL g763 ( .A1(n_764), .A2(n_765), .B1(n_770), .B2(n_771), .Y(n_763) );
OAI33xp33_ASAP7_75t_L g1387 ( .A1(n_764), .A2(n_1388), .A3(n_1394), .B1(n_1397), .B2(n_1398), .B3(n_1399), .Y(n_1387) );
INVx1_ASAP7_75t_L g1110 ( .A(n_770), .Y(n_1110) );
INVx1_ASAP7_75t_L g861 ( .A(n_781), .Y(n_861) );
XNOR2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_828), .Y(n_781) );
INVx1_ASAP7_75t_L g827 ( .A(n_783), .Y(n_827) );
NAND3xp33_ASAP7_75t_L g783 ( .A(n_784), .B(n_805), .C(n_808), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_787), .B(n_789), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_787), .B(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g1133 ( .A(n_787), .Y(n_1133) );
AOI222xp33_ASAP7_75t_L g1469 ( .A1(n_787), .A2(n_1126), .B1(n_1470), .B2(n_1471), .C1(n_1472), .C2(n_1474), .Y(n_1469) );
OAI211xp5_ASAP7_75t_L g790 ( .A1(n_791), .A2(n_792), .B(n_793), .C(n_794), .Y(n_790) );
OAI211xp5_ASAP7_75t_L g834 ( .A1(n_792), .A2(n_835), .B(n_836), .C(n_839), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_813), .Y(n_809) );
INVx2_ASAP7_75t_L g1395 ( .A(n_817), .Y(n_1395) );
INVx1_ASAP7_75t_SL g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g1068 ( .A(n_820), .Y(n_1068) );
INVx3_ASAP7_75t_L g976 ( .A(n_821), .Y(n_976) );
INVx2_ASAP7_75t_SL g824 ( .A(n_825), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_825), .A2(n_1021), .B1(n_1078), .B2(n_1079), .Y(n_1092) );
OAI22xp5_ASAP7_75t_SL g1224 ( .A1(n_826), .A2(n_1225), .B1(n_1226), .B2(n_1227), .Y(n_1224) );
NAND3xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_848), .C(n_851), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_853), .B(n_855), .Y(n_852) );
INVx1_ASAP7_75t_L g1006 ( .A(n_862), .Y(n_1006) );
INVxp67_ASAP7_75t_SL g862 ( .A(n_863), .Y(n_862) );
XNOR2x1_ASAP7_75t_L g863 ( .A(n_864), .B(n_955), .Y(n_863) );
XNOR2x1_ASAP7_75t_L g864 ( .A(n_865), .B(n_954), .Y(n_864) );
OR2x2_ASAP7_75t_L g865 ( .A(n_866), .B(n_914), .Y(n_865) );
NAND3xp33_ASAP7_75t_SL g866 ( .A(n_867), .B(n_895), .C(n_908), .Y(n_866) );
AOI211xp5_ASAP7_75t_SL g867 ( .A1(n_868), .A2(n_871), .B(n_878), .C(n_887), .Y(n_867) );
INVx2_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
OAI221xp5_ASAP7_75t_L g890 ( .A1(n_873), .A2(n_875), .B1(n_891), .B2(n_892), .C(n_893), .Y(n_890) );
INVxp67_ASAP7_75t_SL g874 ( .A(n_875), .Y(n_874) );
INVx2_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g1001 ( .A(n_879), .Y(n_1001) );
NAND2x2_ASAP7_75t_L g879 ( .A(n_880), .B(n_882), .Y(n_879) );
INVx1_ASAP7_75t_L g886 ( .A(n_880), .Y(n_886) );
INVx2_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx2_ASAP7_75t_SL g882 ( .A(n_883), .Y(n_882) );
CKINVDCx5p33_ASAP7_75t_R g1005 ( .A(n_885), .Y(n_1005) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
HB1xp67_ASAP7_75t_L g992 ( .A(n_893), .Y(n_992) );
INVx4_ASAP7_75t_L g1366 ( .A(n_893), .Y(n_1366) );
AOI222xp33_ASAP7_75t_L g895 ( .A1(n_896), .A2(n_899), .B1(n_900), .B2(n_904), .C1(n_905), .C2(n_907), .Y(n_895) );
AOI21xp33_ASAP7_75t_SL g1003 ( .A1(n_896), .A2(n_1004), .B(n_1005), .Y(n_1003) );
AND2x4_ASAP7_75t_L g896 ( .A(n_897), .B(n_898), .Y(n_896) );
AOI222xp33_ASAP7_75t_L g999 ( .A1(n_900), .A2(n_966), .B1(n_978), .B2(n_1000), .C1(n_1001), .C2(n_1002), .Y(n_999) );
AND2x4_ASAP7_75t_L g900 ( .A(n_901), .B(n_903), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
AOI211xp5_ASAP7_75t_L g932 ( .A1(n_904), .A2(n_933), .B(n_936), .C(n_944), .Y(n_932) );
AOI222xp33_ASAP7_75t_L g986 ( .A1(n_905), .A2(n_967), .B1(n_987), .B2(n_992), .C1(n_993), .C2(n_996), .Y(n_986) );
INVx2_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_909), .B(n_910), .Y(n_908) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx3_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
HB1xp67_ASAP7_75t_L g957 ( .A(n_912), .Y(n_957) );
AND2x4_ASAP7_75t_L g952 ( .A(n_913), .B(n_953), .Y(n_952) );
AOI221xp5_ASAP7_75t_L g915 ( .A1(n_916), .A2(n_918), .B1(n_919), .B2(n_923), .C(n_926), .Y(n_915) );
INVx2_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
OAI221xp5_ASAP7_75t_L g969 ( .A1(n_921), .A2(n_970), .B1(n_971), .B2(n_972), .C(n_973), .Y(n_969) );
BUFx2_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
AOI22xp5_ASAP7_75t_L g977 ( .A1(n_928), .A2(n_931), .B1(n_958), .B2(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
INVx2_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx4_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_938), .A2(n_940), .B1(n_966), .B2(n_967), .Y(n_965) );
INVx2_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
OR2x6_ASAP7_75t_L g941 ( .A(n_942), .B(n_943), .Y(n_941) );
INVx2_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx3_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_951), .B(n_952), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_952), .B(n_961), .Y(n_960) );
AOI211x1_ASAP7_75t_L g956 ( .A1(n_957), .A2(n_958), .B(n_959), .C(n_985), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_960), .B(n_962), .Y(n_959) );
NAND3xp33_ASAP7_75t_L g968 ( .A(n_969), .B(n_977), .C(n_979), .Y(n_968) );
INVx3_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
OAI211xp5_ASAP7_75t_L g979 ( .A1(n_980), .A2(n_981), .B(n_983), .C(n_984), .Y(n_979) );
INVx3_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVx2_ASAP7_75t_L g1400 ( .A(n_982), .Y(n_1400) );
NAND3xp33_ASAP7_75t_L g985 ( .A(n_986), .B(n_999), .C(n_1003), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_991), .A2(n_1088), .B1(n_1089), .B2(n_1090), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1382 ( .A1(n_991), .A2(n_1383), .B1(n_1384), .B2(n_1385), .Y(n_1382) );
CKINVDCx5p33_ASAP7_75t_R g1386 ( .A(n_996), .Y(n_1386) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1008), .Y(n_1142) );
AOI22xp5_ASAP7_75t_L g1008 ( .A1(n_1009), .A2(n_1010), .B1(n_1049), .B2(n_1140), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
AND3x1_ASAP7_75t_L g1015 ( .A(n_1016), .B(n_1019), .C(n_1023), .Y(n_1015) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
OAI21xp5_ASAP7_75t_L g1032 ( .A1(n_1033), .A2(n_1042), .B(n_1048), .Y(n_1032) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx1_ASAP7_75t_L g1047 ( .A(n_1037), .Y(n_1047) );
INVx2_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1049), .Y(n_1140) );
AOI22xp5_ASAP7_75t_L g1049 ( .A1(n_1050), .A2(n_1051), .B1(n_1096), .B2(n_1137), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
HB1xp67_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
XOR2xp5_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1095), .Y(n_1052) );
NAND3xp33_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1069), .C(n_1093), .Y(n_1053) );
NAND4xp25_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1077), .C(n_1080), .D(n_1081), .Y(n_1070) );
OAI211xp5_ASAP7_75t_L g1071 ( .A1(n_1072), .A2(n_1073), .B(n_1074), .C(n_1075), .Y(n_1071) );
XNOR2xp5_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1136), .Y(n_1096) );
OAI22xp5_ASAP7_75t_L g1137 ( .A1(n_1097), .A2(n_1136), .B1(n_1138), .B2(n_1139), .Y(n_1137) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1097), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1115), .Y(n_1097) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
AOI222xp33_ASAP7_75t_L g1125 ( .A1(n_1113), .A2(n_1114), .B1(n_1126), .B2(n_1127), .C1(n_1128), .C2(n_1132), .Y(n_1125) );
NAND3xp33_ASAP7_75t_L g1116 ( .A(n_1117), .B(n_1121), .C(n_1125), .Y(n_1116) );
INVx2_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
CKINVDCx5p33_ASAP7_75t_R g1138 ( .A(n_1136), .Y(n_1138) );
OAI221xp5_ASAP7_75t_L g1143 ( .A1(n_1144), .A2(n_1356), .B1(n_1359), .B2(n_1455), .C(n_1458), .Y(n_1143) );
NOR3xp33_ASAP7_75t_L g1144 ( .A(n_1145), .B(n_1293), .C(n_1332), .Y(n_1144) );
NAND3xp33_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1228), .C(n_1260), .Y(n_1145) );
AOI211xp5_ASAP7_75t_L g1146 ( .A1(n_1147), .A2(n_1172), .B(n_1189), .C(n_1208), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1147), .B(n_1207), .Y(n_1206) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1147), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1163), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1148), .B(n_1169), .Y(n_1276) );
NAND3xp33_ASAP7_75t_L g1280 ( .A(n_1148), .B(n_1266), .C(n_1281), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1148), .B(n_1198), .Y(n_1286) );
OR2x2_ASAP7_75t_L g1304 ( .A(n_1148), .B(n_1169), .Y(n_1304) );
NAND2xp5_ASAP7_75t_L g1318 ( .A(n_1148), .B(n_1261), .Y(n_1318) );
CKINVDCx6p67_ASAP7_75t_R g1148 ( .A(n_1149), .Y(n_1148) );
OR2x2_ASAP7_75t_L g1196 ( .A(n_1149), .B(n_1169), .Y(n_1196) );
OR2x2_ASAP7_75t_L g1267 ( .A(n_1149), .B(n_1268), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1296 ( .A(n_1149), .B(n_1198), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1149), .B(n_1169), .Y(n_1297) );
CKINVDCx5p33_ASAP7_75t_R g1320 ( .A(n_1149), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1149), .B(n_1223), .Y(n_1325) );
OR2x6_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1157), .Y(n_1149) );
OR2x2_ASAP7_75t_L g1309 ( .A(n_1150), .B(n_1157), .Y(n_1309) );
INVx2_ASAP7_75t_L g1225 ( .A(n_1151), .Y(n_1225) );
AND2x6_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1153), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1152), .B(n_1156), .Y(n_1155) );
AND2x4_ASAP7_75t_L g1158 ( .A(n_1152), .B(n_1159), .Y(n_1158) );
AND2x6_ASAP7_75t_L g1161 ( .A(n_1152), .B(n_1162), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1152), .B(n_1156), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1152), .B(n_1156), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1358 ( .A(n_1152), .B(n_1159), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1154), .B(n_1160), .Y(n_1159) );
HB1xp67_ASAP7_75t_L g1502 ( .A(n_1159), .Y(n_1502) );
AOI21xp33_ASAP7_75t_L g1245 ( .A1(n_1163), .A2(n_1222), .B(n_1246), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1163), .B(n_1193), .Y(n_1344) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1168), .Y(n_1163) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1164), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1164), .B(n_1169), .Y(n_1210) );
OR2x2_ASAP7_75t_L g1259 ( .A(n_1164), .B(n_1169), .Y(n_1259) );
OR2x2_ASAP7_75t_L g1282 ( .A(n_1164), .B(n_1179), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1165), .B(n_1167), .Y(n_1164) );
INVxp67_ASAP7_75t_L g1227 ( .A(n_1166), .Y(n_1227) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
OAI221xp5_ASAP7_75t_L g1189 ( .A1(n_1169), .A2(n_1190), .B1(n_1194), .B2(n_1200), .C(n_1206), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1169), .B(n_1199), .Y(n_1221) );
A2O1A1Ixp33_ASAP7_75t_L g1228 ( .A1(n_1169), .A2(n_1229), .B(n_1243), .C(n_1244), .Y(n_1228) );
INVx3_ASAP7_75t_L g1289 ( .A(n_1169), .Y(n_1289) );
O2A1O1Ixp33_ASAP7_75t_L g1333 ( .A1(n_1169), .A2(n_1334), .B(n_1335), .C(n_1336), .Y(n_1333) );
NAND2xp5_ASAP7_75t_L g1347 ( .A(n_1169), .B(n_1179), .Y(n_1347) );
AND2x4_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1171), .Y(n_1169) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
AOI21xp5_ASAP7_75t_L g1336 ( .A1(n_1173), .A2(n_1259), .B(n_1337), .Y(n_1336) );
OR2x2_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1178), .Y(n_1173) );
INVx2_ASAP7_75t_L g1191 ( .A(n_1174), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1174), .B(n_1203), .Y(n_1207) );
BUFx2_ASAP7_75t_L g1234 ( .A(n_1174), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1174), .B(n_1182), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1174), .B(n_1248), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1175), .B(n_1176), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1182), .Y(n_1178) );
INVx2_ASAP7_75t_L g1193 ( .A(n_1179), .Y(n_1193) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1179), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1241 ( .A(n_1179), .B(n_1234), .Y(n_1241) );
OR2x2_ASAP7_75t_L g1251 ( .A(n_1179), .B(n_1252), .Y(n_1251) );
NOR2xp33_ASAP7_75t_L g1301 ( .A(n_1179), .B(n_1302), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1179), .B(n_1203), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1181), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_1182), .B(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1182), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g1322 ( .A(n_1182), .B(n_1323), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1182), .B(n_1241), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1186), .Y(n_1182) );
INVx2_ASAP7_75t_L g1204 ( .A(n_1183), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1183), .B(n_1205), .Y(n_1248) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1183), .B(n_1234), .Y(n_1252) );
OR2x2_ASAP7_75t_L g1183 ( .A(n_1184), .B(n_1185), .Y(n_1183) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1186), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1186), .B(n_1191), .Y(n_1214) );
OR2x2_ASAP7_75t_L g1233 ( .A(n_1186), .B(n_1234), .Y(n_1233) );
AND3x1_ASAP7_75t_L g1237 ( .A(n_1186), .B(n_1191), .C(n_1204), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1186), .B(n_1234), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1186), .B(n_1204), .Y(n_1266) );
OAI21xp33_ASAP7_75t_L g1298 ( .A1(n_1186), .A2(n_1299), .B(n_1300), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1188), .Y(n_1186) );
OR2x2_ASAP7_75t_L g1190 ( .A(n_1191), .B(n_1192), .Y(n_1190) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1191), .B(n_1201), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1191), .B(n_1203), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1191), .B(n_1248), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_1191), .B(n_1204), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1323 ( .A(n_1191), .B(n_1193), .Y(n_1323) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1193), .Y(n_1213) );
NAND2xp5_ASAP7_75t_L g1247 ( .A(n_1193), .B(n_1248), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1193), .B(n_1255), .Y(n_1254) );
NOR2xp33_ASAP7_75t_L g1274 ( .A(n_1193), .B(n_1252), .Y(n_1274) );
O2A1O1Ixp33_ASAP7_75t_L g1283 ( .A1(n_1193), .A2(n_1217), .B(n_1284), .C(n_1285), .Y(n_1283) );
NOR2xp33_ASAP7_75t_L g1292 ( .A(n_1193), .B(n_1233), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1307 ( .A(n_1193), .B(n_1198), .Y(n_1307) );
NOR2xp33_ASAP7_75t_L g1194 ( .A(n_1195), .B(n_1197), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
OAI21xp33_ASAP7_75t_L g1277 ( .A1(n_1196), .A2(n_1278), .B(n_1280), .Y(n_1277) );
OAI222xp33_ASAP7_75t_L g1326 ( .A1(n_1196), .A2(n_1285), .B1(n_1327), .B2(n_1328), .C1(n_1329), .C2(n_1331), .Y(n_1326) );
OAI211xp5_ASAP7_75t_L g1229 ( .A1(n_1197), .A2(n_1230), .B(n_1235), .C(n_1238), .Y(n_1229) );
INVx2_ASAP7_75t_L g1291 ( .A(n_1197), .Y(n_1291) );
O2A1O1Ixp33_ASAP7_75t_L g1312 ( .A1(n_1197), .A2(n_1253), .B(n_1279), .C(n_1313), .Y(n_1312) );
NAND2xp5_ASAP7_75t_L g1354 ( .A(n_1197), .B(n_1355), .Y(n_1354) );
INVx2_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
OR2x2_ASAP7_75t_L g1238 ( .A(n_1198), .B(n_1239), .Y(n_1238) );
INVx2_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
OAI211xp5_ASAP7_75t_SL g1303 ( .A1(n_1200), .A2(n_1261), .B(n_1304), .C(n_1305), .Y(n_1303) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1201), .Y(n_1316) );
NAND2xp5_ASAP7_75t_L g1201 ( .A(n_1202), .B(n_1203), .Y(n_1201) );
INVx2_ASAP7_75t_L g1232 ( .A(n_1202), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1202), .B(n_1258), .Y(n_1257) );
NAND2xp5_ASAP7_75t_SL g1299 ( .A(n_1202), .B(n_1210), .Y(n_1299) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1203), .Y(n_1242) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1203), .B(n_1257), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_1203), .B(n_1323), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1205), .Y(n_1203) );
OR2x2_ASAP7_75t_L g1302 ( .A(n_1204), .B(n_1234), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1204), .B(n_1234), .Y(n_1330) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1207), .Y(n_1331) );
O2A1O1Ixp33_ASAP7_75t_SL g1208 ( .A1(n_1209), .A2(n_1211), .B(n_1215), .C(n_1222), .Y(n_1208) );
INVx2_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
OAI21xp5_ASAP7_75t_SL g1314 ( .A1(n_1210), .A2(n_1315), .B(n_1316), .Y(n_1314) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
NOR2xp33_ASAP7_75t_L g1212 ( .A(n_1213), .B(n_1214), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_1213), .B(n_1221), .Y(n_1220) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
AOI21xp33_ASAP7_75t_L g1216 ( .A1(n_1217), .A2(n_1219), .B(n_1220), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
AOI221xp5_ASAP7_75t_L g1305 ( .A1(n_1219), .A2(n_1241), .B1(n_1266), .B2(n_1306), .C(n_1308), .Y(n_1305) );
AOI21xp33_ASAP7_75t_L g1313 ( .A1(n_1219), .A2(n_1220), .B(n_1284), .Y(n_1313) );
OAI21xp5_ASAP7_75t_L g1249 ( .A1(n_1221), .A2(n_1250), .B(n_1253), .Y(n_1249) );
CKINVDCx6p67_ASAP7_75t_R g1268 ( .A(n_1221), .Y(n_1268) );
INVx3_ASAP7_75t_L g1243 ( .A(n_1222), .Y(n_1243) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1222), .B(n_1289), .Y(n_1288) );
INVx2_ASAP7_75t_SL g1222 ( .A(n_1223), .Y(n_1222) );
INVx2_ASAP7_75t_SL g1261 ( .A(n_1223), .Y(n_1261) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
NOR2xp33_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1233), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1232), .B(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1232), .Y(n_1272) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
A2O1A1Ixp33_ASAP7_75t_L g1345 ( .A1(n_1236), .A2(n_1289), .B(n_1324), .C(n_1346), .Y(n_1345) );
AND2x2_ASAP7_75t_SL g1353 ( .A(n_1237), .B(n_1258), .Y(n_1353) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1238), .Y(n_1334) );
OR2x2_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1242), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1241), .B(n_1248), .Y(n_1315) );
O2A1O1Ixp33_ASAP7_75t_L g1321 ( .A1(n_1243), .A2(n_1258), .B(n_1322), .C(n_1324), .Y(n_1321) );
NAND3xp33_ASAP7_75t_L g1244 ( .A(n_1245), .B(n_1249), .C(n_1256), .Y(n_1244) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
OAI211xp5_ASAP7_75t_L g1311 ( .A1(n_1251), .A2(n_1268), .B(n_1312), .C(n_1314), .Y(n_1311) );
AOI211xp5_ASAP7_75t_L g1275 ( .A1(n_1253), .A2(n_1276), .B(n_1277), .C(n_1283), .Y(n_1275) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1255), .Y(n_1351) );
OAI21xp5_ASAP7_75t_L g1269 ( .A1(n_1258), .A2(n_1270), .B(n_1274), .Y(n_1269) );
INVx2_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
AOI22xp5_ASAP7_75t_L g1260 ( .A1(n_1261), .A2(n_1262), .B1(n_1287), .B2(n_1290), .Y(n_1260) );
NAND3xp33_ASAP7_75t_L g1262 ( .A(n_1263), .B(n_1269), .C(n_1275), .Y(n_1262) );
INVxp67_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
NOR2xp33_ASAP7_75t_L g1264 ( .A(n_1265), .B(n_1267), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
AOI211xp5_ASAP7_75t_L g1339 ( .A1(n_1270), .A2(n_1289), .B(n_1340), .C(n_1342), .Y(n_1339) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1272), .B(n_1273), .Y(n_1271) );
NAND2xp5_ASAP7_75t_L g1341 ( .A(n_1273), .B(n_1306), .Y(n_1341) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1273), .Y(n_1350) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
INVxp33_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1291), .B(n_1292), .Y(n_1290) );
AOI21xp5_ASAP7_75t_L g1352 ( .A1(n_1291), .A2(n_1335), .B(n_1353), .Y(n_1352) );
AOI221xp5_ASAP7_75t_SL g1293 ( .A1(n_1294), .A2(n_1309), .B1(n_1310), .B2(n_1317), .C(n_1319), .Y(n_1293) );
O2A1O1Ixp33_ASAP7_75t_L g1294 ( .A1(n_1295), .A2(n_1297), .B(n_1298), .C(n_1303), .Y(n_1294) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
INVxp67_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
AOI211xp5_ASAP7_75t_L g1319 ( .A1(n_1311), .A2(n_1320), .B(n_1321), .C(n_1326), .Y(n_1319) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1315), .Y(n_1327) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
A2O1A1Ixp33_ASAP7_75t_L g1332 ( .A1(n_1320), .A2(n_1333), .B(n_1339), .C(n_1345), .Y(n_1332) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
CKINVDCx14_ASAP7_75t_R g1329 ( .A(n_1330), .Y(n_1329) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_1330), .B(n_1344), .Y(n_1343) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
INVxp67_ASAP7_75t_SL g1342 ( .A(n_1343), .Y(n_1342) );
OAI211xp5_ASAP7_75t_SL g1346 ( .A1(n_1347), .A2(n_1348), .B(n_1352), .C(n_1354), .Y(n_1346) );
INVxp67_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
NAND2xp5_ASAP7_75t_SL g1349 ( .A(n_1350), .B(n_1351), .Y(n_1349) );
CKINVDCx20_ASAP7_75t_R g1356 ( .A(n_1357), .Y(n_1356) );
CKINVDCx5p33_ASAP7_75t_R g1357 ( .A(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
INVx2_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
NAND3xp33_ASAP7_75t_L g1363 ( .A(n_1364), .B(n_1401), .C(n_1428), .Y(n_1363) );
NOR2xp33_ASAP7_75t_L g1364 ( .A(n_1365), .B(n_1387), .Y(n_1364) );
OAI33xp33_ASAP7_75t_L g1365 ( .A1(n_1366), .A2(n_1367), .A3(n_1373), .B1(n_1377), .B2(n_1382), .B3(n_1386), .Y(n_1365) );
OAI22xp33_ASAP7_75t_L g1388 ( .A1(n_1368), .A2(n_1380), .B1(n_1389), .B2(n_1392), .Y(n_1388) );
INVx3_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
BUFx6f_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
OAI22xp33_ASAP7_75t_L g1399 ( .A1(n_1372), .A2(n_1381), .B1(n_1389), .B2(n_1400), .Y(n_1399) );
OAI22xp5_ASAP7_75t_L g1394 ( .A1(n_1374), .A2(n_1384), .B1(n_1395), .B2(n_1396), .Y(n_1394) );
INVx2_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
INVx2_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1393), .Y(n_1435) );
OAI31xp33_ASAP7_75t_L g1401 ( .A1(n_1402), .A2(n_1414), .A3(n_1421), .B(n_1425), .Y(n_1401) );
INVx3_ASAP7_75t_L g1403 ( .A(n_1404), .Y(n_1403) );
AOI22xp33_ASAP7_75t_L g1406 ( .A1(n_1407), .A2(n_1408), .B1(n_1410), .B2(n_1411), .Y(n_1406) );
AOI22xp33_ASAP7_75t_L g1438 ( .A1(n_1407), .A2(n_1439), .B1(n_1442), .B2(n_1443), .Y(n_1438) );
INVx2_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
INVx2_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
BUFx6f_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
INVxp67_ASAP7_75t_SL g1418 ( .A(n_1419), .Y(n_1418) );
INVx2_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
CKINVDCx16_ASAP7_75t_R g1423 ( .A(n_1424), .Y(n_1423) );
BUFx2_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
OAI31xp33_ASAP7_75t_L g1428 ( .A1(n_1429), .A2(n_1434), .A3(n_1445), .B(n_1450), .Y(n_1428) );
BUFx3_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
CKINVDCx8_ASAP7_75t_R g1436 ( .A(n_1437), .Y(n_1436) );
AND2x4_ASAP7_75t_L g1439 ( .A(n_1440), .B(n_1441), .Y(n_1439) );
AND2x4_ASAP7_75t_L g1443 ( .A(n_1440), .B(n_1444), .Y(n_1443) );
INVx2_ASAP7_75t_L g1446 ( .A(n_1447), .Y(n_1446) );
BUFx3_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
AND2x2_ASAP7_75t_L g1450 ( .A(n_1451), .B(n_1453), .Y(n_1450) );
INVx1_ASAP7_75t_SL g1451 ( .A(n_1452), .Y(n_1451) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
INVx2_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
INVxp33_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
HB1xp67_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
NAND3xp33_ASAP7_75t_L g1463 ( .A(n_1464), .B(n_1466), .C(n_1485), .Y(n_1463) );
AOI21xp5_ASAP7_75t_L g1466 ( .A1(n_1467), .A2(n_1468), .B(n_1483), .Y(n_1466) );
NAND3xp33_ASAP7_75t_L g1468 ( .A(n_1469), .B(n_1475), .C(n_1480), .Y(n_1468) );
NAND2xp5_ASAP7_75t_L g1486 ( .A(n_1487), .B(n_1488), .Y(n_1486) );
INVx1_ASAP7_75t_L g1494 ( .A(n_1495), .Y(n_1494) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
HB1xp67_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
BUFx3_ASAP7_75t_L g1497 ( .A(n_1498), .Y(n_1497) );
HB1xp67_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
OAI21xp5_ASAP7_75t_L g1500 ( .A1(n_1501), .A2(n_1502), .B(n_1503), .Y(n_1500) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
endmodule