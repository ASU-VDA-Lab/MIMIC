module fake_jpeg_2987_n_159 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_159);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_7),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_42),
.Y(n_54)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

OR2x2_ASAP7_75t_SL g69 ( 
.A(n_41),
.B(n_16),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_49),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_10),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_48),
.Y(n_57)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_13),
.B1(n_25),
.B2(n_19),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_13),
.Y(n_62)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_24),
.B1(n_30),
.B2(n_15),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_50),
.A2(n_61),
.B1(n_6),
.B2(n_63),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_27),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_53),
.B(n_59),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_23),
.B1(n_43),
.B2(n_40),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_76),
.B1(n_6),
.B2(n_11),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_28),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_34),
.A2(n_23),
.B1(n_28),
.B2(n_27),
.Y(n_61)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_63),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_31),
.B(n_14),
.C(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_64),
.B(n_66),
.Y(n_85)
);

AO22x1_ASAP7_75t_SL g65 ( 
.A1(n_47),
.A2(n_19),
.B1(n_14),
.B2(n_17),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_53),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_29),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_17),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_71),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_69),
.B(n_72),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_33),
.B(n_16),
.Y(n_71)
);

NOR2x1_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_32),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_10),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_54),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_36),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_86),
.B1(n_55),
.B2(n_51),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_84),
.A2(n_50),
.B1(n_65),
.B2(n_76),
.Y(n_102)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_90),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_95),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_64),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_68),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_68),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_86),
.B1(n_85),
.B2(n_80),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_102),
.B1(n_106),
.B2(n_103),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_61),
.B1(n_75),
.B2(n_72),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_103),
.A2(n_96),
.B1(n_97),
.B2(n_91),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_61),
.B1(n_55),
.B2(n_69),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_114),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_80),
.B(n_96),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_111),
.A2(n_112),
.B(n_83),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_96),
.A2(n_98),
.B(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_78),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_119),
.Y(n_138)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NOR3xp33_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_126),
.C(n_128),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_82),
.B1(n_92),
.B2(n_90),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_124),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_99),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_87),
.C(n_111),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_112),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_104),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

HAxp5_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_100),
.CON(n_128),
.SN(n_128)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_125),
.C(n_120),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_134),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_110),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_100),
.B(n_106),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_125),
.B(n_120),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_108),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_135),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_145),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_121),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_141),
.B(n_129),
.Y(n_147)
);

AO221x1_ASAP7_75t_L g142 ( 
.A1(n_136),
.A2(n_119),
.B1(n_115),
.B2(n_126),
.C(n_116),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_145),
.Y(n_150)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_144),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_143),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_140),
.C(n_132),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_152),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_146),
.A2(n_138),
.B1(n_133),
.B2(n_123),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_153),
.A2(n_154),
.B(n_148),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_105),
.A3(n_115),
.B1(n_117),
.B2(n_138),
.C1(n_134),
.C2(n_130),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_155),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_156),
.C(n_152),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);


endmodule