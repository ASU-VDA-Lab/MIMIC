module fake_ibex_1247_n_1588 (n_151, n_147, n_85, n_251, n_167, n_128, n_253, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_247, n_55, n_130, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_8, n_118, n_224, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_264, n_124, n_37, n_256, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_263, n_27, n_165, n_242, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_255, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_262, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_249, n_14, n_0, n_239, n_94, n_134, n_12, n_42, n_77, n_112, n_257, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_258, n_80, n_172, n_215, n_250, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_261, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_260, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_252, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_248, n_92, n_144, n_170, n_213, n_254, n_101, n_190, n_113, n_138, n_230, n_96, n_185, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_265, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_259, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_246, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1588);

input n_151;
input n_147;
input n_85;
input n_251;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_247;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_8;
input n_118;
input n_224;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_264;
input n_124;
input n_37;
input n_256;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_263;
input n_27;
input n_165;
input n_242;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_255;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_262;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_249;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_257;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_258;
input n_80;
input n_172;
input n_215;
input n_250;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_261;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_260;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_252;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_248;
input n_92;
input n_144;
input n_170;
input n_213;
input n_254;
input n_101;
input n_190;
input n_113;
input n_138;
input n_230;
input n_96;
input n_185;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_265;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_259;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_246;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1588;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_280;
wire n_375;
wire n_1391;
wire n_884;
wire n_667;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_1509;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1301;
wire n_869;
wire n_1561;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_562;
wire n_564;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_1506;
wire n_881;
wire n_734;
wire n_1558;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1531;
wire n_1332;
wire n_482;
wire n_282;
wire n_1424;
wire n_870;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_737;
wire n_606;
wire n_1571;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_1577;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_1568;
wire n_325;
wire n_1184;
wire n_1477;
wire n_1364;
wire n_1540;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1522;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_267;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_1545;
wire n_351;
wire n_456;
wire n_1471;
wire n_998;
wire n_1115;
wire n_1395;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1470;
wire n_444;
wire n_986;
wire n_495;
wire n_1420;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_1539;
wire n_712;
wire n_1400;
wire n_650;
wire n_409;
wire n_1575;
wire n_332;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_1439;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_318;
wire n_291;
wire n_268;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_303;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_266;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1560;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1497;
wire n_1578;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_1458;
wire n_1460;
wire n_326;
wire n_270;
wire n_1340;
wire n_339;
wire n_276;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_1491;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1587;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_269;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_1538;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_993;
wire n_851;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_1169;
wire n_571;
wire n_648;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_839;
wire n_768;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_1406;
wire n_1489;
wire n_804;
wire n_484;
wire n_1455;
wire n_480;
wire n_1057;
wire n_354;
wire n_1473;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_277;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1501;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_1513;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1221;
wire n_284;
wire n_1047;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1565;
wire n_1257;
wire n_274;
wire n_387;
wire n_688;
wire n_1542;
wire n_946;
wire n_1547;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_586;
wire n_1330;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1564;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_886;
wire n_383;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1161;
wire n_1103;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_335;
wire n_1499;
wire n_1500;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_305;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1536;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_537;
wire n_1113;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_271;
wire n_1393;
wire n_984;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_244),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_224),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_92),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_107),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_238),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_180),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_263),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_204),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_45),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_213),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_67),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_83),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_129),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_128),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_206),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_162),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_199),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_198),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_84),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_3),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_202),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_242),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_82),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_115),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_5),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_239),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_147),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_78),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_191),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_243),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_183),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_232),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_104),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_212),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_228),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_153),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_88),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_241),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_108),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_157),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_223),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_77),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_80),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_163),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_195),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_252),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_160),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_217),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_120),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_189),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_83),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_185),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_215),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_59),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_255),
.Y(n_320)
);

BUFx10_ASAP7_75t_L g321 ( 
.A(n_230),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_184),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_245),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_112),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_117),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_211),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_37),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_37),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_45),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_176),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_193),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_3),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_210),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_214),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_121),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_133),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_7),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_260),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_33),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_11),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_246),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_178),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_100),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_146),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_218),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_234),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_8),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_19),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_56),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_29),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_110),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_34),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_70),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_124),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_127),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_173),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_231),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_247),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_175),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_150),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_29),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_123),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_161),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_265),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_257),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_48),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_136),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_100),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_253),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_42),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_64),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_229),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_18),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_53),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_159),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_152),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_143),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_61),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_171),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_182),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_220),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_15),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_114),
.Y(n_383)
);

BUFx2_ASAP7_75t_SL g384 ( 
.A(n_30),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_38),
.Y(n_385)
);

INVxp33_ASAP7_75t_L g386 ( 
.A(n_181),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_240),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_256),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_87),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_32),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_33),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_236),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_42),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_21),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_118),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_20),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_145),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_158),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_87),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_119),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_86),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_84),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_137),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_135),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_172),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_219),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_16),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_85),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_207),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_151),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_101),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_166),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_258),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_10),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_122),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_155),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_51),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_65),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_138),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_40),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_235),
.Y(n_421)
);

CKINVDCx14_ASAP7_75t_R g422 ( 
.A(n_0),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_165),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_168),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_126),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_188),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_55),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_80),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_216),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_203),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_156),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_79),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_131),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_237),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_102),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_47),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_34),
.Y(n_437)
);

BUFx2_ASAP7_75t_SL g438 ( 
.A(n_30),
.Y(n_438)
);

BUFx5_ASAP7_75t_L g439 ( 
.A(n_141),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_144),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_130),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_197),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_149),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_4),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_8),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_174),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_262),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_31),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_140),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_225),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_90),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_54),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_62),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_41),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_1),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_57),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_177),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_69),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_192),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_63),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_22),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_264),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_116),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_233),
.Y(n_464)
);

BUFx10_ASAP7_75t_L g465 ( 
.A(n_179),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_125),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_248),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_154),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_113),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_249),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_49),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_91),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_41),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_26),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_164),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_55),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_289),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_339),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_266),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_339),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_269),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_299),
.B(n_2),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_439),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_422),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_349),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_279),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_349),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_371),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_269),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_448),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_448),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_315),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_399),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_437),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_455),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_268),
.Y(n_496)
);

BUFx6f_ASAP7_75t_SL g497 ( 
.A(n_321),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_304),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_444),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_461),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_451),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_299),
.B(n_4),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_472),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_436),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_329),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_436),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_276),
.Y(n_507)
);

NOR2xp67_ASAP7_75t_L g508 ( 
.A(n_293),
.B(n_307),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_328),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_332),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_318),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g512 ( 
.A(n_321),
.Y(n_512)
);

INVxp33_ASAP7_75t_SL g513 ( 
.A(n_268),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_456),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_340),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_330),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_368),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_370),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_274),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_374),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_362),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_364),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_369),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_385),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_274),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_389),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_277),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_377),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_400),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_439),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_405),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_394),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_407),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_418),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_277),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_428),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_458),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_473),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_413),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_284),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_284),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_474),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_271),
.B(n_6),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_465),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_285),
.Y(n_545)
);

NOR2xp67_ASAP7_75t_L g546 ( 
.A(n_273),
.B(n_6),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_465),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_291),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_285),
.Y(n_549)
);

INVxp67_ASAP7_75t_SL g550 ( 
.A(n_386),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_292),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_416),
.Y(n_552)
);

INVxp67_ASAP7_75t_SL g553 ( 
.A(n_282),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_297),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_439),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_439),
.Y(n_556)
);

INVxp67_ASAP7_75t_SL g557 ( 
.A(n_282),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_288),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_300),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_314),
.Y(n_560)
);

CKINVDCx16_ASAP7_75t_R g561 ( 
.A(n_421),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_325),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_288),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_326),
.B(n_7),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_331),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_R g566 ( 
.A(n_305),
.B(n_109),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_290),
.Y(n_567)
);

INVxp33_ASAP7_75t_L g568 ( 
.A(n_311),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_267),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_290),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_333),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_267),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_298),
.B(n_9),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_298),
.B(n_9),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_334),
.Y(n_575)
);

INVxp67_ASAP7_75t_SL g576 ( 
.A(n_294),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_335),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_346),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_302),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_354),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_356),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_302),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_270),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_411),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_357),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_483),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_483),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_530),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_478),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_530),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_480),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_485),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_550),
.B(n_411),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_487),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_555),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_490),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_555),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_556),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_491),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_504),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_506),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_568),
.B(n_414),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_496),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_SL g604 ( 
.A(n_497),
.B(n_568),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_582),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_544),
.B(n_341),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_484),
.B(n_414),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_499),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_513),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_547),
.B(n_341),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_497),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_481),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_477),
.B(n_360),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_489),
.B(n_360),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_507),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_503),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_548),
.B(n_311),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_551),
.Y(n_618)
);

OAI21x1_ASAP7_75t_L g619 ( 
.A1(n_554),
.A2(n_376),
.B(n_355),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_559),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_545),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_553),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_509),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_560),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_557),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_510),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_562),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_576),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_512),
.B(n_427),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_501),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_515),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_517),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_545),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_565),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_519),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_SL g636 ( 
.A(n_497),
.B(n_272),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_518),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_520),
.Y(n_638)
);

AND2x6_ASAP7_75t_L g639 ( 
.A(n_482),
.B(n_363),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_526),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_569),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_532),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_572),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_533),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_524),
.B(n_493),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_505),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_534),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_536),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_493),
.B(n_432),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_571),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_583),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_537),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_538),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_542),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_575),
.B(n_355),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_577),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_502),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_573),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_585),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_578),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_580),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_581),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_508),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_574),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_543),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_492),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_546),
.Y(n_667)
);

AOI22x1_ASAP7_75t_L g668 ( 
.A1(n_492),
.A2(n_433),
.B1(n_468),
.B2(n_376),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_564),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_566),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_494),
.B(n_471),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_494),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_479),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_519),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_525),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_525),
.B(n_471),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_527),
.Y(n_677)
);

BUFx8_ASAP7_75t_L g678 ( 
.A(n_527),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_535),
.Y(n_679)
);

OA21x2_ASAP7_75t_L g680 ( 
.A1(n_486),
.A2(n_468),
.B(n_433),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_535),
.B(n_363),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_540),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_540),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_541),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_541),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_498),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_549),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_511),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_549),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_558),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_558),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_563),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_563),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_567),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_567),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_516),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_570),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_570),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_579),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_579),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_584),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_584),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_521),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_488),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_522),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_523),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_528),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_529),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_531),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_539),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_552),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_561),
.B(n_278),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_488),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_495),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_495),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_500),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_500),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_505),
.B(n_358),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_514),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_514),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_L g721 ( 
.A(n_569),
.B(n_439),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_478),
.Y(n_722)
);

XOR2xp5_ASAP7_75t_L g723 ( 
.A(n_488),
.B(n_308),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_513),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_483),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_478),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_483),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_478),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_496),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_483),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_550),
.B(n_278),
.Y(n_731)
);

BUFx2_ASAP7_75t_L g732 ( 
.A(n_545),
.Y(n_732)
);

OA21x2_ASAP7_75t_L g733 ( 
.A1(n_483),
.A2(n_367),
.B(n_365),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_513),
.A2(n_319),
.B1(n_327),
.B2(n_316),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_483),
.Y(n_735)
);

BUFx2_ASAP7_75t_L g736 ( 
.A(n_545),
.Y(n_736)
);

BUFx8_ASAP7_75t_L g737 ( 
.A(n_497),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_483),
.Y(n_738)
);

NAND2xp33_ASAP7_75t_SL g739 ( 
.A(n_497),
.B(n_280),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_513),
.A2(n_476),
.B1(n_337),
.B2(n_343),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_548),
.B(n_439),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_496),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_478),
.B(n_372),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_478),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_483),
.Y(n_745)
);

INVx4_ASAP7_75t_L g746 ( 
.A(n_497),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_483),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_478),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_483),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_550),
.B(n_281),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_483),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_478),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_478),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_483),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_548),
.B(n_439),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_478),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_608),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_731),
.B(n_281),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_669),
.B(n_380),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_653),
.B(n_283),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_596),
.Y(n_761)
);

AND2x6_ASAP7_75t_L g762 ( 
.A(n_743),
.B(n_387),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_608),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_596),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_645),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_669),
.B(n_397),
.Y(n_766)
);

NAND2x1p5_ASAP7_75t_L g767 ( 
.A(n_611),
.B(n_417),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_726),
.Y(n_768)
);

INVx5_ASAP7_75t_L g769 ( 
.A(n_586),
.Y(n_769)
);

INVx4_ASAP7_75t_L g770 ( 
.A(n_611),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_726),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_746),
.B(n_420),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_608),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_728),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_728),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_608),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_635),
.B(n_384),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_L g778 ( 
.A(n_639),
.B(n_439),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_748),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_602),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_669),
.B(n_403),
.Y(n_781)
);

INVx4_ASAP7_75t_L g782 ( 
.A(n_746),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_750),
.B(n_286),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_619),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_669),
.B(n_404),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_752),
.Y(n_786)
);

AND3x4_ASAP7_75t_L g787 ( 
.A(n_718),
.B(n_438),
.C(n_348),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_657),
.B(n_287),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_613),
.B(n_347),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_613),
.B(n_350),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_658),
.A2(n_353),
.B1(n_361),
.B2(n_352),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_613),
.B(n_366),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_612),
.B(n_287),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_658),
.B(n_664),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_587),
.B(n_410),
.Y(n_795)
);

INVx4_ASAP7_75t_L g796 ( 
.A(n_618),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_587),
.B(n_423),
.Y(n_797)
);

INVx5_ASAP7_75t_L g798 ( 
.A(n_586),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_588),
.B(n_424),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_756),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_756),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_616),
.B(n_295),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_605),
.B(n_373),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_737),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_589),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_618),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_618),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_737),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_664),
.B(n_295),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_622),
.B(n_296),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_620),
.Y(n_811)
);

AO21x2_ASAP7_75t_L g812 ( 
.A1(n_619),
.A2(n_431),
.B(n_426),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_743),
.B(n_378),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_620),
.Y(n_814)
);

INVxp67_ASAP7_75t_SL g815 ( 
.A(n_615),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_656),
.B(n_296),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_591),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_625),
.B(n_301),
.Y(n_818)
);

OR2x6_ASAP7_75t_L g819 ( 
.A(n_686),
.B(n_441),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_628),
.B(n_301),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_678),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_743),
.B(n_630),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_609),
.Y(n_823)
);

BUFx10_ASAP7_75t_L g824 ( 
.A(n_609),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_732),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_593),
.B(n_303),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_605),
.B(n_382),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_624),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_656),
.B(n_303),
.Y(n_829)
);

INVx4_ASAP7_75t_L g830 ( 
.A(n_624),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_631),
.A2(n_391),
.B1(n_393),
.B2(n_390),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_659),
.B(n_412),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_729),
.B(n_396),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_592),
.Y(n_834)
);

AND2x2_ASAP7_75t_SL g835 ( 
.A(n_736),
.B(n_449),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_729),
.B(n_401),
.Y(n_836)
);

BUFx4f_ASAP7_75t_L g837 ( 
.A(n_686),
.Y(n_837)
);

AND2x6_ASAP7_75t_L g838 ( 
.A(n_681),
.B(n_462),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_594),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_607),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_599),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_722),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_588),
.B(n_463),
.Y(n_843)
);

BUFx4f_ASAP7_75t_L g844 ( 
.A(n_686),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_742),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_627),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_672),
.B(n_402),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_627),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_672),
.B(n_408),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_627),
.Y(n_850)
);

NAND2xp33_ASAP7_75t_L g851 ( 
.A(n_639),
.B(n_419),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_665),
.B(n_419),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_SL g853 ( 
.A(n_724),
.B(n_425),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_634),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_659),
.B(n_425),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_665),
.B(n_430),
.Y(n_856)
);

INVx4_ASAP7_75t_L g857 ( 
.A(n_634),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_733),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_662),
.B(n_430),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_621),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_681),
.B(n_435),
.Y(n_861)
);

AO22x2_ASAP7_75t_L g862 ( 
.A1(n_718),
.A2(n_470),
.B1(n_409),
.B2(n_306),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_744),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_650),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_629),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_650),
.Y(n_866)
);

AND2x6_ASAP7_75t_L g867 ( 
.A(n_681),
.B(n_312),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_662),
.B(n_466),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_661),
.B(n_466),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_650),
.Y(n_870)
);

OAI22xp33_ASAP7_75t_L g871 ( 
.A1(n_674),
.A2(n_452),
.B1(n_453),
.B2(n_445),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_660),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_615),
.A2(n_312),
.B1(n_450),
.B2(n_429),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_660),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_688),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_606),
.B(n_454),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_R g877 ( 
.A(n_636),
.B(n_467),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_606),
.B(n_460),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_688),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_688),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_753),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_733),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_600),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_621),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_610),
.B(n_469),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_733),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_623),
.B(n_475),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_603),
.B(n_475),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_633),
.B(n_275),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_590),
.B(n_312),
.Y(n_890)
);

OR2x2_ASAP7_75t_L g891 ( 
.A(n_676),
.B(n_12),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_623),
.B(n_309),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_633),
.B(n_359),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_586),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_678),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_626),
.B(n_637),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_610),
.B(n_381),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_600),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_626),
.A2(n_450),
.B1(n_429),
.B2(n_415),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_601),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_688),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_637),
.B(n_310),
.Y(n_902)
);

NAND2xp33_ASAP7_75t_L g903 ( 
.A(n_639),
.B(n_313),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_638),
.B(n_317),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_641),
.B(n_464),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_595),
.B(n_597),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_638),
.B(n_320),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_696),
.Y(n_908)
);

NAND2xp33_ASAP7_75t_L g909 ( 
.A(n_639),
.B(n_459),
.Y(n_909)
);

BUFx8_ASAP7_75t_SL g910 ( 
.A(n_646),
.Y(n_910)
);

AO22x2_ASAP7_75t_L g911 ( 
.A1(n_787),
.A2(n_723),
.B1(n_719),
.B2(n_720),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_910),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_845),
.A2(n_765),
.B1(n_794),
.B2(n_860),
.Y(n_913)
);

AO22x2_ASAP7_75t_L g914 ( 
.A1(n_787),
.A2(n_791),
.B1(n_862),
.B2(n_861),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_794),
.B(n_666),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_780),
.B(n_610),
.Y(n_916)
);

OAI221xp5_ASAP7_75t_L g917 ( 
.A1(n_865),
.A2(n_734),
.B1(n_671),
.B2(n_674),
.C(n_685),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_805),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_884),
.B(n_641),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_817),
.Y(n_920)
);

OAI221xp5_ASAP7_75t_L g921 ( 
.A1(n_840),
.A2(n_685),
.B1(n_697),
.B2(n_692),
.C(n_679),
.Y(n_921)
);

AO22x2_ASAP7_75t_L g922 ( 
.A1(n_791),
.A2(n_719),
.B1(n_692),
.B2(n_697),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_860),
.B(n_666),
.Y(n_923)
);

OAI221xp5_ASAP7_75t_L g924 ( 
.A1(n_809),
.A2(n_679),
.B1(n_698),
.B2(n_649),
.C(n_740),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_825),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_809),
.B(n_614),
.Y(n_926)
);

NAND3xp33_ASAP7_75t_SL g927 ( 
.A(n_853),
.B(n_691),
.C(n_675),
.Y(n_927)
);

NAND2xp33_ASAP7_75t_L g928 ( 
.A(n_762),
.B(n_604),
.Y(n_928)
);

AO22x2_ASAP7_75t_L g929 ( 
.A1(n_862),
.A2(n_698),
.B1(n_682),
.B2(n_683),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_834),
.Y(n_930)
);

OR2x6_ASAP7_75t_L g931 ( 
.A(n_808),
.B(n_714),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_813),
.B(n_643),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_839),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_804),
.B(n_712),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_852),
.B(n_856),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_822),
.B(n_651),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_841),
.Y(n_937)
);

NAND2xp33_ASAP7_75t_L g938 ( 
.A(n_762),
.B(n_739),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_842),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_823),
.Y(n_940)
);

AO22x2_ASAP7_75t_L g941 ( 
.A1(n_862),
.A2(n_684),
.B1(n_687),
.B2(n_677),
.Y(n_941)
);

NAND2x1p5_ASAP7_75t_L g942 ( 
.A(n_770),
.B(n_782),
.Y(n_942)
);

AO22x2_ASAP7_75t_L g943 ( 
.A1(n_861),
.A2(n_689),
.B1(n_693),
.B2(n_690),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_869),
.B(n_632),
.Y(n_944)
);

AO22x2_ASAP7_75t_L g945 ( 
.A1(n_885),
.A2(n_694),
.B1(n_700),
.B2(n_699),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_863),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_786),
.Y(n_947)
);

XOR2x2_ASAP7_75t_L g948 ( 
.A(n_835),
.B(n_695),
.Y(n_948)
);

AO22x2_ASAP7_75t_L g949 ( 
.A1(n_885),
.A2(n_702),
.B1(n_717),
.B2(n_704),
.Y(n_949)
);

CKINVDCx16_ASAP7_75t_R g950 ( 
.A(n_824),
.Y(n_950)
);

AO22x2_ASAP7_75t_L g951 ( 
.A1(n_831),
.A2(n_713),
.B1(n_716),
.B2(n_715),
.Y(n_951)
);

AO22x2_ASAP7_75t_L g952 ( 
.A1(n_813),
.A2(n_678),
.B1(n_646),
.B2(n_673),
.Y(n_952)
);

AO22x2_ASAP7_75t_L g953 ( 
.A1(n_789),
.A2(n_706),
.B1(n_710),
.B2(n_703),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_803),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_883),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_883),
.Y(n_956)
);

AO22x2_ASAP7_75t_L g957 ( 
.A1(n_789),
.A2(n_792),
.B1(n_790),
.B2(n_876),
.Y(n_957)
);

NOR2xp67_ASAP7_75t_L g958 ( 
.A(n_821),
.B(n_707),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_881),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_900),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_815),
.B(n_640),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_867),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_815),
.Y(n_963)
);

AND2x6_ASAP7_75t_SL g964 ( 
.A(n_895),
.B(n_711),
.Y(n_964)
);

AO22x2_ASAP7_75t_L g965 ( 
.A1(n_790),
.A2(n_667),
.B1(n_701),
.B2(n_695),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_900),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_838),
.A2(n_680),
.B1(n_670),
.B2(n_642),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_896),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_SL g969 ( 
.A1(n_838),
.A2(n_701),
.B1(n_714),
.B2(n_708),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_761),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_764),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_768),
.Y(n_972)
);

AO22x2_ASAP7_75t_L g973 ( 
.A1(n_792),
.A2(n_680),
.B1(n_663),
.B2(n_714),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_771),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_838),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_774),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_782),
.Y(n_977)
);

BUFx6f_ASAP7_75t_SL g978 ( 
.A(n_824),
.Y(n_978)
);

CKINVDCx20_ASAP7_75t_R g979 ( 
.A(n_877),
.Y(n_979)
);

AND2x6_ASAP7_75t_L g980 ( 
.A(n_878),
.B(n_705),
.Y(n_980)
);

AO22x2_ASAP7_75t_L g981 ( 
.A1(n_878),
.A2(n_655),
.B1(n_617),
.B2(n_647),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_775),
.Y(n_982)
);

NAND2x1p5_ASAP7_75t_L g983 ( 
.A(n_837),
.B(n_705),
.Y(n_983)
);

AND2x2_ASAP7_75t_SL g984 ( 
.A(n_837),
.B(n_705),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_779),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_800),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_801),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_898),
.Y(n_988)
);

NAND3xp33_ASAP7_75t_L g989 ( 
.A(n_826),
.B(n_721),
.C(n_668),
.Y(n_989)
);

AO22x2_ASAP7_75t_L g990 ( 
.A1(n_847),
.A2(n_617),
.B1(n_647),
.B2(n_644),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_847),
.B(n_705),
.Y(n_991)
);

AO22x2_ASAP7_75t_L g992 ( 
.A1(n_849),
.A2(n_827),
.B1(n_836),
.B2(n_833),
.Y(n_992)
);

INVxp67_ASAP7_75t_L g993 ( 
.A(n_888),
.Y(n_993)
);

BUFx8_ASAP7_75t_L g994 ( 
.A(n_867),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_760),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_772),
.B(n_708),
.Y(n_996)
);

AO22x2_ASAP7_75t_L g997 ( 
.A1(n_849),
.A2(n_654),
.B1(n_648),
.B2(n_652),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_826),
.B(n_648),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_891),
.B(n_709),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_877),
.Y(n_1000)
);

AO22x2_ASAP7_75t_L g1001 ( 
.A1(n_777),
.A2(n_654),
.B1(n_709),
.B2(n_741),
.Y(n_1001)
);

AO22x2_ASAP7_75t_L g1002 ( 
.A1(n_889),
.A2(n_709),
.B1(n_755),
.B2(n_14),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_796),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_816),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_829),
.Y(n_1005)
);

NAND2x1p5_ASAP7_75t_L g1006 ( 
.A(n_844),
.B(n_598),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_875),
.B(n_13),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_788),
.B(n_758),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_879),
.B(n_880),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_901),
.B(n_14),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_814),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_SL g1012 ( 
.A1(n_767),
.A2(n_323),
.B1(n_324),
.B2(n_322),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_832),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_893),
.B(n_727),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_830),
.Y(n_1015)
);

NAND2x1p5_ASAP7_75t_L g1016 ( 
.A(n_844),
.B(n_735),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_855),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_855),
.Y(n_1018)
);

INVxp67_ASAP7_75t_L g1019 ( 
.A(n_905),
.Y(n_1019)
);

AO22x2_ASAP7_75t_L g1020 ( 
.A1(n_859),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_1020)
);

AO22x2_ASAP7_75t_L g1021 ( 
.A1(n_859),
.A2(n_22),
.B1(n_17),
.B2(n_20),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_762),
.A2(n_747),
.B1(n_745),
.B2(n_754),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_793),
.B(n_23),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_867),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_908),
.B(n_24),
.Y(n_1025)
);

NAND2x1p5_ASAP7_75t_L g1026 ( 
.A(n_769),
.B(n_725),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_868),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_819),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_867),
.Y(n_1029)
);

AO22x2_ASAP7_75t_L g1030 ( 
.A1(n_887),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_1030)
);

AO22x2_ASAP7_75t_L g1031 ( 
.A1(n_759),
.A2(n_28),
.B1(n_25),
.B2(n_27),
.Y(n_1031)
);

AO22x2_ASAP7_75t_L g1032 ( 
.A1(n_759),
.A2(n_31),
.B1(n_27),
.B2(n_28),
.Y(n_1032)
);

AO22x2_ASAP7_75t_L g1033 ( 
.A1(n_766),
.A2(n_785),
.B1(n_781),
.B2(n_795),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_797),
.Y(n_1034)
);

AO22x2_ASAP7_75t_L g1035 ( 
.A1(n_766),
.A2(n_36),
.B1(n_32),
.B2(n_35),
.Y(n_1035)
);

OAI221xp5_ASAP7_75t_L g1036 ( 
.A1(n_802),
.A2(n_406),
.B1(n_338),
.B2(n_342),
.C(n_344),
.Y(n_1036)
);

AO22x2_ASAP7_75t_L g1037 ( 
.A1(n_781),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_1037)
);

NOR3xp33_ASAP7_75t_L g1038 ( 
.A(n_871),
.B(n_345),
.C(n_336),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_858),
.Y(n_1039)
);

INVxp33_ASAP7_75t_SL g1040 ( 
.A(n_783),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_897),
.A2(n_751),
.B(n_749),
.C(n_738),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_968),
.B(n_858),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_1039),
.B(n_882),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_915),
.B(n_810),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_913),
.B(n_810),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_967),
.B(n_886),
.Y(n_1046)
);

XNOR2x2_ASAP7_75t_L g1047 ( 
.A(n_914),
.B(n_897),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_1028),
.B(n_871),
.Y(n_1048)
);

NAND2xp33_ASAP7_75t_SL g1049 ( 
.A(n_975),
.B(n_886),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_923),
.B(n_892),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_940),
.B(n_902),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_936),
.B(n_902),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_1040),
.B(n_904),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_919),
.B(n_907),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_925),
.B(n_907),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_1012),
.B(n_818),
.Y(n_1056)
);

NAND2xp33_ASAP7_75t_SL g1057 ( 
.A(n_979),
.B(n_784),
.Y(n_1057)
);

NAND2xp33_ASAP7_75t_SL g1058 ( 
.A(n_962),
.B(n_784),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_950),
.B(n_818),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_969),
.B(n_820),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_916),
.B(n_769),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_1000),
.B(n_1019),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_963),
.B(n_769),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_932),
.B(n_785),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_961),
.B(n_769),
.Y(n_1065)
);

NAND2xp33_ASAP7_75t_SL g1066 ( 
.A(n_1024),
.B(n_857),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1014),
.B(n_799),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_984),
.B(n_798),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_995),
.B(n_799),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_994),
.B(n_899),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_934),
.B(n_857),
.Y(n_1071)
);

NAND2xp33_ASAP7_75t_SL g1072 ( 
.A(n_1029),
.B(n_843),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_958),
.B(n_351),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_993),
.B(n_375),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_1007),
.B(n_379),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_1007),
.B(n_383),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_1010),
.B(n_388),
.Y(n_1077)
);

NAND2xp33_ASAP7_75t_SL g1078 ( 
.A(n_978),
.B(n_851),
.Y(n_1078)
);

NAND2xp33_ASAP7_75t_SL g1079 ( 
.A(n_926),
.B(n_812),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_1010),
.B(n_392),
.Y(n_1080)
);

NAND2xp33_ASAP7_75t_SL g1081 ( 
.A(n_1008),
.B(n_812),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_1025),
.B(n_395),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_954),
.B(n_906),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_1025),
.B(n_398),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_991),
.B(n_434),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_991),
.B(n_440),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_1009),
.B(n_442),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_1009),
.B(n_443),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1004),
.B(n_903),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_999),
.B(n_446),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_918),
.B(n_806),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1005),
.B(n_909),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_999),
.B(n_447),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_942),
.B(n_1038),
.Y(n_1094)
);

NAND2xp33_ASAP7_75t_SL g1095 ( 
.A(n_944),
.B(n_846),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1013),
.B(n_778),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_1017),
.B(n_457),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1018),
.B(n_806),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1027),
.B(n_854),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_920),
.B(n_854),
.Y(n_1100)
);

NAND2xp33_ASAP7_75t_SL g1101 ( 
.A(n_935),
.B(n_763),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_930),
.B(n_866),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_933),
.B(n_866),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_998),
.B(n_1022),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_937),
.B(n_870),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_939),
.B(n_870),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_1006),
.B(n_894),
.Y(n_1107)
);

NAND2xp33_ASAP7_75t_SL g1108 ( 
.A(n_1023),
.B(n_763),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_1016),
.B(n_872),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_977),
.B(n_872),
.Y(n_1110)
);

NAND2xp33_ASAP7_75t_SL g1111 ( 
.A(n_914),
.B(n_873),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_983),
.B(n_730),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_946),
.B(n_807),
.Y(n_1113)
);

AND2x2_ASAP7_75t_SL g1114 ( 
.A(n_928),
.B(n_938),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_959),
.B(n_811),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_992),
.B(n_39),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_948),
.B(n_828),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_970),
.B(n_757),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_992),
.B(n_40),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_957),
.B(n_911),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_997),
.B(n_957),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_988),
.B(n_848),
.Y(n_1122)
);

NAND2xp33_ASAP7_75t_SL g1123 ( 
.A(n_912),
.B(n_890),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_996),
.B(n_850),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_924),
.B(n_864),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_974),
.B(n_773),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_911),
.B(n_952),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_1003),
.B(n_874),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_953),
.B(n_776),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_952),
.B(n_43),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_953),
.B(n_43),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1011),
.B(n_44),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_1015),
.B(n_44),
.Y(n_1133)
);

XNOR2xp5_ASAP7_75t_L g1134 ( 
.A(n_941),
.B(n_46),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_976),
.B(n_48),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_989),
.B(n_49),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_971),
.B(n_50),
.Y(n_1137)
);

NAND2xp33_ASAP7_75t_SL g1138 ( 
.A(n_947),
.B(n_50),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_972),
.B(n_51),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_955),
.B(n_52),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_956),
.B(n_53),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_960),
.B(n_54),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_922),
.B(n_56),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_966),
.B(n_57),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1026),
.B(n_58),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_982),
.B(n_59),
.Y(n_1146)
);

NAND2xp33_ASAP7_75t_SL g1147 ( 
.A(n_929),
.B(n_60),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_985),
.B(n_60),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_986),
.B(n_61),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_987),
.B(n_62),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_931),
.B(n_1034),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_951),
.B(n_66),
.Y(n_1152)
);

XNOR2x2_ASAP7_75t_L g1153 ( 
.A(n_941),
.B(n_67),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_927),
.B(n_68),
.Y(n_1154)
);

NAND2xp33_ASAP7_75t_SL g1155 ( 
.A(n_973),
.B(n_68),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1041),
.B(n_70),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_980),
.B(n_71),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_980),
.B(n_72),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_949),
.B(n_72),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_949),
.B(n_73),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_981),
.B(n_74),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_945),
.B(n_75),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_921),
.B(n_76),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_943),
.B(n_81),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_945),
.B(n_81),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_943),
.B(n_85),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1033),
.B(n_990),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_981),
.B(n_86),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1033),
.B(n_111),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_965),
.B(n_931),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_965),
.B(n_88),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1044),
.A2(n_917),
.B(n_1036),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1045),
.B(n_990),
.Y(n_1173)
);

INVx3_ASAP7_75t_SL g1174 ( 
.A(n_1062),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1081),
.A2(n_1001),
.B(n_1002),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1135),
.Y(n_1176)
);

INVxp67_ASAP7_75t_SL g1177 ( 
.A(n_1135),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_SL g1178 ( 
.A1(n_1134),
.A2(n_1127),
.B(n_1130),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1135),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1042),
.A2(n_1001),
.B(n_1002),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1042),
.A2(n_1030),
.B(n_1021),
.Y(n_1181)
);

O2A1O1Ixp5_ASAP7_75t_L g1182 ( 
.A1(n_1156),
.A2(n_1030),
.B(n_1020),
.C(n_1021),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1064),
.B(n_1020),
.Y(n_1183)
);

OA21x2_ASAP7_75t_L g1184 ( 
.A1(n_1046),
.A2(n_1037),
.B(n_1035),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1050),
.A2(n_1037),
.B(n_1035),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_1143),
.A2(n_1032),
.A3(n_1031),
.B(n_91),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_1091),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1147),
.A2(n_1032),
.B(n_1031),
.C(n_964),
.Y(n_1188)
);

AO21x1_ASAP7_75t_L g1189 ( 
.A1(n_1111),
.A2(n_89),
.B(n_92),
.Y(n_1189)
);

CKINVDCx11_ASAP7_75t_R g1190 ( 
.A(n_1151),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1123),
.B(n_93),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1083),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1171),
.B(n_93),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_SL g1194 ( 
.A1(n_1121),
.A2(n_1153),
.B(n_1047),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1114),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1117),
.B(n_94),
.Y(n_1196)
);

AOI221x1_ASAP7_75t_L g1197 ( 
.A1(n_1079),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.C(n_97),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1113),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1120),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1054),
.B(n_98),
.Y(n_1200)
);

INVx3_ASAP7_75t_SL g1201 ( 
.A(n_1071),
.Y(n_1201)
);

NAND2x1_ASAP7_75t_SL g1202 ( 
.A(n_1116),
.B(n_99),
.Y(n_1202)
);

NAND3xp33_ASAP7_75t_L g1203 ( 
.A(n_1154),
.B(n_102),
.C(n_103),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1089),
.A2(n_1092),
.B(n_1163),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1094),
.B(n_103),
.Y(n_1205)
);

NOR3xp33_ASAP7_75t_SL g1206 ( 
.A(n_1078),
.B(n_104),
.C(n_105),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1115),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1131),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1104),
.A2(n_105),
.B(n_106),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1170),
.B(n_1075),
.Y(n_1210)
);

AND3x4_ASAP7_75t_L g1211 ( 
.A(n_1151),
.B(n_106),
.C(n_107),
.Y(n_1211)
);

OR2x2_ASAP7_75t_L g1212 ( 
.A(n_1053),
.B(n_1059),
.Y(n_1212)
);

BUFx10_ASAP7_75t_L g1213 ( 
.A(n_1151),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1076),
.B(n_132),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1118),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_SL g1216 ( 
.A(n_1162),
.B(n_134),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_1077),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_1161),
.A2(n_139),
.A3(n_142),
.B(n_148),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_1165),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1119),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1164),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_1168),
.A2(n_167),
.A3(n_169),
.B(n_170),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1152),
.B(n_1051),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1080),
.B(n_186),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1125),
.A2(n_187),
.A3(n_190),
.B(n_194),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1069),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1114),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1056),
.B(n_196),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1166),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1146),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1052),
.B(n_200),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1048),
.B(n_201),
.Y(n_1232)
);

AO31x2_ASAP7_75t_L g1233 ( 
.A1(n_1129),
.A2(n_205),
.A3(n_208),
.B(n_209),
.Y(n_1233)
);

BUFx8_ASAP7_75t_L g1234 ( 
.A(n_1091),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_1082),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1167),
.A2(n_221),
.B1(n_222),
.B2(n_226),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1096),
.A2(n_1060),
.B(n_1067),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1055),
.B(n_227),
.Y(n_1238)
);

BUFx2_ASAP7_75t_SL g1239 ( 
.A(n_1084),
.Y(n_1239)
);

NAND2x1p5_ASAP7_75t_L g1240 ( 
.A(n_1160),
.B(n_261),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1085),
.B(n_1086),
.Y(n_1241)
);

BUFx10_ASAP7_75t_L g1242 ( 
.A(n_1091),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_1087),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1043),
.A2(n_250),
.B(n_251),
.Y(n_1244)
);

AO31x2_ASAP7_75t_L g1245 ( 
.A1(n_1098),
.A2(n_254),
.A3(n_259),
.B(n_1099),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1148),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_SL g1247 ( 
.A(n_1070),
.B(n_1057),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_SL g1248 ( 
.A1(n_1169),
.A2(n_1158),
.B(n_1157),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_1088),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1097),
.B(n_1090),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_1138),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1149),
.Y(n_1252)
);

AO31x2_ASAP7_75t_L g1253 ( 
.A1(n_1100),
.A2(n_1105),
.A3(n_1102),
.B(n_1106),
.Y(n_1253)
);

NAND3xp33_ASAP7_75t_SL g1254 ( 
.A(n_1073),
.B(n_1150),
.C(n_1093),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1137),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1066),
.B(n_1103),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1103),
.B(n_1072),
.Y(n_1257)
);

AO31x2_ASAP7_75t_L g1258 ( 
.A1(n_1101),
.A2(n_1108),
.A3(n_1136),
.B(n_1095),
.Y(n_1258)
);

O2A1O1Ixp33_ASAP7_75t_SL g1259 ( 
.A1(n_1065),
.A2(n_1107),
.B(n_1068),
.C(n_1139),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1074),
.B(n_1126),
.Y(n_1260)
);

CKINVDCx16_ASAP7_75t_R g1261 ( 
.A(n_1049),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1061),
.B(n_1126),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1132),
.B(n_1133),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_1058),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1063),
.Y(n_1265)
);

AOI221xp5_ASAP7_75t_L g1266 ( 
.A1(n_1140),
.A2(n_1144),
.B1(n_1142),
.B2(n_1141),
.C(n_1145),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1110),
.B(n_1124),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_SL g1268 ( 
.A(n_1109),
.B(n_1112),
.Y(n_1268)
);

AO32x2_ASAP7_75t_L g1269 ( 
.A1(n_1122),
.A2(n_1047),
.A3(n_1153),
.B1(n_1167),
.B2(n_1155),
.Y(n_1269)
);

INVx5_ASAP7_75t_L g1270 ( 
.A(n_1128),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1198),
.Y(n_1271)
);

OAI222xp33_ASAP7_75t_L g1272 ( 
.A1(n_1177),
.A2(n_1219),
.B1(n_1183),
.B2(n_1229),
.C1(n_1221),
.C2(n_1205),
.Y(n_1272)
);

AOI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1211),
.A2(n_1223),
.B1(n_1178),
.B2(n_1193),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1182),
.A2(n_1172),
.B(n_1173),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1198),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1216),
.B(n_1205),
.Y(n_1276)
);

INVx2_ASAP7_75t_SL g1277 ( 
.A(n_1234),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1220),
.B(n_1174),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1208),
.A2(n_1185),
.B1(n_1194),
.B2(n_1252),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1188),
.A2(n_1207),
.B1(n_1251),
.B2(n_1175),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1243),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1226),
.B(n_1207),
.Y(n_1282)
);

INVx2_ASAP7_75t_SL g1283 ( 
.A(n_1234),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_SL g1284 ( 
.A1(n_1191),
.A2(n_1247),
.B(n_1256),
.C(n_1209),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1244),
.A2(n_1180),
.B(n_1181),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1192),
.B(n_1190),
.Y(n_1286)
);

OAI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1196),
.A2(n_1197),
.B1(n_1176),
.B2(n_1179),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1264),
.Y(n_1288)
);

A2O1A1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1206),
.A2(n_1228),
.B(n_1232),
.C(n_1202),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1230),
.A2(n_1246),
.B1(n_1254),
.B2(n_1239),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1226),
.B(n_1237),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1249),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1255),
.A2(n_1189),
.B1(n_1227),
.B2(n_1195),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1253),
.B(n_1204),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1212),
.B(n_1210),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1201),
.Y(n_1296)
);

OR2x6_ASAP7_75t_L g1297 ( 
.A(n_1248),
.B(n_1195),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1217),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1200),
.Y(n_1299)
);

AO21x1_ASAP7_75t_L g1300 ( 
.A1(n_1240),
.A2(n_1236),
.B(n_1257),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1235),
.B(n_1241),
.Y(n_1301)
);

O2A1O1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1203),
.A2(n_1260),
.B(n_1250),
.C(n_1199),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1263),
.A2(n_1184),
.B(n_1266),
.Y(n_1303)
);

OR2x6_ASAP7_75t_L g1304 ( 
.A(n_1195),
.B(n_1227),
.Y(n_1304)
);

INVxp67_ASAP7_75t_L g1305 ( 
.A(n_1238),
.Y(n_1305)
);

OR2x6_ASAP7_75t_L g1306 ( 
.A(n_1227),
.B(n_1238),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1262),
.A2(n_1184),
.B1(n_1187),
.B2(n_1215),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1213),
.B(n_1265),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1213),
.A2(n_1267),
.B1(n_1214),
.B2(n_1224),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1242),
.B(n_1231),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1242),
.Y(n_1311)
);

OR2x6_ASAP7_75t_L g1312 ( 
.A(n_1261),
.B(n_1269),
.Y(n_1312)
);

BUFx2_ASAP7_75t_R g1313 ( 
.A(n_1269),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1270),
.A2(n_1268),
.B1(n_1186),
.B2(n_1259),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1258),
.B(n_1245),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1270),
.Y(n_1316)
);

A2O1A1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1218),
.A2(n_1222),
.B(n_1225),
.C(n_1245),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1218),
.B(n_1222),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1222),
.Y(n_1319)
);

AOI21xp33_ASAP7_75t_L g1320 ( 
.A1(n_1258),
.A2(n_1225),
.B(n_1233),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1225),
.A2(n_1127),
.B1(n_914),
.B2(n_911),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1211),
.A2(n_914),
.B1(n_915),
.B2(n_1040),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1219),
.B(n_1220),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1192),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_1190),
.Y(n_1325)
);

O2A1O1Ixp33_ASAP7_75t_SL g1326 ( 
.A1(n_1188),
.A2(n_1159),
.B(n_1160),
.C(n_1191),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1177),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1242),
.Y(n_1328)
);

INVx6_ASAP7_75t_L g1329 ( 
.A(n_1234),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1192),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1219),
.B(n_1220),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1177),
.B(n_1187),
.Y(n_1332)
);

BUFx8_ASAP7_75t_SL g1333 ( 
.A(n_1243),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1192),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1177),
.A2(n_914),
.B1(n_1188),
.B2(n_929),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1242),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1177),
.B(n_1187),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1226),
.B(n_1198),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1271),
.B(n_1275),
.Y(n_1339)
);

OA21x2_ASAP7_75t_L g1340 ( 
.A1(n_1317),
.A2(n_1320),
.B(n_1315),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1327),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1324),
.B(n_1330),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1327),
.Y(n_1343)
);

INVxp67_ASAP7_75t_L g1344 ( 
.A(n_1296),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1294),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1297),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1285),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1294),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1338),
.B(n_1282),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1322),
.A2(n_1335),
.B1(n_1273),
.B2(n_1280),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1311),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1334),
.B(n_1274),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1282),
.Y(n_1353)
);

NAND4xp25_ASAP7_75t_L g1354 ( 
.A(n_1321),
.B(n_1279),
.C(n_1335),
.D(n_1280),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1291),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1311),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1274),
.B(n_1307),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1291),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1305),
.B(n_1303),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1318),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1319),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1312),
.B(n_1299),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1297),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_1276),
.Y(n_1364)
);

OR2x6_ASAP7_75t_L g1365 ( 
.A(n_1312),
.B(n_1306),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1311),
.Y(n_1366)
);

INVx2_ASAP7_75t_SL g1367 ( 
.A(n_1329),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_SL g1368 ( 
.A(n_1305),
.B(n_1272),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1332),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1312),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1297),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1320),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1313),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1306),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1313),
.B(n_1337),
.Y(n_1375)
);

AO21x1_ASAP7_75t_SL g1376 ( 
.A1(n_1314),
.A2(n_1272),
.B(n_1293),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_L g1377 ( 
.A(n_1351),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_R g1378 ( 
.A(n_1367),
.B(n_1325),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1341),
.B(n_1304),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1339),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1342),
.B(n_1286),
.Y(n_1381)
);

XNOR2xp5_ASAP7_75t_L g1382 ( 
.A(n_1367),
.B(n_1281),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1353),
.B(n_1323),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1342),
.B(n_1301),
.Y(n_1384)
);

INVxp67_ASAP7_75t_L g1385 ( 
.A(n_1343),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1339),
.Y(n_1386)
);

XNOR2xp5_ASAP7_75t_L g1387 ( 
.A(n_1350),
.B(n_1292),
.Y(n_1387)
);

INVxp67_ASAP7_75t_L g1388 ( 
.A(n_1341),
.Y(n_1388)
);

INVxp67_ASAP7_75t_L g1389 ( 
.A(n_1351),
.Y(n_1389)
);

NAND2xp33_ASAP7_75t_R g1390 ( 
.A(n_1373),
.B(n_1288),
.Y(n_1390)
);

XNOR2xp5_ASAP7_75t_L g1391 ( 
.A(n_1350),
.B(n_1277),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1365),
.B(n_1371),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1355),
.B(n_1287),
.Y(n_1393)
);

NAND2xp33_ASAP7_75t_R g1394 ( 
.A(n_1373),
.B(n_1298),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_1344),
.Y(n_1395)
);

NAND2xp33_ASAP7_75t_R g1396 ( 
.A(n_1375),
.B(n_1331),
.Y(n_1396)
);

NAND2xp33_ASAP7_75t_R g1397 ( 
.A(n_1375),
.B(n_1278),
.Y(n_1397)
);

INVxp67_ASAP7_75t_L g1398 ( 
.A(n_1356),
.Y(n_1398)
);

NAND2xp33_ASAP7_75t_R g1399 ( 
.A(n_1365),
.B(n_1336),
.Y(n_1399)
);

NAND2xp33_ASAP7_75t_R g1400 ( 
.A(n_1365),
.B(n_1336),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1355),
.B(n_1287),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_R g1402 ( 
.A(n_1368),
.B(n_1329),
.Y(n_1402)
);

INVxp67_ASAP7_75t_L g1403 ( 
.A(n_1356),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1358),
.B(n_1295),
.Y(n_1404)
);

XNOR2xp5_ASAP7_75t_L g1405 ( 
.A(n_1354),
.B(n_1283),
.Y(n_1405)
);

NAND2xp33_ASAP7_75t_R g1406 ( 
.A(n_1365),
.B(n_1328),
.Y(n_1406)
);

INVxp67_ASAP7_75t_L g1407 ( 
.A(n_1366),
.Y(n_1407)
);

NAND2xp33_ASAP7_75t_R g1408 ( 
.A(n_1365),
.B(n_1328),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1366),
.Y(n_1409)
);

NAND2xp33_ASAP7_75t_R g1410 ( 
.A(n_1346),
.B(n_1329),
.Y(n_1410)
);

INVxp67_ASAP7_75t_L g1411 ( 
.A(n_1369),
.Y(n_1411)
);

NAND2xp33_ASAP7_75t_SL g1412 ( 
.A(n_1349),
.B(n_1314),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1358),
.B(n_1302),
.Y(n_1413)
);

XNOR2xp5_ASAP7_75t_L g1414 ( 
.A(n_1354),
.B(n_1333),
.Y(n_1414)
);

NOR2xp67_ASAP7_75t_L g1415 ( 
.A(n_1388),
.B(n_1370),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1380),
.B(n_1360),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1386),
.B(n_1360),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1385),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1413),
.Y(n_1419)
);

AND2x4_ASAP7_75t_SL g1420 ( 
.A(n_1379),
.B(n_1374),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1413),
.B(n_1345),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1393),
.B(n_1345),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1393),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1401),
.B(n_1348),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1392),
.B(n_1372),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1392),
.B(n_1372),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1401),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1404),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1384),
.B(n_1340),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1381),
.B(n_1340),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1379),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1409),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1411),
.B(n_1340),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1377),
.B(n_1347),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1412),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1419),
.B(n_1352),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1434),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1429),
.B(n_1383),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1416),
.Y(n_1439)
);

NAND3xp33_ASAP7_75t_L g1440 ( 
.A(n_1419),
.B(n_1405),
.C(n_1391),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1429),
.B(n_1370),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1416),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1429),
.B(n_1430),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1416),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1428),
.B(n_1352),
.Y(n_1445)
);

OAI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1432),
.A2(n_1396),
.B1(n_1410),
.B2(n_1368),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1432),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1430),
.B(n_1359),
.Y(n_1448)
);

AOI31xp33_ASAP7_75t_L g1449 ( 
.A1(n_1435),
.A2(n_1397),
.A3(n_1390),
.B(n_1414),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1417),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1431),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1417),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1417),
.Y(n_1453)
);

AOI221xp5_ASAP7_75t_SL g1454 ( 
.A1(n_1435),
.A2(n_1387),
.B1(n_1382),
.B2(n_1364),
.C(n_1361),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1428),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1430),
.B(n_1357),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1438),
.B(n_1423),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1443),
.B(n_1425),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1450),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1455),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1455),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1450),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1449),
.B(n_1418),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1443),
.B(n_1425),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1452),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1447),
.Y(n_1466)
);

OAI21xp33_ASAP7_75t_L g1467 ( 
.A1(n_1440),
.A2(n_1378),
.B(n_1418),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1456),
.B(n_1423),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1452),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1439),
.B(n_1425),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1439),
.B(n_1426),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1442),
.B(n_1426),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1442),
.B(n_1426),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1441),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1447),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1441),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1448),
.B(n_1423),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1453),
.B(n_1433),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1478),
.B(n_1454),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_L g1480 ( 
.A(n_1467),
.B(n_1440),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1478),
.B(n_1454),
.Y(n_1481)
);

INVxp33_ASAP7_75t_L g1482 ( 
.A(n_1463),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1476),
.B(n_1433),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1460),
.Y(n_1484)
);

AO221x2_ASAP7_75t_L g1485 ( 
.A1(n_1467),
.A2(n_1446),
.B1(n_1394),
.B2(n_1453),
.C(n_1444),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1476),
.B(n_1433),
.Y(n_1486)
);

INVx2_ASAP7_75t_SL g1487 ( 
.A(n_1475),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1474),
.B(n_1427),
.Y(n_1488)
);

OAI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1466),
.A2(n_1438),
.B1(n_1451),
.B2(n_1408),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1482),
.B(n_1475),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1487),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1484),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1485),
.B(n_1458),
.Y(n_1493)
);

INVxp67_ASAP7_75t_L g1494 ( 
.A(n_1480),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1488),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1483),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1486),
.Y(n_1497)
);

INVx1_ASAP7_75t_SL g1498 ( 
.A(n_1479),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1485),
.B(n_1458),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1481),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_SL g1501 ( 
.A(n_1489),
.B(n_1466),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1487),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1496),
.B(n_1477),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1498),
.A2(n_1474),
.B1(n_1457),
.B2(n_1468),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1494),
.B(n_1464),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1491),
.Y(n_1506)
);

INVxp67_ASAP7_75t_SL g1507 ( 
.A(n_1490),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1500),
.B(n_1464),
.Y(n_1508)
);

OAI321xp33_ASAP7_75t_L g1509 ( 
.A1(n_1501),
.A2(n_1451),
.A3(n_1421),
.B1(n_1477),
.B2(n_1424),
.C(n_1422),
.Y(n_1509)
);

AOI21xp33_ASAP7_75t_L g1510 ( 
.A1(n_1500),
.A2(n_1395),
.B(n_1421),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1502),
.A2(n_1474),
.B1(n_1457),
.B2(n_1448),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1506),
.B(n_1495),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1503),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1507),
.B(n_1496),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1505),
.B(n_1495),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1508),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1511),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1510),
.B(n_1493),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1504),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1509),
.B(n_1492),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1514),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1512),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1514),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1513),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1517),
.B(n_1493),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1512),
.Y(n_1526)
);

BUFx12f_ASAP7_75t_L g1527 ( 
.A(n_1518),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1519),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1515),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1516),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1520),
.B(n_1499),
.Y(n_1531)
);

NOR3xp33_ASAP7_75t_L g1532 ( 
.A(n_1528),
.B(n_1520),
.C(n_1499),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1526),
.A2(n_1531),
.B(n_1528),
.Y(n_1533)
);

NOR3xp33_ASAP7_75t_L g1534 ( 
.A(n_1523),
.B(n_1492),
.C(n_1289),
.Y(n_1534)
);

NAND4xp75_ASAP7_75t_L g1535 ( 
.A(n_1521),
.B(n_1497),
.C(n_1415),
.D(n_1300),
.Y(n_1535)
);

NAND4xp25_ASAP7_75t_SL g1536 ( 
.A(n_1525),
.B(n_1497),
.C(n_1364),
.D(n_1470),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1525),
.B(n_1460),
.Y(n_1537)
);

AOI211xp5_ASAP7_75t_L g1538 ( 
.A1(n_1524),
.A2(n_1402),
.B(n_1326),
.C(n_1308),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1522),
.B(n_1461),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1527),
.B(n_1461),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1533),
.Y(n_1541)
);

NAND3xp33_ASAP7_75t_SL g1542 ( 
.A(n_1532),
.B(n_1521),
.C(n_1522),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1540),
.Y(n_1543)
);

O2A1O1Ixp33_ASAP7_75t_L g1544 ( 
.A1(n_1534),
.A2(n_1530),
.B(n_1529),
.C(n_1527),
.Y(n_1544)
);

NOR3x1_ASAP7_75t_L g1545 ( 
.A(n_1535),
.B(n_1346),
.C(n_1363),
.Y(n_1545)
);

OAI211xp5_ASAP7_75t_L g1546 ( 
.A1(n_1537),
.A2(n_1290),
.B(n_1302),
.C(n_1309),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1539),
.Y(n_1547)
);

XOR2x2_ASAP7_75t_L g1548 ( 
.A(n_1542),
.B(n_1538),
.Y(n_1548)
);

NOR2xp67_ASAP7_75t_L g1549 ( 
.A(n_1543),
.B(n_1536),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1541),
.B(n_1470),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1547),
.B(n_1459),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1544),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1546),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1545),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_SL g1555 ( 
.A(n_1553),
.B(n_1459),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_R g1556 ( 
.A(n_1552),
.B(n_1316),
.Y(n_1556)
);

NAND2x1_ASAP7_75t_SL g1557 ( 
.A(n_1554),
.B(n_1459),
.Y(n_1557)
);

NAND3xp33_ASAP7_75t_L g1558 ( 
.A(n_1549),
.B(n_1309),
.C(n_1465),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_R g1559 ( 
.A(n_1550),
.B(n_1399),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_R g1560 ( 
.A(n_1548),
.B(n_1400),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_R g1561 ( 
.A(n_1551),
.B(n_1406),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1558),
.A2(n_1549),
.B1(n_1551),
.B2(n_1469),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1557),
.Y(n_1563)
);

AO22x2_ASAP7_75t_L g1564 ( 
.A1(n_1555),
.A2(n_1556),
.B1(n_1560),
.B2(n_1559),
.Y(n_1564)
);

INVx3_ASAP7_75t_L g1565 ( 
.A(n_1561),
.Y(n_1565)
);

OAI22xp33_ASAP7_75t_SL g1566 ( 
.A1(n_1555),
.A2(n_1469),
.B1(n_1465),
.B2(n_1462),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1557),
.Y(n_1567)
);

AOI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1558),
.A2(n_1473),
.B1(n_1472),
.B2(n_1471),
.Y(n_1568)
);

INVxp67_ASAP7_75t_L g1569 ( 
.A(n_1555),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1569),
.A2(n_1462),
.B1(n_1407),
.B2(n_1403),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1564),
.B(n_1471),
.Y(n_1571)
);

AND4x2_ASAP7_75t_L g1572 ( 
.A(n_1565),
.B(n_1376),
.C(n_1420),
.D(n_1415),
.Y(n_1572)
);

OAI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1563),
.A2(n_1437),
.B(n_1473),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1567),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1562),
.Y(n_1575)
);

XNOR2x1_ASAP7_75t_L g1576 ( 
.A(n_1574),
.B(n_1571),
.Y(n_1576)
);

CKINVDCx16_ASAP7_75t_R g1577 ( 
.A(n_1575),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_1570),
.Y(n_1578)
);

OAI321xp33_ASAP7_75t_L g1579 ( 
.A1(n_1570),
.A2(n_1568),
.A3(n_1566),
.B1(n_1398),
.B2(n_1389),
.C(n_1472),
.Y(n_1579)
);

AOI31xp33_ASAP7_75t_L g1580 ( 
.A1(n_1576),
.A2(n_1577),
.A3(n_1578),
.B(n_1579),
.Y(n_1580)
);

AOI31xp33_ASAP7_75t_L g1581 ( 
.A1(n_1576),
.A2(n_1572),
.A3(n_1573),
.B(n_1445),
.Y(n_1581)
);

XOR2xp5_ASAP7_75t_L g1582 ( 
.A(n_1580),
.B(n_1377),
.Y(n_1582)
);

OAI322xp33_ASAP7_75t_L g1583 ( 
.A1(n_1581),
.A2(n_1361),
.A3(n_1437),
.B1(n_1444),
.B2(n_1427),
.C1(n_1310),
.C2(n_1436),
.Y(n_1583)
);

AOI32xp33_ASAP7_75t_L g1584 ( 
.A1(n_1582),
.A2(n_1420),
.A3(n_1437),
.B1(n_1362),
.B2(n_1431),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_SL g1585 ( 
.A1(n_1583),
.A2(n_1437),
.B1(n_1431),
.B2(n_1420),
.Y(n_1585)
);

BUFx2_ASAP7_75t_SL g1586 ( 
.A(n_1585),
.Y(n_1586)
);

AOI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1586),
.A2(n_1584),
.B1(n_1377),
.B2(n_1431),
.C(n_1427),
.Y(n_1587)
);

AOI211xp5_ASAP7_75t_L g1588 ( 
.A1(n_1587),
.A2(n_1284),
.B(n_1357),
.C(n_1371),
.Y(n_1588)
);


endmodule