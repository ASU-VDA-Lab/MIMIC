module fake_aes_2099_n_19 (n_1, n_2, n_0, n_19);
input n_1;
input n_2;
input n_0;
output n_19;
wire n_5;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_3;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_6;
wire n_4;
wire n_7;
NAND2xp5_ASAP7_75t_L g3 ( .A(n_1), .B(n_2), .Y(n_3) );
INVx2_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
NAND2xp33_ASAP7_75t_R g5 ( .A(n_0), .B(n_1), .Y(n_5) );
AO31x2_ASAP7_75t_L g6 ( .A1(n_4), .A2(n_0), .A3(n_1), .B(n_2), .Y(n_6) );
AND2x2_ASAP7_75t_L g7 ( .A(n_3), .B(n_0), .Y(n_7) );
NAND2x1p5_ASAP7_75t_L g8 ( .A(n_5), .B(n_0), .Y(n_8) );
OR2x2_ASAP7_75t_L g9 ( .A(n_8), .B(n_1), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_7), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
AOI22xp5_ASAP7_75t_L g12 ( .A1(n_10), .A2(n_8), .B1(n_5), .B2(n_7), .Y(n_12) );
OAI21xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_9), .B(n_6), .Y(n_13) );
AOI211x1_ASAP7_75t_SL g14 ( .A1(n_11), .A2(n_6), .B(n_1), .C(n_2), .Y(n_14) );
OAI211xp5_ASAP7_75t_SL g15 ( .A1(n_14), .A2(n_6), .B(n_0), .C(n_2), .Y(n_15) );
HB1xp67_ASAP7_75t_L g16 ( .A(n_13), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
AOI21xp5_ASAP7_75t_L g18 ( .A1(n_15), .A2(n_14), .B(n_6), .Y(n_18) );
OAI21xp5_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_0), .B(n_17), .Y(n_19) );
endmodule