module fake_jpeg_2390_n_118 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_118);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_43),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_26),
.B(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_48),
.A2(n_30),
.B1(n_37),
.B2(n_39),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_37),
.B1(n_39),
.B2(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_29),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_57),
.Y(n_59)
);

NAND3xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_68),
.C(n_38),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_49),
.B1(n_56),
.B2(n_31),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_67),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_64),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_44),
.B1(n_46),
.B2(n_27),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_42),
.B1(n_4),
.B2(n_7),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_38),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_68),
.B(n_36),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_71),
.B(n_73),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_74),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_32),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_78),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_42),
.B1(n_32),
.B2(n_31),
.Y(n_77)
);

AO22x1_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_2),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_80),
.A2(n_16),
.B1(n_25),
.B2(n_24),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_3),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_3),
.Y(n_86)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_83),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_80),
.A2(n_72),
.B1(n_69),
.B2(n_70),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_86),
.Y(n_103)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_7),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_94),
.Y(n_96)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_12),
.B(n_20),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_92),
.B(n_9),
.Y(n_99)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_14),
.C(n_19),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_93),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_95),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_104),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_103),
.A2(n_93),
.B1(n_92),
.B2(n_87),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_101),
.C(n_97),
.Y(n_109)
);

OA21x2_ASAP7_75t_SL g112 ( 
.A1(n_109),
.A2(n_108),
.B(n_100),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_110),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_112),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_114),
.B(n_98),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_102),
.C(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_96),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_99),
.Y(n_118)
);


endmodule