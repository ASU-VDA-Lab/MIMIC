module fake_jpeg_28149_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx13_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

INVx11_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx12_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_18),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_8),
.Y(n_21)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_15),
.B(n_0),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_15),
.Y(n_24)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_8),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_22),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_25),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_21),
.A2(n_17),
.B(n_13),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_19),
.B(n_13),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_17),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_11),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_8),
.B1(n_10),
.B2(n_20),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_22),
.A2(n_15),
.B1(n_9),
.B2(n_13),
.Y(n_30)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_36),
.Y(n_44)
);

AND2x6_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_2),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_27),
.C(n_20),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_42),
.B(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_36),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_41),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_44),
.C(n_43),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_37),
.B1(n_18),
.B2(n_10),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_46),
.A2(n_47),
.B(n_48),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_42),
.B(n_12),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_51),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_12),
.B(n_14),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_55),
.B(n_12),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_10),
.B1(n_18),
.B2(n_6),
.Y(n_55)
);

AOI322xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_12),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_1),
.C2(n_14),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_12),
.C(n_14),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_58),
.B(n_5),
.Y(n_59)
);


endmodule