module fake_jpeg_16234_n_130 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_130);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx6_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_23),
.B1(n_18),
.B2(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_27),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_26),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_22),
.B1(n_24),
.B2(n_30),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_23),
.Y(n_68)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_58),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_32),
.A2(n_16),
.B1(n_29),
.B2(n_26),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_6),
.B(n_7),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_20),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_22),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_61),
.Y(n_73)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_67),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_33),
.B1(n_32),
.B2(n_47),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_70),
.B1(n_77),
.B2(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_66),
.B(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_21),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_81),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_30),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_11),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_40),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_74),
.B(n_76),
.Y(n_96)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_46),
.Y(n_91)
);

FAx1_ASAP7_75t_SL g76 ( 
.A(n_54),
.B(n_2),
.CI(n_6),
.CON(n_76),
.SN(n_76)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_7),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_84),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_79),
.B1(n_55),
.B2(n_59),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_91),
.Y(n_97)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_51),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_95),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_73),
.Y(n_95)
);

OA21x2_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_70),
.B(n_76),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_101),
.A2(n_96),
.B(n_90),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_79),
.B1(n_87),
.B2(n_88),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_96),
.B(n_90),
.C(n_93),
.D(n_89),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_105),
.B(n_107),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_102),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_108),
.B(n_109),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_100),
.A2(n_82),
.B(n_94),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_111),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_92),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_112),
.A2(n_103),
.B(n_99),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_110),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_117),
.A2(n_84),
.B1(n_78),
.B2(n_75),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_120),
.A2(n_84),
.B1(n_78),
.B2(n_75),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_118),
.B1(n_116),
.B2(n_115),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_124),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_121),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_126),
.B(n_49),
.Y(n_129)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_129),
.Y(n_130)
);


endmodule