module fake_ariane_1999_n_1845 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1845);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1845;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_4),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_63),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_19),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_23),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_35),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_42),
.Y(n_184)
);

BUFx8_ASAP7_75t_SL g185 ( 
.A(n_151),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_75),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_131),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_87),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_141),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_56),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_13),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_77),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_110),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_94),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_20),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_49),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_150),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_178),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_73),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_64),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_114),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_134),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_101),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_4),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_43),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_2),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_71),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_44),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_129),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_78),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_119),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_124),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_102),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_127),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_25),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_37),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_36),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_49),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_108),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_1),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_70),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_45),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_72),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_132),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_12),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_154),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_41),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_121),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_167),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_45),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_172),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_85),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_166),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_158),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_10),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_54),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_157),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_81),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_133),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_26),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_34),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_8),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_115),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_174),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_169),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_60),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_107),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_40),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_46),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_137),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_74),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_68),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_32),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_33),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_95),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_0),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_17),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_8),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_80),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_11),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_159),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_62),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_24),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_109),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_9),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_37),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_116),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_29),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_20),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_51),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_93),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_143),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_99),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_147),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_136),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_50),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_18),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_34),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_22),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_0),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_6),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_13),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_2),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_50),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_46),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_100),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_3),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_18),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_36),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_130),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_31),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_128),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_6),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_33),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_32),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_113),
.Y(n_297)
);

BUFx10_ASAP7_75t_L g298 ( 
.A(n_126),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_105),
.Y(n_299)
);

BUFx10_ASAP7_75t_L g300 ( 
.A(n_162),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_12),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_23),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_148),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_79),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_170),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_51),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_57),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_16),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_24),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_161),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_144),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_29),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_146),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_48),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_27),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_67),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_7),
.Y(n_317)
);

BUFx2_ASAP7_75t_SL g318 ( 
.A(n_152),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_19),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_25),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_160),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_47),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_145),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_90),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_96),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_7),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_176),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_153),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_177),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_139),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_112),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_14),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_149),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_15),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_163),
.Y(n_335)
);

INVxp33_ASAP7_75t_L g336 ( 
.A(n_65),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_140),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_91),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_117),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_44),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_22),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_98),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_47),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_156),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_16),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_142),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_42),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_39),
.Y(n_348)
);

BUFx5_ASAP7_75t_L g349 ( 
.A(n_41),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_55),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_92),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_164),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_58),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_120),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_52),
.Y(n_355)
);

BUFx10_ASAP7_75t_L g356 ( 
.A(n_27),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_185),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_349),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_352),
.B(n_1),
.Y(n_359)
);

INVxp33_ASAP7_75t_SL g360 ( 
.A(n_319),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_279),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_182),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_349),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_349),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_182),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_267),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_288),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_264),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_270),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_189),
.B(n_3),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_349),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_314),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_201),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_225),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_349),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_238),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_260),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_349),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_349),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_299),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_349),
.B(n_5),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_339),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_255),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_219),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_294),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_255),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_197),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_179),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_255),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_179),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_221),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_255),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_295),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_220),
.B(n_5),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_199),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_255),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_223),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_180),
.B(n_9),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_353),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_353),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_337),
.Y(n_401)
);

BUFx2_ASAP7_75t_SL g402 ( 
.A(n_233),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_181),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_353),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_228),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_210),
.B(n_10),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_226),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_233),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_239),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_353),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_233),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_298),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_231),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_353),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_184),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_236),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_294),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_294),
.Y(n_418)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_197),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_237),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_184),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_315),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_298),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_315),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_336),
.B(n_11),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_298),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_181),
.Y(n_427)
);

NOR2xp67_ASAP7_75t_L g428 ( 
.A(n_340),
.B(n_14),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_320),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_320),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_242),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_249),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_300),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_183),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_250),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_211),
.B(n_15),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_350),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_350),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_254),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_300),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_300),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_257),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_201),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_188),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_188),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_247),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_405),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_360),
.A2(n_368),
.B1(n_401),
.B2(n_395),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_358),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_358),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_409),
.Y(n_451)
);

INVx5_ASAP7_75t_L g452 ( 
.A(n_409),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_363),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_363),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_409),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_364),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_441),
.B(n_186),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_409),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_364),
.B(n_213),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_371),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_371),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_409),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_375),
.B(n_215),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_409),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_375),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_378),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_378),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_379),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_379),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_383),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_383),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_441),
.B(n_194),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_386),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_386),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_389),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_389),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_392),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_392),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_396),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_441),
.B(n_194),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_396),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_399),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_399),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_441),
.B(n_229),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_444),
.B(n_232),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_400),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_400),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_404),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_404),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_444),
.B(n_234),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_410),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_410),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_361),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_369),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_414),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_373),
.B(n_252),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_414),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_373),
.B(n_252),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_445),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_445),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_362),
.B(n_212),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_381),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_446),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_446),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_415),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_415),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_365),
.B(n_212),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_421),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_387),
.B(n_240),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_393),
.B(n_183),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_421),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_422),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_422),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_398),
.A2(n_327),
.B(n_247),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_424),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_424),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_429),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_429),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_430),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_430),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_419),
.B(n_240),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_437),
.B(n_276),
.Y(n_522)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_384),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_437),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_469),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_472),
.B(n_402),
.Y(n_526)
);

NAND3xp33_ASAP7_75t_L g527 ( 
.A(n_449),
.B(n_436),
.C(n_406),
.Y(n_527)
);

NAND2xp33_ASAP7_75t_SL g528 ( 
.A(n_523),
.B(n_357),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_469),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_469),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_467),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_522),
.A2(n_359),
.B1(n_370),
.B2(n_394),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_467),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_457),
.B(n_402),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_467),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_467),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_507),
.B(n_388),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_467),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_470),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_470),
.Y(n_540)
);

BUFx10_ASAP7_75t_L g541 ( 
.A(n_501),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_523),
.B(n_391),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_447),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_447),
.B(n_390),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_449),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_471),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_522),
.A2(n_425),
.B1(n_427),
.B2(n_403),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_471),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_522),
.A2(n_434),
.B1(n_428),
.B2(n_443),
.Y(n_549)
);

BUFx10_ASAP7_75t_L g550 ( 
.A(n_501),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_523),
.B(n_397),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_507),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_522),
.A2(n_428),
.B1(n_309),
.B2(n_345),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_493),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_467),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_467),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_L g557 ( 
.A(n_502),
.B(n_407),
.Y(n_557)
);

AND2x6_ASAP7_75t_L g558 ( 
.A(n_502),
.B(n_327),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_501),
.B(n_385),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_472),
.B(n_413),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_473),
.Y(n_561)
);

OAI22xp33_ASAP7_75t_L g562 ( 
.A1(n_523),
.A2(n_417),
.B1(n_418),
.B2(n_243),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_473),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_522),
.A2(n_241),
.B1(n_347),
.B2(n_259),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_474),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_474),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_472),
.B(n_416),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_475),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_450),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_501),
.B(n_438),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_475),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_476),
.Y(n_572)
);

NAND2xp33_ASAP7_75t_L g573 ( 
.A(n_502),
.B(n_420),
.Y(n_573)
);

OAI22xp33_ASAP7_75t_L g574 ( 
.A1(n_523),
.A2(n_290),
.B1(n_334),
.B2(n_367),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_450),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_510),
.B(n_380),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_476),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_507),
.B(n_438),
.Y(n_578)
);

BUFx6f_ASAP7_75t_SL g579 ( 
.A(n_501),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_450),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_450),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_450),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_479),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_461),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_472),
.A2(n_207),
.B1(n_284),
.B2(n_209),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_509),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_479),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_461),
.Y(n_588)
);

INVxp33_ASAP7_75t_L g589 ( 
.A(n_510),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_461),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_509),
.B(n_521),
.Y(n_591)
);

OAI22xp33_ASAP7_75t_L g592 ( 
.A1(n_448),
.A2(n_372),
.B1(n_439),
.B2(n_435),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_472),
.B(n_431),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_461),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_481),
.Y(n_595)
);

OR2x6_ASAP7_75t_L g596 ( 
.A(n_480),
.B(n_318),
.Y(n_596)
);

AND2x6_ASAP7_75t_L g597 ( 
.A(n_502),
.B(n_346),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_480),
.B(n_432),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_480),
.B(n_442),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_481),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_480),
.B(n_187),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_461),
.Y(n_602)
);

NOR2x1p5_ASAP7_75t_L g603 ( 
.A(n_512),
.B(n_374),
.Y(n_603)
);

AND2x6_ASAP7_75t_L g604 ( 
.A(n_502),
.B(n_346),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_480),
.B(n_265),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_509),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_478),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_521),
.Y(n_608)
);

BUFx4f_ASAP7_75t_L g609 ( 
.A(n_502),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_496),
.B(n_498),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_499),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_478),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_477),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_483),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_521),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_499),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_483),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_496),
.B(n_328),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_484),
.B(n_366),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_486),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_496),
.A2(n_269),
.B1(n_277),
.B2(n_278),
.Y(n_621)
);

AND3x1_ASAP7_75t_L g622 ( 
.A(n_448),
.B(n_192),
.C(n_191),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_484),
.B(n_408),
.Y(n_623)
);

INVx5_ASAP7_75t_L g624 ( 
.A(n_455),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_496),
.A2(n_317),
.B1(n_283),
.B2(n_280),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_477),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_486),
.Y(n_627)
);

AND2x2_ASAP7_75t_SL g628 ( 
.A(n_502),
.B(n_239),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_493),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_496),
.B(n_498),
.Y(n_630)
);

AND2x6_ASAP7_75t_L g631 ( 
.A(n_498),
.B(n_499),
.Y(n_631)
);

NAND2xp33_ASAP7_75t_L g632 ( 
.A(n_453),
.B(n_186),
.Y(n_632)
);

INVxp67_ASAP7_75t_SL g633 ( 
.A(n_459),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_499),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_487),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_498),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_499),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_477),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_498),
.B(n_376),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_453),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_506),
.A2(n_440),
.B1(n_433),
.B2(n_426),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_459),
.B(n_377),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_500),
.Y(n_643)
);

AND2x6_ASAP7_75t_L g644 ( 
.A(n_500),
.B(n_276),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_454),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_500),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_454),
.B(n_411),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_456),
.Y(n_648)
);

NAND2xp33_ASAP7_75t_R g649 ( 
.A(n_514),
.B(n_412),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_494),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_456),
.B(n_190),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_460),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_494),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_463),
.B(n_190),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_460),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_500),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_465),
.B(n_195),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_487),
.Y(n_658)
);

BUFx10_ASAP7_75t_L g659 ( 
.A(n_465),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_466),
.B(n_423),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_489),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_463),
.B(n_195),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_512),
.B(n_312),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_500),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_466),
.Y(n_665)
);

NAND2x1p5_ASAP7_75t_L g666 ( 
.A(n_514),
.B(n_245),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_512),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_468),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_468),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_485),
.B(n_198),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_485),
.B(n_198),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_514),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_512),
.B(n_312),
.Y(n_673)
);

OR2x6_ASAP7_75t_L g674 ( 
.A(n_490),
.B(n_193),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_503),
.B(n_200),
.Y(n_675)
);

INVx4_ASAP7_75t_SL g676 ( 
.A(n_455),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_503),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_633),
.B(n_512),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_550),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_659),
.B(n_200),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_659),
.B(n_550),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_623),
.B(n_518),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_545),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_545),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_640),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_663),
.B(n_518),
.Y(n_686)
);

NAND3xp33_ASAP7_75t_L g687 ( 
.A(n_619),
.B(n_205),
.C(n_196),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_550),
.Y(n_688)
);

NOR3xp33_ASAP7_75t_L g689 ( 
.A(n_629),
.B(n_306),
.C(n_205),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_663),
.B(n_518),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_550),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_640),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_659),
.B(n_202),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_645),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_552),
.B(n_518),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_673),
.B(n_518),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_541),
.B(n_609),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_667),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_554),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_667),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_544),
.Y(n_701)
);

INVxp33_ASAP7_75t_L g702 ( 
.A(n_544),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_629),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_541),
.B(n_202),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_673),
.B(n_504),
.Y(n_705)
);

INVx4_ASAP7_75t_L g706 ( 
.A(n_579),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_645),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_543),
.B(n_382),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_591),
.B(n_504),
.Y(n_709)
);

NOR2xp67_ASAP7_75t_L g710 ( 
.A(n_647),
.B(n_490),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_591),
.B(n_506),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_537),
.B(n_508),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_525),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_525),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_552),
.B(n_508),
.Y(n_715)
);

OAI21xp5_ASAP7_75t_L g716 ( 
.A1(n_569),
.A2(n_492),
.B(n_489),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_586),
.B(n_511),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_586),
.B(n_511),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_529),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_537),
.B(n_513),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_606),
.B(n_513),
.Y(n_721)
);

BUFx6f_ASAP7_75t_SL g722 ( 
.A(n_559),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_606),
.B(n_519),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_650),
.B(n_519),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_650),
.B(n_524),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_539),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_608),
.B(n_524),
.Y(n_727)
);

AO22x2_ASAP7_75t_L g728 ( 
.A1(n_576),
.A2(n_520),
.B1(n_517),
.B2(n_516),
.Y(n_728)
);

AOI221xp5_ASAP7_75t_L g729 ( 
.A1(n_562),
.A2(n_322),
.B1(n_196),
.B2(n_206),
.C(n_216),
.Y(n_729)
);

NOR3xp33_ASAP7_75t_L g730 ( 
.A(n_554),
.B(n_216),
.C(n_206),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_576),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_540),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_608),
.A2(n_321),
.B1(n_354),
.B2(n_351),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_615),
.B(n_505),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_540),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_541),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_615),
.B(n_258),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_674),
.A2(n_321),
.B1(n_354),
.B2(n_351),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_674),
.A2(n_325),
.B1(n_214),
.B2(n_208),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_546),
.Y(n_740)
);

INVxp67_ASAP7_75t_SL g741 ( 
.A(n_609),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_648),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_631),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_542),
.B(n_505),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_631),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_656),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_551),
.B(n_505),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_528),
.Y(n_748)
);

INVx8_ASAP7_75t_L g749 ( 
.A(n_579),
.Y(n_749)
);

AND2x4_ASAP7_75t_SL g750 ( 
.A(n_559),
.B(n_312),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_652),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_674),
.A2(n_262),
.B1(n_344),
.B2(n_203),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_630),
.B(n_515),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_677),
.B(n_515),
.Y(n_754)
);

NOR2x1_ASAP7_75t_L g755 ( 
.A(n_660),
.B(n_515),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_548),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_628),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_653),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_653),
.B(n_356),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_656),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_677),
.B(n_578),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_578),
.A2(n_520),
.B(n_517),
.C(n_516),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_570),
.B(n_516),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_548),
.Y(n_764)
);

OAI22xp33_ASAP7_75t_L g765 ( 
.A1(n_674),
.A2(n_217),
.B1(n_218),
.B2(n_266),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_609),
.B(n_203),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_561),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_559),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_674),
.A2(n_262),
.B1(n_344),
.B2(n_204),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_559),
.B(n_517),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_641),
.B(n_217),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_592),
.B(n_218),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_656),
.B(n_204),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_570),
.B(n_520),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_549),
.B(n_356),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_642),
.B(n_560),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_561),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_588),
.B(n_208),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_570),
.B(n_526),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_588),
.B(n_214),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_570),
.B(n_356),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_596),
.A2(n_266),
.B1(n_355),
.B2(n_348),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_563),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_611),
.B(n_492),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_611),
.B(n_497),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_611),
.B(n_497),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_616),
.B(n_634),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_563),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_588),
.B(n_311),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_603),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_590),
.B(n_311),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_567),
.B(n_261),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_649),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_590),
.B(n_316),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_616),
.B(n_316),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_565),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_596),
.B(n_251),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_590),
.B(n_324),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_603),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_636),
.B(n_324),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_529),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_616),
.B(n_325),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_547),
.B(n_322),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_634),
.B(n_329),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_655),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_565),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_636),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_610),
.A2(n_326),
.B(n_332),
.C(n_341),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_598),
.B(n_271),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_636),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_628),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_636),
.B(n_628),
.Y(n_812)
);

BUFx6f_ASAP7_75t_SL g813 ( 
.A(n_596),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_634),
.B(n_329),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_637),
.B(n_333),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_637),
.B(n_333),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_569),
.B(n_335),
.Y(n_817)
);

NAND2x1p5_ASAP7_75t_L g818 ( 
.A(n_637),
.B(n_256),
.Y(n_818)
);

INVx8_ASAP7_75t_L g819 ( 
.A(n_579),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_566),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_566),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_531),
.A2(n_451),
.B(n_458),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_596),
.B(n_326),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_593),
.B(n_281),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_643),
.B(n_335),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_643),
.B(n_338),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_568),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_596),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_643),
.B(n_338),
.Y(n_829)
);

OAI22xp33_ASAP7_75t_L g830 ( 
.A1(n_601),
.A2(n_343),
.B1(n_332),
.B2(n_341),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_599),
.B(n_343),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_646),
.B(n_282),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_622),
.B(n_348),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_534),
.B(n_285),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_639),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_646),
.B(n_286),
.Y(n_836)
);

NAND2xp33_ASAP7_75t_L g837 ( 
.A(n_631),
.B(n_289),
.Y(n_837)
);

INVx8_ASAP7_75t_L g838 ( 
.A(n_631),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_665),
.Y(n_839)
);

O2A1O1Ixp5_ASAP7_75t_L g840 ( 
.A1(n_654),
.A2(n_313),
.B(n_268),
.C(n_275),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_631),
.A2(n_495),
.B1(n_491),
.B2(n_488),
.Y(n_841)
);

NAND2x1_ASAP7_75t_L g842 ( 
.A(n_631),
.B(n_451),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_568),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_665),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_607),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_803),
.A2(n_631),
.B1(n_585),
.B2(n_644),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_726),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_713),
.Y(n_848)
);

OAI321xp33_ASAP7_75t_L g849 ( 
.A1(n_765),
.A2(n_574),
.A3(n_532),
.B1(n_527),
.B2(n_621),
.C(n_625),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_743),
.A2(n_646),
.B1(n_664),
.B2(n_527),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_702),
.B(n_622),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_762),
.A2(n_672),
.B(n_580),
.Y(n_852)
);

INVxp67_ASAP7_75t_L g853 ( 
.A(n_701),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_682),
.B(n_605),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_776),
.B(n_662),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_SL g856 ( 
.A(n_699),
.B(n_589),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_682),
.B(n_618),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_838),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_710),
.B(n_664),
.Y(n_859)
);

AO21x1_ASAP7_75t_L g860 ( 
.A1(n_834),
.A2(n_666),
.B(n_573),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_776),
.B(n_670),
.Y(n_861)
);

NOR3xp33_ASAP7_75t_L g862 ( 
.A(n_765),
.B(n_687),
.C(n_703),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_761),
.B(n_664),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_715),
.B(n_564),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_834),
.A2(n_575),
.B(n_594),
.C(n_602),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_830),
.A2(n_557),
.B(n_632),
.C(n_657),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_775),
.A2(n_644),
.B1(n_668),
.B2(n_669),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_702),
.B(n_553),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_715),
.B(n_675),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_744),
.A2(n_672),
.B(n_580),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_743),
.A2(n_668),
.B1(n_669),
.B2(n_651),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_717),
.B(n_671),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_745),
.A2(n_575),
.B1(n_581),
.B2(n_582),
.Y(n_873)
);

OAI321xp33_ASAP7_75t_L g874 ( 
.A1(n_729),
.A2(n_666),
.A3(n_572),
.B1(n_661),
.B2(n_658),
.C(n_577),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_830),
.A2(n_594),
.B(n_582),
.C(n_584),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_698),
.B(n_700),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_713),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_747),
.A2(n_602),
.B(n_584),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_787),
.A2(n_678),
.B(n_686),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_690),
.A2(n_581),
.B(n_533),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_696),
.A2(n_531),
.B(n_533),
.Y(n_881)
);

INVx11_ASAP7_75t_L g882 ( 
.A(n_758),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_717),
.B(n_644),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_721),
.B(n_644),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_838),
.Y(n_885)
);

O2A1O1Ixp5_ASAP7_75t_L g886 ( 
.A1(n_766),
.A2(n_600),
.B(n_577),
.C(n_661),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_753),
.A2(n_556),
.B(n_538),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_773),
.A2(n_556),
.B(n_538),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_745),
.A2(n_572),
.B1(n_595),
.B2(n_658),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_768),
.B(n_688),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_695),
.A2(n_620),
.B(n_600),
.C(n_587),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_R g892 ( 
.A(n_731),
.B(n_838),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_724),
.B(n_355),
.Y(n_893)
);

NOR2x1p5_ASAP7_75t_L g894 ( 
.A(n_772),
.B(n_823),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_688),
.B(n_607),
.Y(n_895)
);

O2A1O1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_808),
.A2(n_620),
.B(n_627),
.C(n_635),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_725),
.B(n_571),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_773),
.A2(n_535),
.B(n_536),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_792),
.B(n_555),
.Y(n_899)
);

O2A1O1Ixp5_ASAP7_75t_L g900 ( 
.A1(n_766),
.A2(n_583),
.B(n_587),
.C(n_595),
.Y(n_900)
);

OAI21xp33_ASAP7_75t_L g901 ( 
.A1(n_792),
.A2(n_302),
.B(n_296),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_705),
.A2(n_535),
.B(n_536),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_784),
.A2(n_555),
.B(n_617),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_688),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_688),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_757),
.A2(n_644),
.B1(n_530),
.B2(n_614),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_785),
.A2(n_555),
.B(n_617),
.Y(n_907)
);

O2A1O1Ixp5_ASAP7_75t_L g908 ( 
.A1(n_762),
.A2(n_583),
.B(n_571),
.C(n_614),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_721),
.B(n_723),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_759),
.B(n_627),
.Y(n_910)
);

BUFx4f_ASAP7_75t_L g911 ( 
.A(n_749),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_714),
.Y(n_912)
);

O2A1O1Ixp5_ASAP7_75t_L g913 ( 
.A1(n_778),
.A2(n_635),
.B(n_530),
.C(n_613),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_786),
.A2(n_666),
.B(n_607),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_809),
.B(n_613),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_723),
.B(n_644),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_732),
.A2(n_308),
.B1(n_307),
.B2(n_292),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_727),
.B(n_644),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_695),
.A2(n_626),
.B(n_638),
.C(n_330),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_691),
.Y(n_920)
);

NOR2xp67_ASAP7_75t_SL g921 ( 
.A(n_807),
.B(n_301),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_691),
.B(n_736),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_735),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_809),
.B(n_626),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_727),
.B(n_638),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_691),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_691),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_736),
.B(n_607),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_712),
.B(n_558),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_720),
.B(n_558),
.Y(n_930)
);

AND2x6_ASAP7_75t_L g931 ( 
.A(n_757),
.B(n_607),
.Y(n_931)
);

OAI321xp33_ASAP7_75t_L g932 ( 
.A1(n_771),
.A2(n_331),
.A3(n_263),
.B1(n_342),
.B2(n_305),
.C(n_310),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_746),
.A2(n_760),
.B(n_741),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_823),
.B(n_612),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_714),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_779),
.B(n_612),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_709),
.B(n_558),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_740),
.A2(n_612),
.B1(n_323),
.B2(n_624),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_746),
.A2(n_612),
.B(n_624),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_760),
.A2(n_612),
.B(n_624),
.Y(n_940)
);

BUFx4f_ASAP7_75t_L g941 ( 
.A(n_749),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_711),
.B(n_558),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_722),
.A2(n_558),
.B1(n_597),
.B2(n_604),
.Y(n_943)
);

NOR2x1_ASAP7_75t_L g944 ( 
.A(n_706),
.B(n_478),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_831),
.B(n_558),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_831),
.B(n_683),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_697),
.A2(n_624),
.B(n_451),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_697),
.A2(n_624),
.B(n_458),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_681),
.A2(n_624),
.B(n_458),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_716),
.A2(n_604),
.B(n_597),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_681),
.A2(n_462),
.B(n_222),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_754),
.A2(n_462),
.B(n_224),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_795),
.A2(n_462),
.B(n_227),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_802),
.A2(n_297),
.B(n_235),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_804),
.A2(n_303),
.B(n_244),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_770),
.B(n_558),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_679),
.B(n_757),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_770),
.B(n_597),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_814),
.A2(n_304),
.B(n_246),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_737),
.B(n_597),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_737),
.B(n_597),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_756),
.A2(n_488),
.B1(n_482),
.B2(n_478),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_679),
.B(n_676),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_718),
.B(n_755),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_719),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_684),
.B(n_597),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_807),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_815),
.A2(n_825),
.B(n_816),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_719),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_826),
.A2(n_230),
.B(n_248),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_757),
.B(n_676),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_810),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_708),
.B(n_597),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_764),
.B(n_604),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_767),
.B(n_604),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_829),
.A2(n_800),
.B(n_837),
.Y(n_976)
);

NAND2x1p5_ASAP7_75t_L g977 ( 
.A(n_706),
.B(n_478),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_777),
.B(n_783),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_788),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_801),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_763),
.A2(n_604),
.B(n_452),
.Y(n_981)
);

OAI321xp33_ASAP7_75t_L g982 ( 
.A1(n_782),
.A2(n_752),
.A3(n_769),
.B1(n_738),
.B2(n_739),
.C(n_797),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_796),
.B(n_604),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_806),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_810),
.B(n_676),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_680),
.B(n_676),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_820),
.B(n_604),
.Y(n_987)
);

OAI21x1_ASAP7_75t_L g988 ( 
.A1(n_822),
.A2(n_287),
.B(n_491),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_750),
.B(n_495),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_680),
.B(n_293),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_811),
.B(n_495),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_800),
.A2(n_274),
.B(n_253),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_821),
.B(n_272),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_827),
.A2(n_273),
.B(n_291),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_843),
.A2(n_452),
.B(n_464),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_781),
.B(n_495),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_693),
.B(n_495),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_824),
.A2(n_693),
.B(n_774),
.C(n_707),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_749),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_801),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_842),
.A2(n_452),
.B(n_464),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_750),
.B(n_495),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_832),
.A2(n_836),
.B(n_794),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_778),
.A2(n_452),
.B(n_464),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_780),
.A2(n_452),
.B(n_464),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_819),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_819),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_835),
.B(n_17),
.Y(n_1008)
);

NAND2x1_ASAP7_75t_L g1009 ( 
.A(n_845),
.B(n_495),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_685),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_734),
.B(n_491),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_811),
.B(n_491),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_845),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_692),
.A2(n_452),
.B(n_488),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_808),
.B(n_824),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_694),
.B(n_491),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_780),
.A2(n_452),
.B(n_464),
.Y(n_1017)
);

OAI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_797),
.A2(n_491),
.B1(n_488),
.B2(n_482),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_789),
.A2(n_452),
.B(n_464),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_811),
.B(n_491),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_789),
.A2(n_464),
.B(n_455),
.Y(n_1021)
);

INVx4_ASAP7_75t_L g1022 ( 
.A(n_819),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_742),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_722),
.B(n_21),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_751),
.B(n_488),
.Y(n_1025)
);

INVx1_ASAP7_75t_SL g1026 ( 
.A(n_793),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_805),
.B(n_488),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_791),
.A2(n_21),
.B(n_26),
.C(n_28),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_797),
.Y(n_1029)
);

INVx4_ASAP7_75t_L g1030 ( 
.A(n_813),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_791),
.A2(n_455),
.B(n_239),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_839),
.B(n_482),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_844),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_794),
.A2(n_28),
.B(n_30),
.C(n_31),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_848),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_897),
.B(n_728),
.Y(n_1036)
);

INVx8_ASAP7_75t_L g1037 ( 
.A(n_931),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_855),
.B(n_861),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_855),
.A2(n_812),
.B(n_790),
.C(n_799),
.Y(n_1039)
);

NAND2x1p5_ASAP7_75t_L g1040 ( 
.A(n_1022),
.B(n_811),
.Y(n_1040)
);

NOR3xp33_ASAP7_75t_L g1041 ( 
.A(n_982),
.B(n_730),
.C(n_704),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_909),
.A2(n_841),
.B1(n_818),
.B2(n_828),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_910),
.B(n_861),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_853),
.Y(n_1044)
);

NOR3xp33_ASAP7_75t_L g1045 ( 
.A(n_849),
.B(n_704),
.C(n_689),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_854),
.B(n_728),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_1022),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_883),
.A2(n_812),
.B(n_845),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_893),
.B(n_728),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_1015),
.A2(n_798),
.B(n_817),
.C(n_818),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_857),
.B(n_748),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_853),
.B(n_869),
.Y(n_1052)
);

INVxp67_ASAP7_75t_SL g1053 ( 
.A(n_1018),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_847),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_877),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_872),
.A2(n_798),
.B(n_817),
.C(n_840),
.Y(n_1056)
);

CKINVDCx6p67_ASAP7_75t_R g1057 ( 
.A(n_1030),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_882),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_912),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_923),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_864),
.B(n_828),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_846),
.A2(n_841),
.B1(n_733),
.B2(n_813),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_884),
.A2(n_845),
.B(n_455),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_846),
.A2(n_833),
.B1(n_482),
.B2(n_478),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_1008),
.B(n_482),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_916),
.A2(n_455),
.B(n_239),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_979),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_984),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_SL g1069 ( 
.A1(n_921),
.A2(n_30),
.B(n_35),
.C(n_38),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_876),
.B(n_38),
.Y(n_1070)
);

NOR3xp33_ASAP7_75t_L g1071 ( 
.A(n_901),
.B(n_39),
.C(n_40),
.Y(n_1071)
);

NAND2x1p5_ASAP7_75t_L g1072 ( 
.A(n_911),
.B(n_482),
.Y(n_1072)
);

INVxp67_ASAP7_75t_L g1073 ( 
.A(n_946),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_1008),
.B(n_478),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_876),
.B(n_43),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_935),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_856),
.A2(n_287),
.B1(n_239),
.B2(n_455),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_886),
.A2(n_287),
.B(n_52),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_851),
.B(n_48),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_918),
.A2(n_97),
.B(n_175),
.Y(n_1080)
);

AOI22x1_ASAP7_75t_L g1081 ( 
.A1(n_968),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_891),
.A2(n_53),
.B(n_56),
.C(n_57),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_978),
.A2(n_58),
.B1(n_59),
.B2(n_287),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_R g1084 ( 
.A(n_911),
.B(n_106),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_941),
.B(n_287),
.Y(n_1085)
);

O2A1O1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_862),
.A2(n_59),
.B(n_287),
.C(n_66),
.Y(n_1086)
);

CKINVDCx10_ASAP7_75t_R g1087 ( 
.A(n_892),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_925),
.A2(n_61),
.B(n_69),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_870),
.A2(n_76),
.B(n_82),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_965),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_915),
.A2(n_287),
.B(n_84),
.C(n_86),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1010),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_879),
.A2(n_83),
.B(n_88),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_969),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_915),
.A2(n_89),
.B(n_103),
.C(n_104),
.Y(n_1095)
);

NOR3xp33_ASAP7_75t_L g1096 ( 
.A(n_862),
.B(n_111),
.C(n_118),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_868),
.B(n_122),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_914),
.A2(n_899),
.B(n_924),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_946),
.B(n_123),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_SL g1100 ( 
.A(n_1030),
.B(n_125),
.Y(n_1100)
);

OAI21xp33_ASAP7_75t_SL g1101 ( 
.A1(n_899),
.A2(n_135),
.B(n_138),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_1026),
.B(n_155),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_924),
.A2(n_168),
.B(n_171),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_964),
.B(n_1029),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_858),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_980),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_904),
.B(n_173),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_892),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_858),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_894),
.B(n_1024),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_904),
.B(n_920),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_874),
.A2(n_866),
.B(n_998),
.C(n_936),
.Y(n_1112)
);

AOI221x1_ASAP7_75t_L g1113 ( 
.A1(n_1003),
.A2(n_976),
.B1(n_960),
.B2(n_961),
.C(n_871),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_885),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_973),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1023),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_989),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_852),
.A2(n_887),
.B(n_933),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1033),
.Y(n_1119)
);

OR2x6_ASAP7_75t_L g1120 ( 
.A(n_934),
.B(n_956),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_936),
.A2(n_896),
.B(n_1034),
.C(n_1028),
.Y(n_1121)
);

O2A1O1Ixp5_ASAP7_75t_L g1122 ( 
.A1(n_860),
.A2(n_997),
.B(n_886),
.C(n_900),
.Y(n_1122)
);

NAND2xp33_ASAP7_75t_L g1123 ( 
.A(n_904),
.B(n_920),
.Y(n_1123)
);

OA22x2_ASAP7_75t_L g1124 ( 
.A1(n_990),
.A2(n_943),
.B1(n_958),
.B2(n_930),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_859),
.B(n_945),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_920),
.B(n_926),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_945),
.B(n_863),
.Y(n_1127)
);

NAND3xp33_ASAP7_75t_L g1128 ( 
.A(n_992),
.B(n_919),
.C(n_994),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_881),
.A2(n_878),
.B(n_880),
.Y(n_1129)
);

INVxp33_ASAP7_75t_SL g1130 ( 
.A(n_1024),
.Y(n_1130)
);

NAND2xp33_ASAP7_75t_SL g1131 ( 
.A(n_926),
.B(n_999),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1000),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_926),
.B(n_1018),
.Y(n_1133)
);

CKINVDCx8_ASAP7_75t_R g1134 ( 
.A(n_931),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_889),
.A2(n_867),
.B1(n_993),
.B2(n_929),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_850),
.A2(n_1002),
.B1(n_867),
.B2(n_917),
.Y(n_1136)
);

AOI221xp5_ASAP7_75t_L g1137 ( 
.A1(n_932),
.A2(n_908),
.B1(n_875),
.B2(n_996),
.C(n_873),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_902),
.A2(n_907),
.B(n_903),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_999),
.B(n_1006),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_888),
.A2(n_898),
.B(n_865),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_908),
.A2(n_942),
.B(n_937),
.C(n_900),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1016),
.Y(n_1142)
);

NAND2xp33_ASAP7_75t_R g1143 ( 
.A(n_1006),
.B(n_1007),
.Y(n_1143)
);

OR2x2_ASAP7_75t_L g1144 ( 
.A(n_1007),
.B(n_927),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_913),
.A2(n_966),
.B(n_950),
.C(n_974),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1025),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_967),
.B(n_972),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_913),
.A2(n_957),
.B(n_987),
.C(n_983),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_885),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_SL g1150 ( 
.A1(n_967),
.A2(n_972),
.B(n_953),
.C(n_959),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_939),
.A2(n_940),
.B(n_1011),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_926),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_905),
.B(n_927),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_952),
.A2(n_963),
.B(n_895),
.Y(n_1154)
);

OA21x2_ASAP7_75t_L g1155 ( 
.A1(n_988),
.A2(n_1021),
.B(n_1031),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1013),
.B(n_906),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1013),
.B(n_906),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1013),
.B(n_957),
.Y(n_1158)
);

AO21x1_ASAP7_75t_L g1159 ( 
.A1(n_991),
.A2(n_1020),
.B(n_986),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_963),
.A2(n_949),
.B(n_948),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_931),
.B(n_922),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_931),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_947),
.A2(n_985),
.B(n_975),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_971),
.B(n_931),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_966),
.A2(n_995),
.B(n_1014),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_890),
.A2(n_928),
.B(n_962),
.C(n_970),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1027),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_977),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_977),
.Y(n_1169)
);

HB1xp67_ASAP7_75t_L g1170 ( 
.A(n_991),
.Y(n_1170)
);

NAND3xp33_ASAP7_75t_L g1171 ( 
.A(n_954),
.B(n_955),
.C(n_938),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1020),
.B(n_1012),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_971),
.A2(n_944),
.B1(n_1009),
.B2(n_981),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1032),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_951),
.A2(n_1004),
.B(n_1005),
.C(n_1017),
.Y(n_1175)
);

AOI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1019),
.A2(n_860),
.B(n_976),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1001),
.B(n_701),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_848),
.Y(n_1178)
);

BUFx4f_ASAP7_75t_L g1179 ( 
.A(n_999),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_909),
.A2(n_884),
.B(n_883),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_853),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_909),
.A2(n_1015),
.B(n_857),
.C(n_854),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_853),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_882),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_1013),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_897),
.B(n_591),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_897),
.B(n_591),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_897),
.B(n_591),
.Y(n_1188)
);

NOR2xp67_ASAP7_75t_L g1189 ( 
.A(n_1058),
.B(n_1184),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1182),
.A2(n_1098),
.B(n_1180),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1108),
.B(n_1047),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_SL g1192 ( 
.A1(n_1130),
.A2(n_1038),
.B1(n_1079),
.B2(n_1070),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_1044),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1038),
.A2(n_1182),
.B(n_1041),
.C(n_1045),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_1113),
.A2(n_1112),
.A3(n_1159),
.B(n_1145),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1051),
.B(n_1043),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1186),
.B(n_1187),
.Y(n_1197)
);

AOI31xp67_ASAP7_75t_L g1198 ( 
.A1(n_1124),
.A2(n_1158),
.A3(n_1133),
.B(n_1136),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1118),
.A2(n_1138),
.B(n_1129),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_1181),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1151),
.A2(n_1160),
.B(n_1140),
.Y(n_1201)
);

INVx5_ASAP7_75t_L g1202 ( 
.A(n_1037),
.Y(n_1202)
);

NOR2xp67_ASAP7_75t_L g1203 ( 
.A(n_1073),
.B(n_1104),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1188),
.B(n_1073),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1054),
.Y(n_1205)
);

AOI221x1_ASAP7_75t_L g1206 ( 
.A1(n_1071),
.A2(n_1041),
.B1(n_1045),
.B2(n_1096),
.C(n_1078),
.Y(n_1206)
);

O2A1O1Ixp5_ASAP7_75t_L g1207 ( 
.A1(n_1065),
.A2(n_1074),
.B(n_1122),
.C(n_1121),
.Y(n_1207)
);

AO32x2_ASAP7_75t_L g1208 ( 
.A1(n_1083),
.A2(n_1135),
.A3(n_1042),
.B1(n_1064),
.B2(n_1062),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1175),
.A2(n_1141),
.B(n_1127),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1141),
.A2(n_1127),
.B(n_1053),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_SL g1211 ( 
.A1(n_1050),
.A2(n_1053),
.B(n_1125),
.Y(n_1211)
);

O2A1O1Ixp33_ASAP7_75t_SL g1212 ( 
.A1(n_1150),
.A2(n_1075),
.B(n_1039),
.C(n_1091),
.Y(n_1212)
);

BUFx10_ASAP7_75t_L g1213 ( 
.A(n_1102),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_SL g1214 ( 
.A1(n_1052),
.A2(n_1069),
.B(n_1095),
.C(n_1147),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_SL g1215 ( 
.A1(n_1082),
.A2(n_1107),
.B(n_1111),
.C(n_1126),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1104),
.B(n_1183),
.Y(n_1216)
);

NAND3xp33_ASAP7_75t_L g1217 ( 
.A(n_1071),
.B(n_1086),
.C(n_1096),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1061),
.B(n_1079),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1110),
.B(n_1060),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1063),
.A2(n_1066),
.B(n_1163),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1050),
.A2(n_1165),
.B(n_1154),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_R g1222 ( 
.A(n_1087),
.B(n_1143),
.Y(n_1222)
);

AO31x2_ASAP7_75t_L g1223 ( 
.A1(n_1046),
.A2(n_1048),
.A3(n_1174),
.B(n_1146),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1067),
.B(n_1068),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1049),
.B(n_1036),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1125),
.B(n_1092),
.Y(n_1226)
);

BUFx2_ASAP7_75t_SL g1227 ( 
.A(n_1134),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1055),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1093),
.A2(n_1101),
.B(n_1123),
.Y(n_1229)
);

INVx2_ASAP7_75t_SL g1230 ( 
.A(n_1057),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1137),
.A2(n_1103),
.B(n_1171),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1116),
.B(n_1119),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1084),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1176),
.A2(n_1122),
.B(n_1148),
.Y(n_1234)
);

OR2x6_ASAP7_75t_L g1235 ( 
.A(n_1037),
.B(n_1040),
.Y(n_1235)
);

AOI221x1_ASAP7_75t_L g1236 ( 
.A1(n_1128),
.A2(n_1172),
.B1(n_1097),
.B2(n_1089),
.C(n_1080),
.Y(n_1236)
);

AO22x1_ASAP7_75t_L g1237 ( 
.A1(n_1102),
.A2(n_1099),
.B1(n_1164),
.B2(n_1047),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1037),
.A2(n_1148),
.B(n_1155),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1059),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1076),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1155),
.A2(n_1056),
.B(n_1166),
.Y(n_1241)
);

O2A1O1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1086),
.A2(n_1082),
.B(n_1056),
.C(n_1177),
.Y(n_1242)
);

INVxp67_ASAP7_75t_L g1243 ( 
.A(n_1117),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1170),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1166),
.A2(n_1088),
.B(n_1173),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1115),
.B(n_1094),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1170),
.A2(n_1142),
.B(n_1167),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1144),
.B(n_1139),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1157),
.Y(n_1249)
);

INVx5_ASAP7_75t_SL g1250 ( 
.A(n_1185),
.Y(n_1250)
);

OAI22x1_ASAP7_75t_L g1251 ( 
.A1(n_1081),
.A2(n_1077),
.B1(n_1164),
.B2(n_1156),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1090),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1161),
.A2(n_1178),
.B(n_1106),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1179),
.A2(n_1072),
.B1(n_1120),
.B2(n_1149),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1179),
.A2(n_1072),
.B1(n_1120),
.B2(n_1149),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1152),
.B(n_1040),
.Y(n_1256)
);

INVx4_ASAP7_75t_L g1257 ( 
.A(n_1162),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1162),
.A2(n_1168),
.B(n_1153),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1120),
.B(n_1169),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1168),
.A2(n_1109),
.B(n_1114),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1105),
.A2(n_1109),
.B(n_1114),
.Y(n_1261)
);

AO31x2_ASAP7_75t_L g1262 ( 
.A1(n_1185),
.A2(n_1100),
.A3(n_1131),
.B(n_1085),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1182),
.A2(n_1098),
.B(n_909),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1038),
.B(n_1043),
.Y(n_1264)
);

OAI22x1_ASAP7_75t_L g1265 ( 
.A1(n_1038),
.A2(n_894),
.B1(n_576),
.B2(n_1079),
.Y(n_1265)
);

OR2x6_ASAP7_75t_L g1266 ( 
.A(n_1037),
.B(n_749),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1038),
.A2(n_855),
.B(n_861),
.C(n_1182),
.Y(n_1267)
);

INVx2_ASAP7_75t_SL g1268 ( 
.A(n_1087),
.Y(n_1268)
);

O2A1O1Ixp5_ASAP7_75t_L g1269 ( 
.A1(n_1038),
.A2(n_1078),
.B(n_860),
.C(n_1098),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1113),
.A2(n_1129),
.B(n_1138),
.Y(n_1270)
);

OAI22x1_ASAP7_75t_L g1271 ( 
.A1(n_1038),
.A2(n_894),
.B1(n_576),
.B2(n_1079),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1038),
.A2(n_855),
.B(n_861),
.C(n_1182),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1134),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1038),
.B(n_1043),
.Y(n_1274)
);

BUFx10_ASAP7_75t_L g1275 ( 
.A(n_1184),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1035),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1182),
.A2(n_1098),
.B(n_909),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1134),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1108),
.B(n_1022),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1108),
.B(n_1022),
.Y(n_1280)
);

AO32x2_ASAP7_75t_L g1281 ( 
.A1(n_1083),
.A2(n_1135),
.A3(n_1042),
.B1(n_1064),
.B2(n_1062),
.Y(n_1281)
);

OA21x2_ASAP7_75t_L g1282 ( 
.A1(n_1113),
.A2(n_1129),
.B(n_1138),
.Y(n_1282)
);

INVx2_ASAP7_75t_SL g1283 ( 
.A(n_1087),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1038),
.B(n_1043),
.Y(n_1284)
);

NOR2x1_ASAP7_75t_R g1285 ( 
.A(n_1184),
.B(n_699),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1038),
.B(n_699),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1184),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1037),
.Y(n_1288)
);

O2A1O1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1038),
.A2(n_861),
.B(n_855),
.C(n_1051),
.Y(n_1289)
);

BUFx10_ASAP7_75t_L g1290 ( 
.A(n_1184),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1118),
.A2(n_1140),
.B(n_1129),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1182),
.A2(n_1098),
.B(n_909),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1134),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1038),
.A2(n_909),
.B1(n_1051),
.B2(n_1053),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_SL g1295 ( 
.A(n_1184),
.B(n_699),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1035),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1038),
.A2(n_909),
.B1(n_1051),
.B2(n_1053),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1182),
.A2(n_1098),
.B(n_909),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1054),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1038),
.A2(n_699),
.B1(n_554),
.B2(n_1130),
.Y(n_1300)
);

OR2x6_ASAP7_75t_L g1301 ( 
.A(n_1037),
.B(n_749),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1038),
.B(n_699),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_1044),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1038),
.B(n_699),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1054),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1038),
.B(n_1051),
.Y(n_1306)
);

INVx4_ASAP7_75t_L g1307 ( 
.A(n_1184),
.Y(n_1307)
);

A2O1A1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1038),
.A2(n_855),
.B(n_861),
.C(n_1182),
.Y(n_1308)
);

O2A1O1Ixp5_ASAP7_75t_L g1309 ( 
.A1(n_1038),
.A2(n_1078),
.B(n_860),
.C(n_1098),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_1044),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1038),
.A2(n_855),
.B(n_861),
.C(n_1182),
.Y(n_1311)
);

O2A1O1Ixp33_ASAP7_75t_SL g1312 ( 
.A1(n_1038),
.A2(n_909),
.B(n_1182),
.C(n_869),
.Y(n_1312)
);

INVx5_ASAP7_75t_L g1313 ( 
.A(n_1037),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1182),
.A2(n_1098),
.B(n_909),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1054),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1132),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1038),
.B(n_1043),
.Y(n_1317)
);

A2O1A1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1038),
.A2(n_855),
.B(n_861),
.C(n_1182),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1045),
.A2(n_728),
.B1(n_775),
.B2(n_382),
.Y(n_1319)
);

BUFx10_ASAP7_75t_L g1320 ( 
.A(n_1184),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1182),
.A2(n_1098),
.B(n_909),
.Y(n_1321)
);

BUFx10_ASAP7_75t_L g1322 ( 
.A(n_1184),
.Y(n_1322)
);

OA21x2_ASAP7_75t_L g1323 ( 
.A1(n_1113),
.A2(n_1129),
.B(n_1138),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_1184),
.Y(n_1324)
);

AO21x1_ASAP7_75t_L g1325 ( 
.A1(n_1086),
.A2(n_1041),
.B(n_1182),
.Y(n_1325)
);

OAI21xp33_ASAP7_75t_L g1326 ( 
.A1(n_1038),
.A2(n_861),
.B(n_855),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1182),
.A2(n_1098),
.B(n_909),
.Y(n_1327)
);

A2O1A1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1038),
.A2(n_855),
.B(n_861),
.C(n_1182),
.Y(n_1328)
);

BUFx10_ASAP7_75t_L g1329 ( 
.A(n_1184),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_SL g1330 ( 
.A1(n_1182),
.A2(n_909),
.B(n_745),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1182),
.A2(n_1098),
.B(n_909),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1182),
.A2(n_1098),
.B(n_909),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1043),
.B(n_701),
.Y(n_1333)
);

O2A1O1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1038),
.A2(n_861),
.B(n_855),
.C(n_1051),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1038),
.B(n_1043),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1182),
.A2(n_1098),
.B(n_909),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1182),
.A2(n_1098),
.B(n_909),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1038),
.B(n_1043),
.Y(n_1338)
);

AO31x2_ASAP7_75t_L g1339 ( 
.A1(n_1113),
.A2(n_860),
.A3(n_1112),
.B(n_1159),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1035),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1288),
.Y(n_1341)
);

CKINVDCx11_ASAP7_75t_R g1342 ( 
.A(n_1275),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1319),
.A2(n_1192),
.B1(n_1217),
.B2(n_1265),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1224),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1267),
.A2(n_1308),
.B1(n_1311),
.B2(n_1318),
.Y(n_1345)
);

CKINVDCx16_ASAP7_75t_R g1346 ( 
.A(n_1222),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1324),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1205),
.Y(n_1348)
);

INVx3_ASAP7_75t_L g1349 ( 
.A(n_1288),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1272),
.A2(n_1328),
.B1(n_1326),
.B2(n_1194),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1288),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1275),
.Y(n_1352)
);

INVx4_ASAP7_75t_L g1353 ( 
.A(n_1307),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1302),
.B(n_1304),
.Y(n_1354)
);

BUFx4_ASAP7_75t_R g1355 ( 
.A(n_1213),
.Y(n_1355)
);

INVx5_ASAP7_75t_L g1356 ( 
.A(n_1266),
.Y(n_1356)
);

BUFx4_ASAP7_75t_SL g1357 ( 
.A(n_1233),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1299),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1305),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1264),
.A2(n_1284),
.B1(n_1317),
.B2(n_1274),
.Y(n_1360)
);

CKINVDCx6p67_ASAP7_75t_R g1361 ( 
.A(n_1290),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_1193),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1200),
.Y(n_1363)
);

BUFx4f_ASAP7_75t_L g1364 ( 
.A(n_1273),
.Y(n_1364)
);

INVx3_ASAP7_75t_L g1365 ( 
.A(n_1202),
.Y(n_1365)
);

OAI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1218),
.A2(n_1300),
.B1(n_1338),
.B2(n_1335),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1271),
.A2(n_1325),
.B1(n_1213),
.B2(n_1294),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_SL g1368 ( 
.A1(n_1297),
.A2(n_1226),
.B1(n_1219),
.B2(n_1206),
.Y(n_1368)
);

INVx4_ASAP7_75t_L g1369 ( 
.A(n_1307),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1249),
.A2(n_1306),
.B1(n_1196),
.B2(n_1225),
.Y(n_1370)
);

BUFx2_ASAP7_75t_SL g1371 ( 
.A(n_1189),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1228),
.A2(n_1340),
.B1(n_1296),
.B2(n_1276),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1290),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1216),
.B(n_1333),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1315),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_1268),
.Y(n_1376)
);

BUFx12f_ASAP7_75t_L g1377 ( 
.A(n_1283),
.Y(n_1377)
);

BUFx8_ASAP7_75t_L g1378 ( 
.A(n_1230),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1239),
.A2(n_1240),
.B1(n_1252),
.B2(n_1246),
.Y(n_1379)
);

CKINVDCx11_ASAP7_75t_R g1380 ( 
.A(n_1320),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1316),
.Y(n_1381)
);

BUFx8_ASAP7_75t_L g1382 ( 
.A(n_1191),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1210),
.B(n_1289),
.Y(n_1383)
);

CKINVDCx11_ASAP7_75t_R g1384 ( 
.A(n_1320),
.Y(n_1384)
);

OAI22xp33_ASAP7_75t_SL g1385 ( 
.A1(n_1204),
.A2(n_1197),
.B1(n_1232),
.B2(n_1243),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1316),
.Y(n_1386)
);

BUFx4f_ASAP7_75t_SL g1387 ( 
.A(n_1322),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1334),
.A2(n_1211),
.B1(n_1263),
.B2(n_1337),
.Y(n_1388)
);

AOI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1203),
.A2(n_1295),
.B1(n_1303),
.B2(n_1310),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1231),
.A2(n_1253),
.B1(n_1247),
.B2(n_1227),
.Y(n_1390)
);

OAI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1273),
.A2(n_1293),
.B1(n_1278),
.B2(n_1313),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1312),
.B(n_1277),
.Y(n_1392)
);

CKINVDCx6p67_ASAP7_75t_R g1393 ( 
.A(n_1322),
.Y(n_1393)
);

INVx6_ASAP7_75t_L g1394 ( 
.A(n_1202),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_SL g1395 ( 
.A1(n_1208),
.A2(n_1281),
.B1(n_1209),
.B2(n_1278),
.Y(n_1395)
);

NAND2x1p5_ASAP7_75t_L g1396 ( 
.A(n_1202),
.B(n_1313),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1208),
.A2(n_1281),
.B1(n_1293),
.B2(n_1198),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1244),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1292),
.A2(n_1327),
.B1(n_1298),
.B2(n_1314),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1253),
.A2(n_1251),
.B1(n_1259),
.B2(n_1248),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1329),
.Y(n_1401)
);

OAI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1313),
.A2(n_1301),
.B1(n_1235),
.B2(n_1254),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1321),
.A2(n_1331),
.B1(n_1332),
.B2(n_1336),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_SL g1404 ( 
.A1(n_1208),
.A2(n_1281),
.B1(n_1259),
.B2(n_1245),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_SL g1405 ( 
.A(n_1191),
.Y(n_1405)
);

INVx8_ASAP7_75t_L g1406 ( 
.A(n_1301),
.Y(n_1406)
);

BUFx12f_ASAP7_75t_L g1407 ( 
.A(n_1329),
.Y(n_1407)
);

BUFx4f_ASAP7_75t_SL g1408 ( 
.A(n_1279),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1250),
.Y(n_1409)
);

BUFx12f_ASAP7_75t_L g1410 ( 
.A(n_1279),
.Y(n_1410)
);

BUFx2_ASAP7_75t_L g1411 ( 
.A(n_1280),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_SL g1412 ( 
.A1(n_1221),
.A2(n_1190),
.B1(n_1229),
.B2(n_1237),
.Y(n_1412)
);

INVx6_ASAP7_75t_L g1413 ( 
.A(n_1257),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1255),
.A2(n_1215),
.B1(n_1212),
.B2(n_1256),
.Y(n_1414)
);

INVx4_ASAP7_75t_SL g1415 ( 
.A(n_1262),
.Y(n_1415)
);

INVx4_ASAP7_75t_L g1416 ( 
.A(n_1257),
.Y(n_1416)
);

INVxp67_ASAP7_75t_SL g1417 ( 
.A(n_1270),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1242),
.A2(n_1241),
.B1(n_1330),
.B2(n_1309),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1238),
.A2(n_1258),
.B1(n_1250),
.B2(n_1260),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1223),
.B(n_1195),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1261),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1234),
.A2(n_1270),
.B1(n_1282),
.B2(n_1323),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1339),
.Y(n_1423)
);

CKINVDCx11_ASAP7_75t_R g1424 ( 
.A(n_1285),
.Y(n_1424)
);

OAI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1236),
.A2(n_1269),
.B1(n_1207),
.B2(n_1323),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1199),
.A2(n_1282),
.B1(n_1201),
.B2(n_1220),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1339),
.B(n_1291),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1214),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1319),
.A2(n_728),
.B1(n_1045),
.B2(n_1041),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1319),
.A2(n_728),
.B1(n_1045),
.B2(n_1041),
.Y(n_1430)
);

OAI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1218),
.A2(n_982),
.B1(n_1038),
.B2(n_1300),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1324),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1267),
.A2(n_1038),
.B1(n_1308),
.B2(n_1272),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1319),
.A2(n_728),
.B1(n_1045),
.B2(n_1041),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1267),
.A2(n_1038),
.B1(n_1308),
.B2(n_1272),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1192),
.A2(n_1130),
.B1(n_1038),
.B2(n_1286),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1319),
.A2(n_728),
.B1(n_1045),
.B2(n_1041),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_1275),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1216),
.B(n_1249),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1224),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1319),
.A2(n_728),
.B1(n_1045),
.B2(n_1041),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1192),
.A2(n_1130),
.B1(n_1038),
.B2(n_1286),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1288),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1224),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_1287),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1224),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1319),
.A2(n_728),
.B1(n_1045),
.B2(n_1041),
.Y(n_1447)
);

OAI22x1_ASAP7_75t_SL g1448 ( 
.A1(n_1268),
.A2(n_731),
.B1(n_1283),
.B2(n_699),
.Y(n_1448)
);

BUFx10_ASAP7_75t_L g1449 ( 
.A(n_1324),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1319),
.A2(n_728),
.B1(n_1045),
.B2(n_1041),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1267),
.A2(n_1038),
.B1(n_1308),
.B2(n_1272),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_SL g1452 ( 
.A1(n_1192),
.A2(n_728),
.B1(n_1038),
.B2(n_1053),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1218),
.A2(n_982),
.B1(n_1038),
.B2(n_1300),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_SL g1454 ( 
.A(n_1268),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_1275),
.Y(n_1455)
);

INVx2_ASAP7_75t_SL g1456 ( 
.A(n_1275),
.Y(n_1456)
);

INVx8_ASAP7_75t_L g1457 ( 
.A(n_1266),
.Y(n_1457)
);

OAI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1218),
.A2(n_982),
.B1(n_1038),
.B2(n_1300),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1192),
.A2(n_728),
.B1(n_1038),
.B2(n_1053),
.Y(n_1459)
);

INVxp67_ASAP7_75t_SL g1460 ( 
.A(n_1270),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1288),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1324),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1224),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1415),
.B(n_1421),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1381),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1386),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1399),
.A2(n_1403),
.B(n_1426),
.Y(n_1467)
);

INVx2_ASAP7_75t_SL g1468 ( 
.A(n_1398),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1363),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1404),
.B(n_1395),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1360),
.B(n_1374),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1439),
.B(n_1420),
.Y(n_1472)
);

BUFx3_ASAP7_75t_L g1473 ( 
.A(n_1382),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1354),
.B(n_1436),
.Y(n_1474)
);

OA21x2_ASAP7_75t_L g1475 ( 
.A1(n_1383),
.A2(n_1392),
.B(n_1422),
.Y(n_1475)
);

OA21x2_ASAP7_75t_L g1476 ( 
.A1(n_1383),
.A2(n_1392),
.B(n_1417),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1404),
.B(n_1395),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1348),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1452),
.A2(n_1459),
.B1(n_1429),
.B2(n_1434),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1411),
.Y(n_1480)
);

NAND3xp33_ASAP7_75t_L g1481 ( 
.A(n_1350),
.B(n_1451),
.C(n_1435),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1347),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1427),
.B(n_1358),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1359),
.B(n_1375),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1423),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1362),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1417),
.A2(n_1460),
.B(n_1426),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1360),
.B(n_1344),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1406),
.Y(n_1489)
);

CKINVDCx6p67_ASAP7_75t_R g1490 ( 
.A(n_1424),
.Y(n_1490)
);

AOI21xp33_ASAP7_75t_L g1491 ( 
.A1(n_1431),
.A2(n_1458),
.B(n_1453),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_SL g1492 ( 
.A1(n_1350),
.A2(n_1451),
.B1(n_1433),
.B2(n_1435),
.Y(n_1492)
);

INVx2_ASAP7_75t_SL g1493 ( 
.A(n_1406),
.Y(n_1493)
);

AOI21xp33_ASAP7_75t_SL g1494 ( 
.A1(n_1366),
.A2(n_1433),
.B(n_1442),
.Y(n_1494)
);

BUFx2_ASAP7_75t_SL g1495 ( 
.A(n_1356),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1399),
.Y(n_1496)
);

AOI21xp33_ASAP7_75t_L g1497 ( 
.A1(n_1385),
.A2(n_1367),
.B(n_1343),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1403),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1388),
.A2(n_1419),
.B(n_1345),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1457),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1440),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1388),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1444),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1446),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1463),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1397),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1397),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1428),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1345),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1405),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1418),
.B(n_1368),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1390),
.A2(n_1414),
.B(n_1400),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1405),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1412),
.Y(n_1514)
);

O2A1O1Ixp5_ASAP7_75t_L g1515 ( 
.A1(n_1425),
.A2(n_1391),
.B(n_1364),
.C(n_1416),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1412),
.Y(n_1516)
);

OR2x6_ASAP7_75t_L g1517 ( 
.A(n_1457),
.B(n_1396),
.Y(n_1517)
);

INVx4_ASAP7_75t_SL g1518 ( 
.A(n_1394),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1418),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1365),
.A2(n_1370),
.B(n_1341),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1368),
.Y(n_1521)
);

AOI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1355),
.A2(n_1455),
.B(n_1438),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1452),
.B(n_1459),
.Y(n_1523)
);

AO21x2_ASAP7_75t_L g1524 ( 
.A1(n_1402),
.A2(n_1389),
.B(n_1437),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1413),
.Y(n_1525)
);

INVx2_ASAP7_75t_SL g1526 ( 
.A(n_1457),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1379),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1372),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_1413),
.Y(n_1529)
);

OAI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1408),
.A2(n_1364),
.B1(n_1346),
.B2(n_1410),
.Y(n_1530)
);

INVx4_ASAP7_75t_L g1531 ( 
.A(n_1356),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1445),
.Y(n_1532)
);

INVx2_ASAP7_75t_SL g1533 ( 
.A(n_1356),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1430),
.B(n_1441),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1447),
.B(n_1450),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1349),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1351),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1443),
.Y(n_1538)
);

AOI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1401),
.A2(n_1456),
.B(n_1461),
.Y(n_1539)
);

BUFx12f_ASAP7_75t_L g1540 ( 
.A(n_1342),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1353),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1471),
.B(n_1369),
.Y(n_1542)
);

OAI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1481),
.A2(n_1409),
.B(n_1352),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1539),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1494),
.B(n_1353),
.Y(n_1545)
);

A2O1A1Ixp33_ASAP7_75t_L g1546 ( 
.A1(n_1491),
.A2(n_1371),
.B(n_1373),
.C(n_1462),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1539),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1501),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1480),
.B(n_1369),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1480),
.B(n_1432),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1464),
.B(n_1361),
.Y(n_1551)
);

A2O1A1Ixp33_ASAP7_75t_L g1552 ( 
.A1(n_1494),
.A2(n_1481),
.B(n_1511),
.C(n_1521),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1469),
.B(n_1393),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1488),
.B(n_1378),
.Y(n_1554)
);

A2O1A1Ixp33_ASAP7_75t_L g1555 ( 
.A1(n_1511),
.A2(n_1521),
.B(n_1492),
.C(n_1497),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1486),
.B(n_1449),
.Y(n_1556)
);

O2A1O1Ixp33_ASAP7_75t_L g1557 ( 
.A1(n_1514),
.A2(n_1376),
.B(n_1448),
.C(n_1387),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1478),
.Y(n_1558)
);

AOI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1523),
.A2(n_1454),
.B1(n_1407),
.B2(n_1380),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1480),
.B(n_1384),
.Y(n_1560)
);

A2O1A1Ixp33_ASAP7_75t_L g1561 ( 
.A1(n_1523),
.A2(n_1470),
.B(n_1477),
.C(n_1499),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1532),
.B(n_1377),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1483),
.B(n_1454),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1478),
.Y(n_1564)
);

BUFx6f_ASAP7_75t_SL g1565 ( 
.A(n_1473),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1509),
.A2(n_1357),
.B1(n_1474),
.B2(n_1519),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1479),
.A2(n_1535),
.B1(n_1470),
.B2(n_1477),
.Y(n_1567)
);

OA21x2_ASAP7_75t_L g1568 ( 
.A1(n_1467),
.A2(n_1499),
.B(n_1512),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1483),
.B(n_1484),
.Y(n_1569)
);

OA21x2_ASAP7_75t_L g1570 ( 
.A1(n_1467),
.A2(n_1512),
.B(n_1496),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1468),
.B(n_1472),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1464),
.B(n_1518),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1503),
.B(n_1504),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1519),
.A2(n_1514),
.B1(n_1516),
.B2(n_1502),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1490),
.Y(n_1575)
);

BUFx4f_ASAP7_75t_SL g1576 ( 
.A(n_1540),
.Y(n_1576)
);

OR2x6_ASAP7_75t_L g1577 ( 
.A(n_1495),
.B(n_1510),
.Y(n_1577)
);

OAI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1516),
.A2(n_1515),
.B(n_1502),
.Y(n_1578)
);

A2O1A1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1535),
.A2(n_1506),
.B(n_1507),
.C(n_1534),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1508),
.B(n_1522),
.Y(n_1580)
);

AOI221xp5_ASAP7_75t_L g1581 ( 
.A1(n_1506),
.A2(n_1507),
.B1(n_1504),
.B2(n_1503),
.C(n_1505),
.Y(n_1581)
);

INVxp33_ASAP7_75t_L g1582 ( 
.A(n_1525),
.Y(n_1582)
);

O2A1O1Ixp33_ASAP7_75t_SL g1583 ( 
.A1(n_1530),
.A2(n_1496),
.B(n_1498),
.C(n_1541),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1522),
.B(n_1541),
.Y(n_1584)
);

A2O1A1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1527),
.A2(n_1520),
.B(n_1513),
.C(n_1510),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1476),
.A2(n_1487),
.B(n_1475),
.Y(n_1586)
);

BUFx4f_ASAP7_75t_L g1587 ( 
.A(n_1517),
.Y(n_1587)
);

A2O1A1Ixp33_ASAP7_75t_L g1588 ( 
.A1(n_1527),
.A2(n_1520),
.B(n_1489),
.C(n_1500),
.Y(n_1588)
);

AO32x2_ASAP7_75t_L g1589 ( 
.A1(n_1533),
.A2(n_1531),
.A3(n_1526),
.B1(n_1493),
.B2(n_1475),
.Y(n_1589)
);

OAI211xp5_ASAP7_75t_L g1590 ( 
.A1(n_1475),
.A2(n_1536),
.B(n_1537),
.C(n_1476),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1529),
.B(n_1538),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1464),
.B(n_1518),
.Y(n_1592)
);

AO32x2_ASAP7_75t_L g1593 ( 
.A1(n_1533),
.A2(n_1531),
.A3(n_1526),
.B1(n_1475),
.B2(n_1476),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1558),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1589),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1564),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1580),
.B(n_1476),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1569),
.B(n_1487),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1571),
.B(n_1487),
.Y(n_1599)
);

INVxp67_ASAP7_75t_L g1600 ( 
.A(n_1580),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1589),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1570),
.B(n_1568),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1572),
.B(n_1592),
.Y(n_1603)
);

INVxp67_ASAP7_75t_SL g1604 ( 
.A(n_1586),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1568),
.B(n_1487),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1589),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1568),
.B(n_1465),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1593),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1548),
.B(n_1465),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1593),
.B(n_1466),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1593),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1593),
.B(n_1485),
.Y(n_1612)
);

BUFx2_ASAP7_75t_L g1613 ( 
.A(n_1549),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1573),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1590),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1584),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1567),
.A2(n_1524),
.B1(n_1528),
.B2(n_1540),
.Y(n_1617)
);

OAI221xp5_ASAP7_75t_SL g1618 ( 
.A1(n_1615),
.A2(n_1552),
.B1(n_1555),
.B2(n_1561),
.C(n_1567),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1599),
.B(n_1542),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1598),
.B(n_1582),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1617),
.A2(n_1552),
.B1(n_1561),
.B2(n_1555),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1605),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1605),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1614),
.B(n_1615),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1617),
.A2(n_1524),
.B1(n_1574),
.B2(n_1578),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1603),
.B(n_1592),
.Y(n_1626)
);

AOI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1595),
.A2(n_1524),
.B1(n_1579),
.B2(n_1566),
.Y(n_1627)
);

INVx5_ASAP7_75t_L g1628 ( 
.A(n_1605),
.Y(n_1628)
);

OAI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1604),
.A2(n_1579),
.B1(n_1546),
.B2(n_1581),
.C(n_1588),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1614),
.B(n_1544),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1595),
.A2(n_1563),
.B1(n_1528),
.B2(n_1565),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1607),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1594),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1594),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1594),
.Y(n_1635)
);

NOR2x1_ASAP7_75t_SL g1636 ( 
.A(n_1599),
.B(n_1577),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1596),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1601),
.B(n_1591),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1597),
.B(n_1544),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1601),
.B(n_1585),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1599),
.B(n_1547),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1600),
.B(n_1554),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1603),
.B(n_1551),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1609),
.Y(n_1644)
);

AOI221xp5_ASAP7_75t_L g1645 ( 
.A1(n_1600),
.A2(n_1546),
.B1(n_1583),
.B2(n_1557),
.C(n_1543),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1608),
.A2(n_1611),
.B1(n_1606),
.B2(n_1604),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1612),
.Y(n_1647)
);

NAND2x1p5_ASAP7_75t_L g1648 ( 
.A(n_1628),
.B(n_1587),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1622),
.Y(n_1649)
);

INVxp67_ASAP7_75t_SL g1650 ( 
.A(n_1624),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1647),
.B(n_1610),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1633),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1624),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1644),
.B(n_1610),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1628),
.B(n_1606),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1647),
.B(n_1597),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1644),
.B(n_1610),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1619),
.B(n_1616),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1634),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1630),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1647),
.B(n_1608),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1639),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1628),
.B(n_1606),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1628),
.B(n_1636),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1628),
.B(n_1606),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1619),
.B(n_1616),
.Y(n_1666)
);

INVx1_ASAP7_75t_SL g1667 ( 
.A(n_1630),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1622),
.B(n_1611),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1635),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1623),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1646),
.B(n_1611),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_SL g1672 ( 
.A(n_1629),
.B(n_1575),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1620),
.B(n_1613),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1637),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1653),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1674),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1674),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1670),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1659),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1653),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1664),
.B(n_1626),
.Y(n_1681)
);

AND2x4_ASAP7_75t_SL g1682 ( 
.A(n_1664),
.B(n_1643),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1664),
.B(n_1626),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1671),
.B(n_1646),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1668),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1671),
.B(n_1658),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1668),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1671),
.B(n_1619),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1668),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1659),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1659),
.Y(n_1691)
);

INVxp67_ASAP7_75t_SL g1692 ( 
.A(n_1672),
.Y(n_1692)
);

OR2x2_ASAP7_75t_SL g1693 ( 
.A(n_1656),
.B(n_1632),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1672),
.A2(n_1629),
.B(n_1621),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1652),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1652),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1649),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1664),
.B(n_1626),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1649),
.Y(n_1699)
);

OAI221xp5_ASAP7_75t_L g1700 ( 
.A1(n_1650),
.A2(n_1618),
.B1(n_1627),
.B2(n_1621),
.C(n_1640),
.Y(n_1700)
);

NAND2xp33_ASAP7_75t_L g1701 ( 
.A(n_1648),
.B(n_1575),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1664),
.B(n_1626),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1664),
.B(n_1626),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1658),
.B(n_1639),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1666),
.B(n_1641),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1666),
.B(n_1650),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1662),
.B(n_1638),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1662),
.B(n_1576),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1651),
.B(n_1643),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1656),
.B(n_1641),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1686),
.B(n_1656),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1682),
.B(n_1651),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1694),
.B(n_1660),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1676),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1686),
.B(n_1654),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1692),
.B(n_1645),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1682),
.B(n_1709),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1676),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1675),
.B(n_1660),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1700),
.A2(n_1618),
.B(n_1640),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1682),
.B(n_1651),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1677),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1680),
.B(n_1706),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1706),
.B(n_1654),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1704),
.B(n_1657),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1708),
.B(n_1576),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1688),
.B(n_1667),
.Y(n_1727)
);

INVx1_ASAP7_75t_SL g1728 ( 
.A(n_1684),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1709),
.B(n_1673),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1681),
.B(n_1673),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1681),
.B(n_1673),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1704),
.B(n_1657),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1693),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1677),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1683),
.B(n_1661),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1688),
.B(n_1667),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1695),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1705),
.B(n_1640),
.Y(n_1738)
);

INVx2_ASAP7_75t_SL g1739 ( 
.A(n_1705),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1684),
.B(n_1669),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1683),
.B(n_1661),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1707),
.B(n_1638),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1693),
.B(n_1661),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_R g1744 ( 
.A(n_1701),
.B(n_1482),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1710),
.B(n_1642),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1710),
.B(n_1670),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1739),
.B(n_1685),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1726),
.B(n_1642),
.Y(n_1748)
);

OAI32xp33_ASAP7_75t_L g1749 ( 
.A1(n_1733),
.A2(n_1743),
.A3(n_1716),
.B1(n_1713),
.B2(n_1738),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1714),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1745),
.B(n_1685),
.Y(n_1751)
);

AOI221xp5_ASAP7_75t_L g1752 ( 
.A1(n_1716),
.A2(n_1645),
.B1(n_1678),
.B2(n_1602),
.C(n_1627),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1712),
.Y(n_1753)
);

OAI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1720),
.A2(n_1559),
.B(n_1625),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1718),
.Y(n_1755)
);

INVxp67_ASAP7_75t_L g1756 ( 
.A(n_1723),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1722),
.Y(n_1757)
);

INVx1_ASAP7_75t_SL g1758 ( 
.A(n_1728),
.Y(n_1758)
);

NAND4xp25_ASAP7_75t_L g1759 ( 
.A(n_1733),
.B(n_1545),
.C(n_1702),
.D(n_1698),
.Y(n_1759)
);

OAI21xp33_ASAP7_75t_L g1760 ( 
.A1(n_1743),
.A2(n_1689),
.B(n_1687),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1712),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1734),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1744),
.B(n_1698),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1737),
.Y(n_1764)
);

INVx6_ASAP7_75t_L g1765 ( 
.A(n_1717),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1739),
.A2(n_1625),
.B1(n_1631),
.B2(n_1655),
.Y(n_1766)
);

INVx2_ASAP7_75t_SL g1767 ( 
.A(n_1717),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1711),
.B(n_1565),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1740),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1740),
.B(n_1695),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1711),
.B(n_1687),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1727),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1758),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1767),
.B(n_1721),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1758),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1770),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1756),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1770),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1769),
.B(n_1736),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1747),
.B(n_1719),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1749),
.A2(n_1752),
.B(n_1754),
.Y(n_1781)
);

AOI22xp5_ASAP7_75t_SL g1782 ( 
.A1(n_1754),
.A2(n_1560),
.B1(n_1721),
.B2(n_1655),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1753),
.B(n_1729),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1765),
.A2(n_1729),
.B1(n_1731),
.B2(n_1730),
.Y(n_1784)
);

NAND3xp33_ASAP7_75t_L g1785 ( 
.A(n_1766),
.B(n_1724),
.C(n_1715),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1750),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1751),
.B(n_1735),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1755),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1761),
.B(n_1735),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_SL g1790 ( 
.A(n_1748),
.B(n_1730),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1772),
.B(n_1741),
.Y(n_1791)
);

A2O1A1Ixp33_ASAP7_75t_L g1792 ( 
.A1(n_1766),
.A2(n_1724),
.B(n_1655),
.C(n_1663),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1783),
.B(n_1765),
.Y(n_1793)
);

INVx1_ASAP7_75t_SL g1794 ( 
.A(n_1777),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1773),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1775),
.B(n_1771),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1777),
.Y(n_1797)
);

AOI221x1_ASAP7_75t_L g1798 ( 
.A1(n_1781),
.A2(n_1764),
.B1(n_1757),
.B2(n_1762),
.C(n_1759),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1783),
.B(n_1790),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1779),
.Y(n_1800)
);

OAI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1785),
.A2(n_1768),
.B1(n_1763),
.B2(n_1742),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1791),
.B(n_1725),
.Y(n_1802)
);

XNOR2xp5_ASAP7_75t_L g1803 ( 
.A(n_1782),
.B(n_1560),
.Y(n_1803)
);

AOI221xp5_ASAP7_75t_L g1804 ( 
.A1(n_1794),
.A2(n_1776),
.B1(n_1778),
.B2(n_1792),
.C(n_1788),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1794),
.A2(n_1790),
.B(n_1792),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1793),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1799),
.B(n_1774),
.Y(n_1807)
);

OAI21xp5_ASAP7_75t_SL g1808 ( 
.A1(n_1798),
.A2(n_1784),
.B(n_1789),
.Y(n_1808)
);

NAND4xp25_ASAP7_75t_L g1809 ( 
.A(n_1796),
.B(n_1787),
.C(n_1780),
.D(n_1786),
.Y(n_1809)
);

OAI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1797),
.A2(n_1760),
.B(n_1731),
.Y(n_1810)
);

AOI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1801),
.A2(n_1746),
.B(n_1690),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1802),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1800),
.B(n_1741),
.Y(n_1813)
);

NOR2x1_ASAP7_75t_L g1814 ( 
.A(n_1812),
.B(n_1809),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1806),
.Y(n_1815)
);

OAI21xp33_ASAP7_75t_L g1816 ( 
.A1(n_1808),
.A2(n_1803),
.B(n_1795),
.Y(n_1816)
);

AOI211xp5_ASAP7_75t_L g1817 ( 
.A1(n_1805),
.A2(n_1746),
.B(n_1725),
.C(n_1732),
.Y(n_1817)
);

AOI221xp5_ASAP7_75t_L g1818 ( 
.A1(n_1804),
.A2(n_1678),
.B1(n_1665),
.B2(n_1663),
.C(n_1655),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1815),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1814),
.Y(n_1820)
);

AOI211xp5_ASAP7_75t_L g1821 ( 
.A1(n_1816),
.A2(n_1807),
.B(n_1810),
.C(n_1811),
.Y(n_1821)
);

OAI31xp33_ASAP7_75t_L g1822 ( 
.A1(n_1817),
.A2(n_1813),
.A3(n_1678),
.B(n_1665),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_SL g1823 ( 
.A1(n_1818),
.A2(n_1689),
.B1(n_1665),
.B2(n_1655),
.Y(n_1823)
);

INVx1_ASAP7_75t_SL g1824 ( 
.A(n_1814),
.Y(n_1824)
);

XNOR2x1_ASAP7_75t_L g1825 ( 
.A(n_1824),
.B(n_1562),
.Y(n_1825)
);

INVx3_ASAP7_75t_L g1826 ( 
.A(n_1819),
.Y(n_1826)
);

AOI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1820),
.A2(n_1821),
.B1(n_1823),
.B2(n_1655),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1822),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1819),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1826),
.B(n_1696),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1826),
.B(n_1702),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1825),
.Y(n_1832)
);

AOI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1832),
.A2(n_1828),
.B1(n_1829),
.B2(n_1831),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1833),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1834),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1834),
.A2(n_1830),
.B(n_1827),
.Y(n_1836)
);

OAI22xp33_ASAP7_75t_SL g1837 ( 
.A1(n_1835),
.A2(n_1697),
.B1(n_1699),
.B2(n_1691),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1836),
.B(n_1679),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1838),
.Y(n_1839)
);

INVx2_ASAP7_75t_SL g1840 ( 
.A(n_1837),
.Y(n_1840)
);

AO21x2_ASAP7_75t_L g1841 ( 
.A1(n_1839),
.A2(n_1699),
.B(n_1697),
.Y(n_1841)
);

AOI21x1_ASAP7_75t_L g1842 ( 
.A1(n_1841),
.A2(n_1840),
.B(n_1690),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1842),
.Y(n_1843)
);

OAI221xp5_ASAP7_75t_R g1844 ( 
.A1(n_1843),
.A2(n_1703),
.B1(n_1631),
.B2(n_1691),
.C(n_1679),
.Y(n_1844)
);

AOI211xp5_ASAP7_75t_L g1845 ( 
.A1(n_1844),
.A2(n_1553),
.B(n_1550),
.C(n_1556),
.Y(n_1845)
);


endmodule