module fake_netlist_6_2212_n_1839 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_186, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1839);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_186;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1839;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_220;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_153),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_14),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_81),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_78),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_60),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_124),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_9),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_80),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_138),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_36),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_62),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_118),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_87),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_169),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_182),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_108),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_82),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_50),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_143),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_21),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_46),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_54),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_181),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_25),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_51),
.Y(n_214)
);

INVxp33_ASAP7_75t_SL g215 ( 
.A(n_93),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_111),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_21),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_103),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_163),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_129),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_9),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_86),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_7),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_32),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_171),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_183),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_123),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_148),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_116),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_37),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_135),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_133),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_2),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_184),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_50),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_79),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_150),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_22),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_71),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_130),
.Y(n_240)
);

INVxp67_ASAP7_75t_SL g241 ( 
.A(n_134),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_69),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_25),
.Y(n_243)
);

BUFx8_ASAP7_75t_SL g244 ( 
.A(n_65),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_0),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_185),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_168),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_106),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_152),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_114),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_63),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_156),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_46),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_120),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_84),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_75),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_110),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_2),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_101),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_146),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_104),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_77),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_42),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_141),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_186),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_19),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_162),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_149),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_44),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_24),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_1),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_147),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_14),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_157),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_85),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_100),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_139),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_30),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_30),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_128),
.Y(n_280)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_24),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_26),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_45),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_7),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_57),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_136),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_131),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_119),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_54),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_55),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_12),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_59),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_127),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_98),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_91),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_41),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_115),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_83),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_137),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_27),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_92),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_160),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_97),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_10),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_172),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_170),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_52),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_112),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_32),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_37),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_105),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_74),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_154),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_11),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_96),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_177),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_113),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_45),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_176),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_39),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_88),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_47),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_70),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_26),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_73),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_57),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_175),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_13),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_20),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_58),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_180),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_52),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_42),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_20),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_17),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_28),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_11),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_27),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_166),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_34),
.Y(n_340)
);

CKINVDCx11_ASAP7_75t_R g341 ( 
.A(n_95),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_6),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_36),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_94),
.Y(n_344)
);

BUFx10_ASAP7_75t_L g345 ( 
.A(n_125),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_12),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_126),
.Y(n_347)
);

BUFx10_ASAP7_75t_L g348 ( 
.A(n_107),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_158),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_13),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_89),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_4),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_173),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_17),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_23),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_102),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_6),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_38),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_72),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_31),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_76),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_15),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_38),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_151),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_142),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_159),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_39),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_122),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_99),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_178),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_5),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_121),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_15),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_187),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_10),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_144),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_23),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_281),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_281),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_281),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_268),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_281),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_308),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_262),
.Y(n_384)
);

INVxp33_ASAP7_75t_L g385 ( 
.A(n_230),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_296),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_233),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_281),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_351),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_281),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_281),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_235),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_373),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_196),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_281),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_189),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_189),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_243),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_194),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_194),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_256),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_199),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_199),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_286),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_209),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_238),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_209),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_287),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_293),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_368),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_211),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_288),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_271),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_221),
.Y(n_414)
);

BUFx2_ASAP7_75t_SL g415 ( 
.A(n_198),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_245),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_265),
.Y(n_417)
);

INVxp33_ASAP7_75t_SL g418 ( 
.A(n_196),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_258),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_266),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_273),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_265),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_271),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_369),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_331),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g426 ( 
.A(n_331),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_244),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_286),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_339),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_278),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_339),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_207),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_283),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_286),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_284),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_289),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_284),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_341),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_317),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_300),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_234),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_263),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_269),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_240),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_364),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_242),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_304),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_246),
.Y(n_448)
);

CKINVDCx14_ASAP7_75t_R g449 ( 
.A(n_190),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_270),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_247),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_282),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_207),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_304),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_364),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_218),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_290),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_291),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_309),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_292),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_375),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_213),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_320),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_326),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_328),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_330),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_334),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_213),
.Y(n_468)
);

INVxp33_ASAP7_75t_SL g469 ( 
.A(n_217),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_350),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_375),
.Y(n_471)
);

BUFx5_ASAP7_75t_L g472 ( 
.A(n_192),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_249),
.Y(n_473)
);

BUFx2_ASAP7_75t_SL g474 ( 
.A(n_198),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_354),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_355),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_357),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_362),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_363),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_214),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_394),
.B(n_432),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_386),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_413),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_387),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_404),
.Y(n_485)
);

OAI21x1_ASAP7_75t_L g486 ( 
.A1(n_390),
.A2(n_218),
.B(n_226),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_386),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_390),
.A2(n_218),
.B(n_226),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_381),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_413),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_404),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_393),
.A2(n_343),
.B1(n_279),
.B2(n_253),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_404),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_423),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_404),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_423),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_404),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_417),
.B(n_214),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_435),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_415),
.B(n_215),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_387),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_428),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_427),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_425),
.B(n_251),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_435),
.Y(n_505)
);

NOR2x1_ASAP7_75t_L g506 ( 
.A(n_415),
.B(n_239),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_441),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_444),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_428),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_392),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_461),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_428),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_461),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_428),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_471),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_471),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_456),
.B(n_251),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_428),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_392),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_434),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_434),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_385),
.A2(n_210),
.B1(n_377),
.B2(n_285),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_388),
.Y(n_523)
);

NOR2x1_ASAP7_75t_L g524 ( 
.A(n_474),
.B(n_239),
.Y(n_524)
);

NOR2x1_ASAP7_75t_L g525 ( 
.A(n_474),
.B(n_250),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_446),
.Y(n_526)
);

AOI22x1_ASAP7_75t_SL g527 ( 
.A1(n_383),
.A2(n_377),
.B1(n_285),
.B2(n_310),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_434),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_398),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_388),
.Y(n_530)
);

AND2x4_ASAP7_75t_SL g531 ( 
.A(n_438),
.B(n_448),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_422),
.B(n_223),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_434),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_398),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_412),
.B(n_190),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_391),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_389),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_425),
.B(n_366),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_434),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_425),
.B(n_366),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_391),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_426),
.B(n_223),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_451),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_395),
.B(n_250),
.Y(n_544)
);

OR2x6_ASAP7_75t_L g545 ( 
.A(n_414),
.B(n_307),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_429),
.B(n_307),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_395),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_378),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_379),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_442),
.Y(n_550)
);

AND2x2_ASAP7_75t_SL g551 ( 
.A(n_380),
.B(n_252),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_382),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_396),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_431),
.B(n_190),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_396),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_455),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_397),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_397),
.Y(n_558)
);

INVx6_ASAP7_75t_L g559 ( 
.A(n_472),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_445),
.B(n_455),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_472),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_424),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_560),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_498),
.B(n_384),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_523),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_549),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_523),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_485),
.Y(n_568)
);

INVxp67_ASAP7_75t_R g569 ( 
.A(n_484),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_517),
.B(n_472),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_530),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_530),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_536),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_498),
.B(n_401),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_560),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_507),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_485),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_549),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_500),
.B(n_418),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_541),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_556),
.Y(n_581)
);

AND2x6_ASAP7_75t_L g582 ( 
.A(n_517),
.B(n_252),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_549),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_541),
.Y(n_584)
);

AO21x2_ASAP7_75t_L g585 ( 
.A1(n_486),
.A2(n_201),
.B(n_197),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_547),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_551),
.A2(n_409),
.B1(n_410),
.B2(n_408),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_556),
.B(n_418),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_553),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_554),
.B(n_439),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_553),
.Y(n_591)
);

NAND2xp33_ASAP7_75t_L g592 ( 
.A(n_532),
.B(n_442),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_554),
.B(n_443),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_547),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_552),
.Y(n_595)
);

NOR2x1p5_ASAP7_75t_L g596 ( 
.A(n_481),
.B(n_217),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_517),
.B(n_472),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_556),
.B(n_469),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_552),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_544),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_551),
.B(n_532),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_508),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g603 ( 
.A1(n_545),
.A2(n_473),
.B1(n_449),
.B2(n_469),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_553),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_545),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_L g606 ( 
.A(n_542),
.B(n_443),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_553),
.Y(n_607)
);

CKINVDCx6p67_ASAP7_75t_R g608 ( 
.A(n_489),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_544),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_557),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_544),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_526),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_548),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_544),
.Y(n_614)
);

OR2x6_ASAP7_75t_L g615 ( 
.A(n_545),
.B(n_421),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_548),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_542),
.B(n_472),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_485),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_546),
.B(n_472),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_548),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_548),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_548),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_557),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_546),
.A2(n_264),
.B1(n_297),
.B2(n_453),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_557),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_557),
.Y(n_626)
);

AOI21x1_ASAP7_75t_L g627 ( 
.A1(n_504),
.A2(n_297),
.B(n_264),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_548),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_485),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_537),
.Y(n_630)
);

NAND3xp33_ASAP7_75t_L g631 ( 
.A(n_481),
.B(n_452),
.C(n_450),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_486),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_485),
.Y(n_633)
);

BUFx4f_ASAP7_75t_L g634 ( 
.A(n_557),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_488),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_488),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_555),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_558),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_506),
.Y(n_639)
);

OR2x6_ASAP7_75t_L g640 ( 
.A(n_545),
.B(n_478),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_485),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_555),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_558),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_558),
.Y(n_644)
);

AND2x2_ASAP7_75t_SL g645 ( 
.A(n_501),
.B(n_286),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_558),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_543),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_492),
.A2(n_224),
.B1(n_314),
.B2(n_310),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_504),
.B(n_399),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_558),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_538),
.B(n_399),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_524),
.B(n_472),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_524),
.B(n_450),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_558),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_495),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_491),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_562),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_525),
.B(n_452),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_495),
.Y(n_659)
);

AND2x2_ASAP7_75t_SL g660 ( 
.A(n_501),
.B(n_286),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_483),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_535),
.B(n_457),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_559),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_525),
.B(n_457),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_495),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_545),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_559),
.Y(n_667)
);

OR2x6_ASAP7_75t_L g668 ( 
.A(n_538),
.B(n_540),
.Y(n_668)
);

AO22x2_ASAP7_75t_L g669 ( 
.A1(n_492),
.A2(n_406),
.B1(n_227),
.B2(n_202),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_497),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_540),
.B(n_458),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_490),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_491),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_490),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_497),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_497),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_491),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_529),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_494),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_539),
.B(n_458),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_509),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_494),
.A2(n_462),
.B1(n_468),
.B2(n_215),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_R g683 ( 
.A(n_510),
.B(n_460),
.Y(n_683)
);

INVx5_ASAP7_75t_L g684 ( 
.A(n_559),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_509),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_491),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_539),
.B(n_460),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_496),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_559),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_491),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_496),
.A2(n_419),
.B1(n_430),
.B2(n_477),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_509),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_534),
.B(n_550),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_510),
.B(n_479),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_493),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_493),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_493),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_519),
.B(n_193),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_519),
.B(n_193),
.Y(n_699)
);

BUFx8_ASAP7_75t_SL g700 ( 
.A(n_503),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_499),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_512),
.B(n_225),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_512),
.Y(n_703)
);

BUFx4f_ASAP7_75t_L g704 ( 
.A(n_493),
.Y(n_704)
);

BUFx6f_ASAP7_75t_SL g705 ( 
.A(n_499),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_630),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_R g707 ( 
.A(n_576),
.B(n_482),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_645),
.A2(n_660),
.B1(n_579),
.B2(n_639),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_694),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_671),
.B(n_482),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_645),
.A2(n_216),
.B1(n_229),
.B2(n_228),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_566),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_563),
.B(n_487),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_645),
.B(n_660),
.Y(n_714)
);

BUFx4f_ASAP7_75t_L g715 ( 
.A(n_660),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_566),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_581),
.B(n_411),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_600),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_609),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_601),
.B(n_561),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_563),
.B(n_512),
.Y(n_721)
);

NOR2x1p5_ASAP7_75t_L g722 ( 
.A(n_608),
.B(n_224),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_575),
.B(n_514),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_653),
.B(n_658),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_611),
.Y(n_725)
);

NOR2xp67_ASAP7_75t_L g726 ( 
.A(n_631),
.B(n_522),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_565),
.B(n_514),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_565),
.B(n_518),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_567),
.B(n_518),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_567),
.B(n_518),
.Y(n_730)
);

OR2x6_ASAP7_75t_L g731 ( 
.A(n_605),
.B(n_487),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_680),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_592),
.A2(n_241),
.B1(n_294),
.B2(n_374),
.Y(n_733)
);

BUFx8_ASAP7_75t_L g734 ( 
.A(n_705),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_617),
.B(n_232),
.Y(n_735)
);

OAI221xp5_ASAP7_75t_L g736 ( 
.A1(n_624),
.A2(n_299),
.B1(n_260),
.B2(n_522),
.C(n_416),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_581),
.B(n_420),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_578),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_611),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_582),
.A2(n_302),
.B1(n_303),
.B2(n_353),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_668),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_687),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_664),
.B(n_188),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_618),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_571),
.B(n_572),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_583),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_587),
.A2(n_301),
.B1(n_327),
.B2(n_323),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_606),
.A2(n_295),
.B1(n_254),
.B2(n_259),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_574),
.B(n_188),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_572),
.B(n_520),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_583),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_573),
.B(n_520),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_573),
.B(n_521),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_614),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_SL g755 ( 
.A(n_576),
.B(n_531),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_661),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_580),
.B(n_533),
.Y(n_757)
);

INVx5_ASAP7_75t_L g758 ( 
.A(n_582),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_619),
.B(n_236),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_618),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_580),
.B(n_533),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_637),
.B(n_433),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_570),
.B(n_237),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_593),
.B(n_191),
.Y(n_764)
);

NOR2xp67_ASAP7_75t_L g765 ( 
.A(n_662),
.B(n_505),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_584),
.B(n_533),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_642),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_584),
.B(n_559),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_586),
.B(n_255),
.Y(n_769)
);

O2A1O1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_586),
.A2(n_466),
.B(n_436),
.C(n_440),
.Y(n_770)
);

OR2x6_ASAP7_75t_L g771 ( 
.A(n_605),
.B(n_480),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_594),
.B(n_257),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_564),
.B(n_191),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_594),
.B(n_261),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_564),
.B(n_531),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_595),
.B(n_267),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_595),
.B(n_272),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_599),
.B(n_275),
.Y(n_778)
);

OR2x2_ASAP7_75t_L g779 ( 
.A(n_682),
.B(n_531),
.Y(n_779)
);

NAND2xp33_ASAP7_75t_SL g780 ( 
.A(n_596),
.B(n_314),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_599),
.B(n_668),
.Y(n_781)
);

BUFx6f_ASAP7_75t_SL g782 ( 
.A(n_615),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_668),
.B(n_321),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_649),
.B(n_651),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_615),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_651),
.B(n_597),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_672),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_674),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_588),
.B(n_195),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_582),
.B(n_511),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_666),
.B(n_679),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_582),
.B(n_513),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_679),
.Y(n_793)
);

OR2x4_ASAP7_75t_L g794 ( 
.A(n_598),
.B(n_480),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_702),
.B(n_513),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_688),
.B(n_515),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_701),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_652),
.B(n_274),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_701),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_655),
.Y(n_800)
);

NAND2xp33_ASAP7_75t_L g801 ( 
.A(n_632),
.B(n_276),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_663),
.B(n_515),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_663),
.B(n_516),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_590),
.A2(n_277),
.B1(n_344),
.B2(n_347),
.Y(n_804)
);

INVxp67_ASAP7_75t_L g805 ( 
.A(n_693),
.Y(n_805)
);

NAND2x1p5_ASAP7_75t_L g806 ( 
.A(n_667),
.B(n_516),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_678),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_659),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_666),
.A2(n_699),
.B1(n_698),
.B2(n_705),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_684),
.B(n_298),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_667),
.B(n_493),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_689),
.B(n_616),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_659),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_689),
.B(n_493),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_665),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_620),
.B(n_621),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_620),
.B(n_502),
.Y(n_817)
);

NAND3xp33_ASAP7_75t_L g818 ( 
.A(n_683),
.B(n_346),
.C(n_360),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_665),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_615),
.B(n_459),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_670),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_618),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_621),
.B(n_622),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_670),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_615),
.B(n_195),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_675),
.Y(n_826)
);

AND2x2_ASAP7_75t_SL g827 ( 
.A(n_648),
.B(n_463),
.Y(n_827)
);

INVx8_ASAP7_75t_L g828 ( 
.A(n_705),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_640),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_675),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_640),
.A2(n_349),
.B1(n_305),
.B2(n_356),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_676),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_640),
.B(n_200),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_640),
.B(n_603),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_569),
.B(n_464),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_648),
.B(n_200),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_632),
.B(n_465),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_676),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_622),
.B(n_502),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_628),
.B(n_203),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_681),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_635),
.A2(n_212),
.B1(n_203),
.B2(n_205),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_700),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_643),
.B(n_502),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_643),
.B(n_502),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_706),
.Y(n_846)
);

BUFx4f_ASAP7_75t_L g847 ( 
.A(n_828),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_718),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_744),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_807),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_843),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_724),
.B(n_784),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_741),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_719),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_744),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_707),
.Y(n_856)
);

INVx4_ASAP7_75t_L g857 ( 
.A(n_828),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_725),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_709),
.B(n_657),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_708),
.B(n_709),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_732),
.B(n_568),
.Y(n_861)
);

OR2x2_ASAP7_75t_SL g862 ( 
.A(n_779),
.B(n_527),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_775),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_791),
.B(n_467),
.Y(n_864)
);

NOR3xp33_ASAP7_75t_SL g865 ( 
.A(n_836),
.B(n_322),
.C(n_318),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_741),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_791),
.B(n_470),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_742),
.B(n_568),
.Y(n_868)
);

BUFx4f_ASAP7_75t_L g869 ( 
.A(n_828),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_739),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_711),
.A2(n_669),
.B1(n_636),
.B2(n_585),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_754),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_707),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_805),
.B(n_602),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_711),
.A2(n_669),
.B1(n_585),
.B2(n_371),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_794),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_789),
.B(n_786),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_756),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_805),
.B(n_602),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_788),
.Y(n_880)
);

INVxp67_ASAP7_75t_L g881 ( 
.A(n_713),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_714),
.A2(n_569),
.B1(n_646),
.B2(n_669),
.Y(n_882)
);

INVx5_ASAP7_75t_L g883 ( 
.A(n_758),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_715),
.A2(n_669),
.B1(n_612),
.B2(n_647),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_734),
.Y(n_885)
);

NOR2x1_ASAP7_75t_R g886 ( 
.A(n_820),
.B(n_647),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_744),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_710),
.B(n_527),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_710),
.B(n_713),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_794),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_743),
.B(n_577),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_743),
.B(n_577),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_714),
.B(n_629),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_787),
.Y(n_894)
);

INVx3_ASAP7_75t_L g895 ( 
.A(n_837),
.Y(n_895)
);

NOR2x2_ASAP7_75t_L g896 ( 
.A(n_731),
.B(n_608),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_820),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_773),
.B(n_629),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_773),
.B(n_629),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_793),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_835),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_781),
.B(n_684),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_782),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_749),
.B(n_691),
.Y(n_904)
);

INVx6_ASAP7_75t_L g905 ( 
.A(n_717),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_SL g906 ( 
.A1(n_834),
.A2(n_324),
.B1(n_318),
.B2(n_322),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_765),
.B(n_684),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_797),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_799),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_771),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_767),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_749),
.B(n_633),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_782),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_721),
.Y(n_914)
);

NOR3xp33_ASAP7_75t_SL g915 ( 
.A(n_780),
.B(n_329),
.C(n_324),
.Y(n_915)
);

NOR3xp33_ASAP7_75t_SL g916 ( 
.A(n_736),
.B(n_332),
.C(n_329),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_771),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_745),
.B(n_641),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_795),
.B(n_641),
.Y(n_919)
);

BUFx4f_ASAP7_75t_L g920 ( 
.A(n_731),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_837),
.B(n_641),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_744),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_764),
.B(n_613),
.Y(n_923)
);

INVx4_ASAP7_75t_L g924 ( 
.A(n_760),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_764),
.B(n_613),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_760),
.Y(n_926)
);

INVxp67_ASAP7_75t_L g927 ( 
.A(n_717),
.Y(n_927)
);

BUFx2_ASAP7_75t_L g928 ( 
.A(n_731),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_737),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_827),
.A2(n_585),
.B1(n_367),
.B2(n_332),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_762),
.B(n_475),
.Y(n_931)
);

OR2x4_ASAP7_75t_L g932 ( 
.A(n_825),
.B(n_476),
.Y(n_932)
);

NOR2x2_ASAP7_75t_L g933 ( 
.A(n_771),
.B(n_681),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_762),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_838),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_720),
.A2(n_634),
.B(n_704),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_827),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_809),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_723),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_726),
.A2(n_646),
.B1(n_638),
.B2(n_589),
.Y(n_940)
);

INVx4_ASAP7_75t_L g941 ( 
.A(n_760),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_760),
.Y(n_942)
);

NOR3xp33_ASAP7_75t_SL g943 ( 
.A(n_818),
.B(n_367),
.C(n_333),
.Y(n_943)
);

INVx2_ASAP7_75t_SL g944 ( 
.A(n_785),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_800),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_840),
.B(n_673),
.Y(n_946)
);

NAND3xp33_ASAP7_75t_SL g947 ( 
.A(n_733),
.B(n_205),
.C(n_204),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_840),
.B(n_677),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_783),
.Y(n_949)
);

INVx4_ASAP7_75t_L g950 ( 
.A(n_822),
.Y(n_950)
);

AOI21x1_ASAP7_75t_L g951 ( 
.A1(n_811),
.A2(n_627),
.B(n_607),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_808),
.Y(n_952)
);

OAI22xp33_ASAP7_75t_L g953 ( 
.A1(n_755),
.A2(n_333),
.B1(n_371),
.B2(n_336),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_740),
.A2(n_685),
.B1(n_703),
.B2(n_692),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_785),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_776),
.B(n_677),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_777),
.B(n_677),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_747),
.A2(n_280),
.B1(n_306),
.B2(n_248),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_822),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_829),
.B(n_589),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_834),
.B(n_613),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_842),
.B(n_335),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_819),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_727),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_821),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_829),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_825),
.B(n_833),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_SL g968 ( 
.A(n_833),
.B(n_338),
.C(n_337),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_778),
.B(n_340),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_826),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_769),
.B(n_772),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_796),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_831),
.B(n_342),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_832),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_748),
.B(n_804),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_728),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_822),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_722),
.B(n_812),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_L g979 ( 
.A1(n_740),
.A2(n_193),
.B1(n_248),
.B2(n_280),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_774),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_735),
.B(n_686),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_735),
.B(n_686),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_759),
.B(n_686),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_798),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_729),
.Y(n_985)
);

BUFx4f_ASAP7_75t_L g986 ( 
.A(n_806),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_816),
.B(n_591),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_759),
.B(n_690),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_730),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_823),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_841),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_790),
.A2(n_685),
.B1(n_604),
.B2(n_654),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_798),
.A2(n_763),
.B1(n_801),
.B2(n_792),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_806),
.Y(n_994)
);

AND3x2_ASAP7_75t_SL g995 ( 
.A(n_712),
.B(n_248),
.C(n_280),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_716),
.B(n_690),
.Y(n_996)
);

INVx1_ASAP7_75t_SL g997 ( 
.A(n_763),
.Y(n_997)
);

BUFx4f_ASAP7_75t_L g998 ( 
.A(n_813),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_750),
.Y(n_999)
);

INVxp67_ASAP7_75t_L g1000 ( 
.A(n_752),
.Y(n_1000)
);

INVxp67_ASAP7_75t_L g1001 ( 
.A(n_753),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_738),
.B(n_697),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_746),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_849),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_852),
.A2(n_761),
.B1(n_766),
.B2(n_757),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_849),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_889),
.A2(n_770),
.B(n_803),
.C(n_802),
.Y(n_1007)
);

BUFx12f_ASAP7_75t_L g1008 ( 
.A(n_885),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_877),
.B(n_751),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_914),
.B(n_939),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_883),
.A2(n_704),
.B(n_768),
.Y(n_1011)
);

OAI21xp33_ASAP7_75t_L g1012 ( 
.A1(n_962),
.A2(n_352),
.B(n_358),
.Y(n_1012)
);

INVx6_ASAP7_75t_L g1013 ( 
.A(n_846),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_858),
.Y(n_1014)
);

AND2x4_ASAP7_75t_SL g1015 ( 
.A(n_857),
.B(n_815),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_881),
.B(n_810),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_SL g1017 ( 
.A1(n_923),
.A2(n_626),
.B(n_610),
.C(n_623),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_881),
.B(n_810),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_870),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_883),
.A2(n_704),
.B(n_814),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_849),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_853),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_875),
.A2(n_824),
.B1(n_830),
.B2(n_845),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_990),
.B(n_964),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_971),
.A2(n_839),
.B(n_817),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_872),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_SL g1027 ( 
.A1(n_975),
.A2(n_844),
.B(n_650),
.C(n_644),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_904),
.B(n_400),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_863),
.B(n_901),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_951),
.A2(n_610),
.B(n_625),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_972),
.B(n_625),
.Y(n_1031)
);

NAND3xp33_ASAP7_75t_SL g1032 ( 
.A(n_967),
.B(n_313),
.C(n_312),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_873),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_936),
.A2(n_695),
.B(n_656),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_949),
.B(n_206),
.Y(n_1035)
);

NAND3xp33_ASAP7_75t_L g1036 ( 
.A(n_962),
.B(n_206),
.C(n_208),
.Y(n_1036)
);

BUFx4f_ASAP7_75t_L g1037 ( 
.A(n_978),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_1003),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_856),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_849),
.Y(n_1040)
);

OAI21xp33_ASAP7_75t_L g1041 ( 
.A1(n_967),
.A2(n_208),
.B(n_212),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_976),
.B(n_618),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_1003),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_848),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_985),
.B(n_656),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_875),
.A2(n_365),
.B1(n_220),
.B2(n_222),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_860),
.B(n_400),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_859),
.B(n_219),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_855),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_935),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_854),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_945),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_984),
.A2(n_359),
.B1(n_361),
.B2(n_219),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_947),
.A2(n_306),
.B1(n_345),
.B2(n_348),
.Y(n_1054)
);

OR2x6_ASAP7_75t_L g1055 ( 
.A(n_857),
.B(n_402),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_992),
.A2(n_437),
.B(n_403),
.Y(n_1056)
);

BUFx8_ASAP7_75t_L g1057 ( 
.A(n_928),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_961),
.A2(n_365),
.B1(n_222),
.B2(n_231),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_989),
.B(n_656),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_952),
.Y(n_1060)
);

OR2x2_ASAP7_75t_L g1061 ( 
.A(n_859),
.B(n_937),
.Y(n_1061)
);

OAI221xp5_ASAP7_75t_L g1062 ( 
.A1(n_958),
.A2(n_220),
.B1(n_231),
.B2(n_312),
.C(n_313),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_999),
.B(n_696),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_871),
.A2(n_376),
.B1(n_311),
.B2(n_315),
.Y(n_1064)
);

INVxp67_ASAP7_75t_L g1065 ( 
.A(n_966),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_923),
.A2(n_696),
.B(n_528),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_874),
.B(n_402),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_853),
.Y(n_1068)
);

O2A1O1Ixp5_ASAP7_75t_SL g1069 ( 
.A1(n_884),
.A2(n_454),
.B(n_447),
.C(n_407),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_917),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_949),
.B(n_696),
.Y(n_1071)
);

INVx4_ASAP7_75t_L g1072 ( 
.A(n_855),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_925),
.A2(n_528),
.B(n_370),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_SL g1074 ( 
.A1(n_893),
.A2(n_454),
.B(n_407),
.C(n_405),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_963),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_851),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_855),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_SL g1078 ( 
.A1(n_888),
.A2(n_306),
.B1(n_348),
.B2(n_345),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1000),
.B(n_325),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_925),
.A2(n_528),
.B(n_325),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_965),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_903),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_891),
.A2(n_528),
.B(n_376),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_916),
.A2(n_927),
.B(n_929),
.C(n_953),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1000),
.B(n_372),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_855),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_913),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_961),
.A2(n_316),
.B(n_372),
.C(n_370),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_850),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_887),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_SL g1091 ( 
.A1(n_969),
.A2(n_403),
.B(n_348),
.C(n_345),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_871),
.A2(n_319),
.B1(n_316),
.B2(n_3),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_892),
.A2(n_528),
.B(n_179),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_970),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_974),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_916),
.A2(n_0),
.B(n_1),
.C(n_3),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_991),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1001),
.B(n_174),
.Y(n_1098)
);

NOR3xp33_ASAP7_75t_L g1099 ( 
.A(n_879),
.B(n_4),
.C(n_5),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_866),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1001),
.B(n_167),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_898),
.A2(n_164),
.B(n_161),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_880),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_899),
.A2(n_155),
.B(n_145),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_879),
.B(n_8),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_912),
.B(n_140),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_911),
.B(n_980),
.Y(n_1107)
);

O2A1O1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_953),
.A2(n_8),
.B(n_16),
.C(n_18),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_895),
.B(n_132),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_878),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_979),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_987),
.B(n_109),
.Y(n_1112)
);

BUFx4f_ASAP7_75t_L g1113 ( 
.A(n_978),
.Y(n_1113)
);

INVx1_ASAP7_75t_SL g1114 ( 
.A(n_866),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_955),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_987),
.B(n_90),
.Y(n_1116)
);

NAND2x2_ASAP7_75t_L g1117 ( 
.A(n_910),
.B(n_22),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_876),
.A2(n_68),
.B1(n_67),
.B2(n_66),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_938),
.B(n_64),
.Y(n_1119)
);

AO21x1_ASAP7_75t_L g1120 ( 
.A1(n_993),
.A2(n_28),
.B(n_29),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_890),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_918),
.B(n_61),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_979),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_969),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_905),
.A2(n_60),
.B1(n_40),
.B2(n_41),
.Y(n_1125)
);

INVx4_ASAP7_75t_L g1126 ( 
.A(n_887),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_997),
.B(n_35),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_998),
.B(n_934),
.Y(n_1128)
);

AOI21x1_ASAP7_75t_L g1129 ( 
.A1(n_902),
.A2(n_40),
.B(n_43),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_909),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_894),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_R g1132 ( 
.A(n_847),
.B(n_59),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_998),
.B(n_47),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_931),
.B(n_48),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_SL g1135 ( 
.A(n_847),
.B(n_48),
.Y(n_1135)
);

BUFx8_ASAP7_75t_L g1136 ( 
.A(n_1008),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1007),
.A2(n_882),
.B(n_940),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1025),
.A2(n_946),
.B(n_948),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1106),
.A2(n_986),
.B(n_957),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1061),
.B(n_920),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_1029),
.B(n_920),
.Y(n_1141)
);

INVxp67_ASAP7_75t_SL g1142 ( 
.A(n_1022),
.Y(n_1142)
);

CKINVDCx16_ASAP7_75t_R g1143 ( 
.A(n_1115),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1024),
.B(n_944),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1051),
.Y(n_1145)
);

NOR2xp67_ASAP7_75t_L g1146 ( 
.A(n_1047),
.B(n_994),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1016),
.A2(n_1018),
.B(n_1069),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1106),
.A2(n_986),
.B(n_956),
.Y(n_1148)
);

NAND2x1p5_ASAP7_75t_L g1149 ( 
.A(n_1089),
.B(n_869),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1048),
.B(n_932),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1005),
.A2(n_907),
.B(n_919),
.Y(n_1151)
);

AO32x2_ASAP7_75t_L g1152 ( 
.A1(n_1092),
.A2(n_906),
.A3(n_954),
.B1(n_941),
.B2(n_924),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1005),
.A2(n_1066),
.B(n_1122),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1024),
.B(n_905),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1010),
.B(n_932),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1010),
.B(n_930),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1067),
.B(n_930),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1028),
.B(n_864),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_1039),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1134),
.B(n_867),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1033),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1009),
.B(n_864),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1020),
.A2(n_1002),
.B(n_996),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_1076),
.Y(n_1164)
);

NAND3xp33_ASAP7_75t_L g1165 ( 
.A(n_1078),
.B(n_958),
.C(n_865),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1107),
.B(n_867),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1084),
.A2(n_865),
.B(n_968),
.C(n_973),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1011),
.A2(n_1093),
.B(n_1122),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_1013),
.Y(n_1169)
);

AOI221x1_ASAP7_75t_L g1170 ( 
.A1(n_1092),
.A2(n_982),
.B1(n_988),
.B2(n_983),
.C(n_981),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_1072),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1009),
.B(n_960),
.Y(n_1172)
);

NOR2xp67_ASAP7_75t_L g1173 ( 
.A(n_1112),
.B(n_994),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_1004),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_1120),
.A2(n_921),
.A3(n_908),
.B(n_900),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_SL g1176 ( 
.A(n_1121),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1111),
.A2(n_943),
.B1(n_917),
.B2(n_968),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1105),
.B(n_960),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1079),
.B(n_966),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_1023),
.A2(n_868),
.A3(n_861),
.B(n_950),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_1036),
.A2(n_943),
.B(n_915),
.C(n_869),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1079),
.B(n_897),
.Y(n_1182)
);

NAND3x1_ASAP7_75t_L g1183 ( 
.A(n_1099),
.B(n_896),
.C(n_995),
.Y(n_1183)
);

AO21x2_ASAP7_75t_L g1184 ( 
.A1(n_1017),
.A2(n_915),
.B(n_995),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1085),
.B(n_977),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_1004),
.Y(n_1186)
);

INVx1_ASAP7_75t_SL g1187 ( 
.A(n_1114),
.Y(n_1187)
);

INVx3_ASAP7_75t_L g1188 ( 
.A(n_1072),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1116),
.A2(n_977),
.B(n_942),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1098),
.A2(n_942),
.B(n_950),
.Y(n_1190)
);

AND2x6_ASAP7_75t_L g1191 ( 
.A(n_1077),
.B(n_959),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1023),
.A2(n_1063),
.B(n_1042),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_1077),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1068),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1098),
.A2(n_933),
.B(n_862),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1111),
.A2(n_959),
.B1(n_926),
.B2(n_922),
.Y(n_1196)
);

OR2x2_ASAP7_75t_L g1197 ( 
.A(n_1085),
.B(n_926),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1103),
.B(n_886),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_1083),
.A2(n_926),
.A3(n_922),
.B(n_887),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_SL g1200 ( 
.A1(n_1101),
.A2(n_887),
.B(n_922),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1130),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1045),
.A2(n_922),
.B(n_51),
.Y(n_1202)
);

NAND3xp33_ASAP7_75t_SL g1203 ( 
.A(n_1054),
.B(n_49),
.C(n_53),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1027),
.A2(n_53),
.B(n_55),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1035),
.B(n_56),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1031),
.B(n_56),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1037),
.A2(n_1113),
.B1(n_1026),
.B2(n_1014),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1037),
.B(n_1113),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1114),
.B(n_1070),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1045),
.A2(n_1063),
.B(n_1059),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1019),
.B(n_1041),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1101),
.A2(n_1088),
.B(n_1073),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1110),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1123),
.A2(n_1135),
.B1(n_1127),
.B2(n_1133),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1059),
.A2(n_1129),
.B(n_1071),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1131),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1126),
.Y(n_1217)
);

OAI22x1_ASAP7_75t_L g1218 ( 
.A1(n_1125),
.A2(n_1119),
.B1(n_1100),
.B2(n_1065),
.Y(n_1218)
);

INVx4_ASAP7_75t_L g1219 ( 
.A(n_1013),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1080),
.A2(n_1071),
.B(n_1102),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_1053),
.B(n_1135),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_1124),
.A2(n_1123),
.A3(n_1104),
.B(n_1064),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1109),
.A2(n_1128),
.B(n_1015),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1052),
.A2(n_1075),
.B(n_1097),
.Y(n_1224)
);

INVx3_ASAP7_75t_SL g1225 ( 
.A(n_1082),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1012),
.B(n_1058),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1038),
.B(n_1043),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1057),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1032),
.A2(n_1062),
.B1(n_1046),
.B2(n_1064),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1060),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1081),
.A2(n_1095),
.B(n_1094),
.Y(n_1231)
);

INVx2_ASAP7_75t_SL g1232 ( 
.A(n_1057),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1050),
.B(n_1046),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1055),
.B(n_1087),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1055),
.B(n_1132),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1006),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1021),
.A2(n_1040),
.B(n_1049),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1086),
.B(n_1090),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1086),
.Y(n_1239)
);

BUFx12f_ASAP7_75t_L g1240 ( 
.A(n_1055),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1049),
.Y(n_1241)
);

INVx5_ASAP7_75t_L g1242 ( 
.A(n_1086),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1090),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1090),
.A2(n_1074),
.B(n_1091),
.Y(n_1244)
);

AO31x2_ASAP7_75t_L g1245 ( 
.A1(n_1096),
.A2(n_1108),
.A3(n_1117),
.B(n_1118),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1024),
.B(n_889),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1024),
.B(n_889),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1048),
.A2(n_889),
.B(n_967),
.C(n_852),
.Y(n_1248)
);

AOI221xp5_ASAP7_75t_L g1249 ( 
.A1(n_1092),
.A2(n_889),
.B1(n_888),
.B2(n_669),
.C(n_492),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1010),
.A2(n_889),
.B1(n_715),
.B2(n_708),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_SL g1251 ( 
.A1(n_1078),
.A2(n_889),
.B(n_967),
.Y(n_1251)
);

AOI21x1_ASAP7_75t_SL g1252 ( 
.A1(n_1106),
.A2(n_877),
.B(n_1105),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_1033),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1024),
.B(n_889),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1044),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1072),
.Y(n_1256)
);

A2O1A1Ixp33_ASAP7_75t_L g1257 ( 
.A1(n_1048),
.A2(n_889),
.B(n_967),
.C(n_852),
.Y(n_1257)
);

AO31x2_ASAP7_75t_L g1258 ( 
.A1(n_1120),
.A2(n_1092),
.A3(n_1023),
.B(n_1005),
.Y(n_1258)
);

AO32x2_ASAP7_75t_L g1259 ( 
.A1(n_1092),
.A2(n_1123),
.A3(n_1111),
.B1(n_1023),
.B2(n_1064),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1004),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1128),
.B(n_955),
.Y(n_1261)
);

AOI221x1_ASAP7_75t_L g1262 ( 
.A1(n_1092),
.A2(n_1099),
.B1(n_889),
.B2(n_967),
.C(n_1111),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1128),
.B(n_955),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1010),
.A2(n_889),
.B1(n_715),
.B2(n_708),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1010),
.A2(n_889),
.B1(n_715),
.B2(n_708),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1044),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1030),
.A2(n_1034),
.B(n_951),
.Y(n_1267)
);

NAND3xp33_ASAP7_75t_L g1268 ( 
.A(n_1048),
.B(n_889),
.C(n_789),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1120),
.A2(n_1092),
.A3(n_1023),
.B(n_1005),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1030),
.A2(n_1056),
.B(n_1106),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1024),
.B(n_889),
.Y(n_1271)
);

AOI21xp33_ASAP7_75t_SL g1272 ( 
.A1(n_1150),
.A2(n_1165),
.B(n_1155),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1267),
.A2(n_1163),
.B(n_1189),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1246),
.B(n_1271),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1268),
.A2(n_1257),
.B(n_1248),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1187),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1266),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1247),
.B(n_1254),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_SL g1279 ( 
.A(n_1219),
.B(n_1159),
.Y(n_1279)
);

AND2x4_ASAP7_75t_SL g1280 ( 
.A(n_1219),
.B(n_1164),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1153),
.A2(n_1137),
.B(n_1138),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1268),
.A2(n_1251),
.B1(n_1249),
.B2(n_1229),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1145),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_SL g1284 ( 
.A1(n_1165),
.A2(n_1157),
.B1(n_1156),
.B2(n_1265),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1160),
.B(n_1158),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1162),
.B(n_1179),
.Y(n_1286)
);

AOI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1244),
.A2(n_1148),
.B(n_1139),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1251),
.A2(n_1262),
.B(n_1229),
.Y(n_1288)
);

OA21x2_ASAP7_75t_L g1289 ( 
.A1(n_1168),
.A2(n_1192),
.B(n_1151),
.Y(n_1289)
);

A2O1A1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1214),
.A2(n_1264),
.B(n_1250),
.C(n_1167),
.Y(n_1290)
);

INVx6_ASAP7_75t_L g1291 ( 
.A(n_1242),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1220),
.A2(n_1204),
.A3(n_1210),
.B(n_1170),
.Y(n_1292)
);

AOI221xp5_ASAP7_75t_L g1293 ( 
.A1(n_1203),
.A2(n_1221),
.B1(n_1214),
.B2(n_1147),
.C(n_1218),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1154),
.B(n_1178),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1201),
.Y(n_1295)
);

O2A1O1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1226),
.A2(n_1205),
.B(n_1166),
.C(n_1181),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1215),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1177),
.A2(n_1195),
.B1(n_1212),
.B2(n_1233),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1213),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1161),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1194),
.B(n_1182),
.Y(n_1301)
);

CKINVDCx6p67_ASAP7_75t_R g1302 ( 
.A(n_1225),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1253),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1200),
.A2(n_1270),
.B(n_1190),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1169),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1216),
.Y(n_1306)
);

NAND2xp33_ASAP7_75t_L g1307 ( 
.A(n_1191),
.B(n_1172),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1136),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1230),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1236),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1149),
.Y(n_1311)
);

AO21x2_ASAP7_75t_L g1312 ( 
.A1(n_1173),
.A2(n_1196),
.B(n_1202),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1206),
.A2(n_1140),
.B1(n_1146),
.B2(n_1185),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1252),
.A2(n_1270),
.B(n_1237),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1180),
.Y(n_1315)
);

INVx1_ASAP7_75t_SL g1316 ( 
.A(n_1143),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1180),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1224),
.A2(n_1231),
.B(n_1223),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1196),
.A2(n_1211),
.B(n_1207),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1197),
.A2(n_1144),
.B(n_1183),
.Y(n_1320)
);

INVxp67_ASAP7_75t_L g1321 ( 
.A(n_1142),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1171),
.Y(n_1322)
);

INVx4_ASAP7_75t_L g1323 ( 
.A(n_1242),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1261),
.Y(n_1324)
);

BUFx2_ASAP7_75t_R g1325 ( 
.A(n_1208),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1238),
.A2(n_1141),
.B(n_1227),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1241),
.A2(n_1256),
.B(n_1217),
.Y(n_1327)
);

AOI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1243),
.A2(n_1239),
.B(n_1198),
.Y(n_1328)
);

INVxp67_ASAP7_75t_L g1329 ( 
.A(n_1176),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1188),
.A2(n_1217),
.B(n_1256),
.Y(n_1330)
);

AO32x2_ASAP7_75t_L g1331 ( 
.A1(n_1259),
.A2(n_1269),
.A3(n_1258),
.B1(n_1180),
.B2(n_1175),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1242),
.A2(n_1184),
.B(n_1259),
.Y(n_1332)
);

OA21x2_ASAP7_75t_L g1333 ( 
.A1(n_1258),
.A2(n_1269),
.B(n_1175),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1258),
.A2(n_1269),
.B(n_1222),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1184),
.A2(n_1259),
.B(n_1188),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1263),
.A2(n_1235),
.B1(n_1176),
.B2(n_1240),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1199),
.A2(n_1234),
.B(n_1222),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1174),
.Y(n_1338)
);

AO31x2_ASAP7_75t_L g1339 ( 
.A1(n_1222),
.A2(n_1152),
.A3(n_1199),
.B(n_1245),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1228),
.A2(n_1232),
.B1(n_1136),
.B2(n_1245),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1152),
.A2(n_1199),
.A3(n_1245),
.B(n_1191),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1152),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1186),
.B(n_1193),
.Y(n_1343)
);

A2O1A1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1193),
.A2(n_889),
.B(n_1257),
.C(n_1248),
.Y(n_1344)
);

NAND2x1_ASAP7_75t_L g1345 ( 
.A(n_1260),
.B(n_1200),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1260),
.A2(n_1267),
.B(n_1163),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1179),
.B(n_1162),
.Y(n_1347)
);

OR2x6_ASAP7_75t_L g1348 ( 
.A(n_1200),
.B(n_1208),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1267),
.A2(n_1163),
.B(n_1189),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1267),
.A2(n_1163),
.B(n_1189),
.Y(n_1350)
);

BUFx2_ASAP7_75t_SL g1351 ( 
.A(n_1164),
.Y(n_1351)
);

AOI21xp33_ASAP7_75t_L g1352 ( 
.A1(n_1268),
.A2(n_889),
.B(n_967),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_1209),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1267),
.A2(n_1163),
.B(n_1189),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1268),
.A2(n_889),
.B1(n_1257),
.B2(n_1248),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1267),
.A2(n_1163),
.B(n_1189),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1255),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1271),
.B(n_1246),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1242),
.Y(n_1359)
);

NAND2x1p5_ASAP7_75t_L g1360 ( 
.A(n_1208),
.B(n_1242),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1255),
.Y(n_1361)
);

O2A1O1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1251),
.A2(n_1257),
.B(n_1248),
.C(n_1268),
.Y(n_1362)
);

OAI221xp5_ASAP7_75t_L g1363 ( 
.A1(n_1249),
.A2(n_1078),
.B1(n_1251),
.B2(n_662),
.C(n_1268),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1255),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1267),
.A2(n_1163),
.B(n_1189),
.Y(n_1365)
);

INVx4_ASAP7_75t_SL g1366 ( 
.A(n_1191),
.Y(n_1366)
);

OA21x2_ASAP7_75t_L g1367 ( 
.A1(n_1153),
.A2(n_1137),
.B(n_1267),
.Y(n_1367)
);

BUFx2_ASAP7_75t_R g1368 ( 
.A(n_1159),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1138),
.A2(n_1153),
.B(n_1220),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1267),
.A2(n_1163),
.B(n_1189),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1219),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_1219),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1268),
.A2(n_1092),
.B1(n_889),
.B2(n_1111),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1209),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1251),
.B(n_1268),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1255),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_1219),
.Y(n_1377)
);

AOI21xp33_ASAP7_75t_L g1378 ( 
.A1(n_1268),
.A2(n_889),
.B(n_967),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1267),
.A2(n_1163),
.B(n_1189),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1208),
.B(n_1261),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1179),
.B(n_1162),
.Y(n_1381)
);

NAND3xp33_ASAP7_75t_L g1382 ( 
.A(n_1268),
.B(n_889),
.C(n_967),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1187),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1160),
.B(n_1158),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1268),
.A2(n_889),
.B(n_1248),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1187),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1268),
.A2(n_967),
.B1(n_1251),
.B2(n_383),
.Y(n_1387)
);

OR2x6_ASAP7_75t_L g1388 ( 
.A(n_1200),
.B(n_1208),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1208),
.B(n_1261),
.Y(n_1389)
);

AOI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1268),
.A2(n_967),
.B1(n_1251),
.B2(n_383),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1255),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1255),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1209),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1271),
.B(n_1246),
.Y(n_1394)
);

O2A1O1Ixp33_ASAP7_75t_SL g1395 ( 
.A1(n_1248),
.A2(n_1257),
.B(n_1124),
.C(n_714),
.Y(n_1395)
);

O2A1O1Ixp33_ASAP7_75t_L g1396 ( 
.A1(n_1251),
.A2(n_1257),
.B(n_1248),
.C(n_1268),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1209),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1179),
.B(n_1162),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1268),
.A2(n_889),
.B(n_1248),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1255),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1285),
.B(n_1384),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1363),
.A2(n_1387),
.B1(n_1390),
.B2(n_1373),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1300),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1286),
.B(n_1347),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1280),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1380),
.B(n_1389),
.Y(n_1406)
);

NOR2x1_ASAP7_75t_SL g1407 ( 
.A(n_1348),
.B(n_1388),
.Y(n_1407)
);

O2A1O1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1282),
.A2(n_1378),
.B(n_1352),
.C(n_1355),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1341),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1281),
.A2(n_1399),
.B(n_1385),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1397),
.B(n_1353),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1373),
.A2(n_1298),
.B1(n_1382),
.B2(n_1274),
.Y(n_1412)
);

O2A1O1Ixp5_ASAP7_75t_L g1413 ( 
.A1(n_1288),
.A2(n_1275),
.B(n_1375),
.C(n_1290),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1381),
.B(n_1398),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1278),
.B(n_1358),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_SL g1416 ( 
.A1(n_1296),
.A2(n_1344),
.B(n_1290),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1394),
.B(n_1294),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1324),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_1303),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1368),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1367),
.A2(n_1396),
.B(n_1362),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1301),
.B(n_1276),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1280),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1375),
.B(n_1284),
.Y(n_1424)
);

O2A1O1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1272),
.A2(n_1395),
.B(n_1344),
.C(n_1296),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1284),
.B(n_1276),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1383),
.B(n_1386),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1298),
.A2(n_1340),
.B1(n_1313),
.B2(n_1293),
.Y(n_1428)
);

O2A1O1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1293),
.A2(n_1320),
.B(n_1307),
.C(n_1321),
.Y(n_1429)
);

CKINVDCx16_ASAP7_75t_R g1430 ( 
.A(n_1279),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1305),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1383),
.B(n_1386),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1289),
.A2(n_1318),
.B(n_1319),
.Y(n_1433)
);

OA21x2_ASAP7_75t_L g1434 ( 
.A1(n_1314),
.A2(n_1332),
.B(n_1379),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1340),
.A2(n_1313),
.B1(n_1325),
.B2(n_1305),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1283),
.B(n_1299),
.Y(n_1436)
);

AOI221x1_ASAP7_75t_SL g1437 ( 
.A1(n_1336),
.A2(n_1295),
.B1(n_1392),
.B2(n_1277),
.C(n_1357),
.Y(n_1437)
);

AOI221x1_ASAP7_75t_SL g1438 ( 
.A1(n_1361),
.A2(n_1400),
.B1(n_1391),
.B2(n_1364),
.C(n_1376),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1311),
.B(n_1366),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1329),
.A2(n_1360),
.B1(n_1371),
.B2(n_1348),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_SL g1441 ( 
.A1(n_1359),
.A2(n_1388),
.B(n_1348),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1306),
.B(n_1309),
.Y(n_1442)
);

INVxp67_ASAP7_75t_L g1443 ( 
.A(n_1310),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1359),
.A2(n_1388),
.B(n_1323),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1316),
.B(n_1337),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1328),
.B(n_1326),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1332),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1326),
.B(n_1322),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_1335),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1329),
.A2(n_1360),
.B1(n_1371),
.B2(n_1377),
.Y(n_1450)
);

OAI22x1_ASAP7_75t_L g1451 ( 
.A1(n_1334),
.A2(n_1333),
.B1(n_1342),
.B2(n_1287),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1366),
.B(n_1338),
.Y(n_1452)
);

AOI221xp5_ASAP7_75t_L g1453 ( 
.A1(n_1335),
.A2(n_1342),
.B1(n_1351),
.B2(n_1372),
.C(n_1308),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1327),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1302),
.A2(n_1291),
.B1(n_1345),
.B2(n_1323),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1334),
.B(n_1339),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1339),
.B(n_1330),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1333),
.B(n_1312),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1315),
.A2(n_1317),
.B1(n_1297),
.B2(n_1333),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1292),
.B(n_1312),
.Y(n_1460)
);

INVx3_ASAP7_75t_L g1461 ( 
.A(n_1346),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_1331),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1273),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1349),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1350),
.A2(n_1370),
.B(n_1354),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1292),
.B(n_1356),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1365),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1285),
.B(n_1384),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1369),
.A2(n_1281),
.B(n_1153),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1280),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1374),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_1359),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_SL g1473 ( 
.A1(n_1296),
.A2(n_1257),
.B(n_1248),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1286),
.B(n_1347),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1286),
.B(n_1347),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1285),
.B(n_1384),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1304),
.A2(n_1153),
.B(n_1369),
.Y(n_1477)
);

AOI21xp5_ASAP7_75t_SL g1478 ( 
.A1(n_1296),
.A2(n_1257),
.B(n_1248),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1300),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1296),
.A2(n_1257),
.B(n_1248),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1374),
.B(n_1393),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1285),
.B(n_1384),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1285),
.B(n_1384),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1363),
.A2(n_1268),
.B1(n_1390),
.B2(n_1387),
.Y(n_1484)
);

O2A1O1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1363),
.A2(n_1251),
.B(n_1257),
.C(n_1248),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1286),
.B(n_1347),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1363),
.A2(n_1268),
.B1(n_1390),
.B2(n_1387),
.Y(n_1487)
);

OA22x2_ASAP7_75t_L g1488 ( 
.A1(n_1387),
.A2(n_1390),
.B1(n_1251),
.B2(n_1229),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1341),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1286),
.B(n_1347),
.Y(n_1490)
);

BUFx8_ASAP7_75t_L g1491 ( 
.A(n_1343),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1285),
.B(n_1384),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1374),
.B(n_1393),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_SL g1494 ( 
.A1(n_1296),
.A2(n_1257),
.B(n_1248),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1460),
.B(n_1447),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1451),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1457),
.B(n_1466),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1434),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1464),
.B(n_1454),
.Y(n_1499)
);

OAI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1408),
.A2(n_1485),
.B(n_1413),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1449),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1427),
.B(n_1404),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1461),
.B(n_1467),
.Y(n_1503)
);

BUFx4f_ASAP7_75t_SL g1504 ( 
.A(n_1419),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_1491),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1458),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1434),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1474),
.B(n_1475),
.Y(n_1508)
);

BUFx2_ASAP7_75t_L g1509 ( 
.A(n_1409),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1459),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1461),
.B(n_1463),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1446),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1402),
.A2(n_1488),
.B1(n_1484),
.B2(n_1487),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1446),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1433),
.A2(n_1469),
.B(n_1465),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1486),
.B(n_1490),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1489),
.B(n_1410),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1489),
.B(n_1410),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1421),
.B(n_1477),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_1432),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1443),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1443),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1456),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1445),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_SL g1525 ( 
.A1(n_1488),
.A2(n_1428),
.B1(n_1412),
.B2(n_1424),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1436),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1426),
.B(n_1422),
.Y(n_1527)
);

AO21x2_ASAP7_75t_L g1528 ( 
.A1(n_1473),
.A2(n_1494),
.B(n_1478),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1442),
.Y(n_1529)
);

AO21x2_ASAP7_75t_L g1530 ( 
.A1(n_1480),
.A2(n_1416),
.B(n_1408),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1448),
.Y(n_1531)
);

AO21x2_ASAP7_75t_L g1532 ( 
.A1(n_1485),
.A2(n_1425),
.B(n_1429),
.Y(n_1532)
);

AO21x2_ASAP7_75t_L g1533 ( 
.A1(n_1425),
.A2(n_1429),
.B(n_1407),
.Y(n_1533)
);

BUFx6f_ASAP7_75t_L g1534 ( 
.A(n_1406),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1491),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1414),
.B(n_1493),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1462),
.B(n_1413),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_SL g1538 ( 
.A(n_1500),
.B(n_1430),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1498),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1506),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1498),
.Y(n_1541)
);

BUFx2_ASAP7_75t_L g1542 ( 
.A(n_1511),
.Y(n_1542)
);

NOR2x1_ASAP7_75t_L g1543 ( 
.A(n_1528),
.B(n_1441),
.Y(n_1543)
);

NAND2x1_ASAP7_75t_L g1544 ( 
.A(n_1499),
.B(n_1444),
.Y(n_1544)
);

BUFx3_ASAP7_75t_L g1545 ( 
.A(n_1505),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1506),
.Y(n_1546)
);

NAND4xp25_ASAP7_75t_SL g1547 ( 
.A(n_1513),
.B(n_1453),
.C(n_1415),
.D(n_1417),
.Y(n_1547)
);

INVx3_ASAP7_75t_L g1548 ( 
.A(n_1511),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1512),
.B(n_1481),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1512),
.B(n_1438),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1513),
.A2(n_1435),
.B1(n_1406),
.B2(n_1471),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1497),
.B(n_1401),
.Y(n_1552)
);

INVxp67_ASAP7_75t_L g1553 ( 
.A(n_1514),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1517),
.B(n_1518),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1514),
.B(n_1453),
.Y(n_1555)
);

INVxp67_ASAP7_75t_L g1556 ( 
.A(n_1501),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1501),
.B(n_1437),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1509),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1507),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_1511),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1505),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1524),
.B(n_1411),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1525),
.A2(n_1492),
.B1(n_1468),
.B2(n_1483),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1517),
.B(n_1482),
.Y(n_1564)
);

BUFx3_ASAP7_75t_L g1565 ( 
.A(n_1505),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1525),
.A2(n_1431),
.B1(n_1440),
.B2(n_1418),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1518),
.B(n_1476),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1521),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1502),
.B(n_1450),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1558),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1539),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1545),
.B(n_1536),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1558),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1540),
.Y(n_1574)
);

AND2x2_ASAP7_75t_SL g1575 ( 
.A(n_1538),
.B(n_1537),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1540),
.B(n_1518),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1539),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1546),
.B(n_1524),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_R g1579 ( 
.A(n_1538),
.B(n_1420),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1549),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1547),
.A2(n_1530),
.B1(n_1528),
.B2(n_1532),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1546),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1541),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1545),
.B(n_1536),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1547),
.A2(n_1530),
.B1(n_1528),
.B2(n_1532),
.Y(n_1585)
);

AOI211xp5_ASAP7_75t_L g1586 ( 
.A1(n_1563),
.A2(n_1537),
.B(n_1530),
.C(n_1528),
.Y(n_1586)
);

NAND3xp33_ASAP7_75t_L g1587 ( 
.A(n_1550),
.B(n_1510),
.C(n_1496),
.Y(n_1587)
);

NAND3xp33_ASAP7_75t_SL g1588 ( 
.A(n_1566),
.B(n_1563),
.C(n_1557),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1548),
.Y(n_1589)
);

AOI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1557),
.A2(n_1530),
.B1(n_1510),
.B2(n_1532),
.C(n_1516),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_1545),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1569),
.B(n_1536),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1561),
.Y(n_1593)
);

OA222x2_ASAP7_75t_L g1594 ( 
.A1(n_1555),
.A2(n_1530),
.B1(n_1532),
.B2(n_1496),
.C1(n_1495),
.C2(n_1527),
.Y(n_1594)
);

OAI221xp5_ASAP7_75t_L g1595 ( 
.A1(n_1551),
.A2(n_1516),
.B1(n_1508),
.B2(n_1502),
.C(n_1527),
.Y(n_1595)
);

OAI321xp33_ASAP7_75t_L g1596 ( 
.A1(n_1555),
.A2(n_1519),
.A3(n_1495),
.B1(n_1524),
.B2(n_1531),
.C(n_1455),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1549),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1548),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1543),
.A2(n_1532),
.B1(n_1533),
.B2(n_1531),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1548),
.B(n_1503),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1548),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1554),
.B(n_1520),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1569),
.B(n_1520),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_R g1604 ( 
.A(n_1561),
.B(n_1403),
.Y(n_1604)
);

OAI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1543),
.A2(n_1508),
.B1(n_1527),
.B2(n_1423),
.C(n_1405),
.Y(n_1605)
);

NAND2x1p5_ASAP7_75t_SL g1606 ( 
.A(n_1554),
.B(n_1519),
.Y(n_1606)
);

AOI222xp33_ASAP7_75t_L g1607 ( 
.A1(n_1553),
.A2(n_1504),
.B1(n_1519),
.B2(n_1531),
.C1(n_1526),
.C2(n_1535),
.Y(n_1607)
);

AOI221xp5_ASAP7_75t_L g1608 ( 
.A1(n_1553),
.A2(n_1526),
.B1(n_1531),
.B2(n_1522),
.C(n_1521),
.Y(n_1608)
);

INVxp67_ASAP7_75t_L g1609 ( 
.A(n_1562),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1571),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1590),
.A2(n_1533),
.B(n_1544),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1574),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1574),
.Y(n_1613)
);

AND2x2_ASAP7_75t_SL g1614 ( 
.A(n_1575),
.B(n_1534),
.Y(n_1614)
);

INVx1_ASAP7_75t_SL g1615 ( 
.A(n_1604),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1582),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1606),
.B(n_1554),
.Y(n_1617)
);

INVxp67_ASAP7_75t_SL g1618 ( 
.A(n_1578),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1579),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1571),
.Y(n_1620)
);

INVx4_ASAP7_75t_SL g1621 ( 
.A(n_1591),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1582),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1600),
.B(n_1601),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1592),
.B(n_1564),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1578),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1570),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1581),
.A2(n_1533),
.B(n_1544),
.Y(n_1627)
);

BUFx2_ASAP7_75t_L g1628 ( 
.A(n_1606),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1570),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1600),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1573),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1573),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1600),
.B(n_1542),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1571),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1600),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1589),
.B(n_1560),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1577),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1577),
.Y(n_1638)
);

OR2x6_ASAP7_75t_L g1639 ( 
.A(n_1591),
.B(n_1561),
.Y(n_1639)
);

INVx2_ASAP7_75t_SL g1640 ( 
.A(n_1591),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1606),
.B(n_1562),
.Y(n_1641)
);

OA21x2_ASAP7_75t_L g1642 ( 
.A1(n_1599),
.A2(n_1515),
.B(n_1559),
.Y(n_1642)
);

BUFx2_ASAP7_75t_L g1643 ( 
.A(n_1575),
.Y(n_1643)
);

NAND3xp33_ASAP7_75t_L g1644 ( 
.A(n_1586),
.B(n_1556),
.C(n_1531),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1576),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1583),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1583),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1572),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1591),
.Y(n_1649)
);

NAND2xp33_ASAP7_75t_L g1650 ( 
.A(n_1619),
.B(n_1585),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1648),
.B(n_1587),
.Y(n_1651)
);

NOR2x1_ASAP7_75t_L g1652 ( 
.A(n_1644),
.B(n_1587),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1626),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1643),
.B(n_1594),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1643),
.B(n_1594),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1614),
.B(n_1575),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1624),
.B(n_1603),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1614),
.B(n_1589),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1618),
.B(n_1597),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_SL g1660 ( 
.A(n_1614),
.B(n_1586),
.Y(n_1660)
);

AOI33xp33_ASAP7_75t_L g1661 ( 
.A1(n_1615),
.A2(n_1608),
.A3(n_1580),
.B1(n_1568),
.B2(n_1529),
.B3(n_1567),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1626),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1625),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1631),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1640),
.B(n_1584),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1610),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1621),
.B(n_1589),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1631),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1649),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1632),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1621),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1621),
.B(n_1589),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1640),
.B(n_1609),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1632),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1621),
.B(n_1598),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1612),
.Y(n_1676)
);

INVx1_ASAP7_75t_SL g1677 ( 
.A(n_1621),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_SL g1678 ( 
.A1(n_1644),
.A2(n_1533),
.B1(n_1595),
.B2(n_1605),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1628),
.B(n_1598),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_1639),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1610),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1617),
.B(n_1576),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1628),
.B(n_1598),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1612),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1613),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1617),
.B(n_1602),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1613),
.Y(n_1687)
);

OAI31xp33_ASAP7_75t_L g1688 ( 
.A1(n_1611),
.A2(n_1593),
.A3(n_1565),
.B(n_1588),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1633),
.B(n_1598),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1649),
.B(n_1504),
.Y(n_1690)
);

OAI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1627),
.A2(n_1596),
.B(n_1607),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1616),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1641),
.B(n_1591),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1641),
.B(n_1564),
.Y(n_1694)
);

INVxp67_ASAP7_75t_L g1695 ( 
.A(n_1629),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1653),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1653),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1656),
.B(n_1649),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1656),
.B(n_1671),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1663),
.B(n_1616),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1662),
.Y(n_1701)
);

AOI322xp5_ASAP7_75t_L g1702 ( 
.A1(n_1652),
.A2(n_1660),
.A3(n_1650),
.B1(n_1678),
.B2(n_1654),
.C1(n_1655),
.C2(n_1651),
.Y(n_1702)
);

BUFx3_ASAP7_75t_L g1703 ( 
.A(n_1669),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1677),
.B(n_1680),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1667),
.B(n_1639),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1686),
.B(n_1622),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1661),
.B(n_1645),
.Y(n_1707)
);

INVx1_ASAP7_75t_SL g1708 ( 
.A(n_1669),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1695),
.B(n_1552),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1662),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1686),
.B(n_1622),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1664),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1664),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1690),
.B(n_1535),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1657),
.B(n_1552),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1667),
.B(n_1639),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1672),
.B(n_1639),
.Y(n_1717)
);

NOR2x1_ASAP7_75t_L g1718 ( 
.A(n_1654),
.B(n_1639),
.Y(n_1718)
);

INVxp33_ASAP7_75t_L g1719 ( 
.A(n_1688),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1672),
.B(n_1623),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1679),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1675),
.B(n_1630),
.Y(n_1722)
);

INVxp67_ASAP7_75t_L g1723 ( 
.A(n_1665),
.Y(n_1723)
);

INVx2_ASAP7_75t_SL g1724 ( 
.A(n_1675),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1659),
.B(n_1535),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1668),
.Y(n_1726)
);

NOR5xp2_ASAP7_75t_L g1727 ( 
.A(n_1691),
.B(n_1556),
.C(n_1523),
.D(n_1638),
.E(n_1637),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1673),
.B(n_1564),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1658),
.B(n_1689),
.Y(n_1729)
);

INVxp67_ASAP7_75t_SL g1730 ( 
.A(n_1693),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1668),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1670),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1720),
.B(n_1658),
.Y(n_1733)
);

INVx1_ASAP7_75t_SL g1734 ( 
.A(n_1708),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1721),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1713),
.Y(n_1736)
);

INVx1_ASAP7_75t_SL g1737 ( 
.A(n_1703),
.Y(n_1737)
);

BUFx3_ASAP7_75t_L g1738 ( 
.A(n_1703),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1723),
.B(n_1704),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1706),
.B(n_1682),
.Y(n_1740)
);

INVx1_ASAP7_75t_SL g1741 ( 
.A(n_1699),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1720),
.B(n_1679),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1706),
.B(n_1682),
.Y(n_1743)
);

INVxp67_ASAP7_75t_L g1744 ( 
.A(n_1718),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1732),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1699),
.B(n_1683),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1724),
.B(n_1670),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1714),
.B(n_1479),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1698),
.B(n_1683),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1732),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1696),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1704),
.B(n_1655),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1698),
.B(n_1705),
.Y(n_1753)
);

AOI21xp33_ASAP7_75t_L g1754 ( 
.A1(n_1719),
.A2(n_1676),
.B(n_1674),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1697),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1729),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1705),
.B(n_1689),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1711),
.B(n_1694),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1711),
.B(n_1674),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1744),
.A2(n_1719),
.B1(n_1741),
.B2(n_1752),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1735),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_SL g1762 ( 
.A1(n_1753),
.A2(n_1730),
.B1(n_1707),
.B2(n_1702),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1734),
.B(n_1725),
.Y(n_1763)
);

AOI21xp33_ASAP7_75t_L g1764 ( 
.A1(n_1737),
.A2(n_1724),
.B(n_1717),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1738),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1753),
.B(n_1721),
.Y(n_1766)
);

AOI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1754),
.A2(n_1717),
.B(n_1716),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1738),
.B(n_1709),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1756),
.Y(n_1769)
);

AOI31xp33_ASAP7_75t_L g1770 ( 
.A1(n_1739),
.A2(n_1716),
.A3(n_1717),
.B(n_1700),
.Y(n_1770)
);

AOI31xp33_ASAP7_75t_L g1771 ( 
.A1(n_1736),
.A2(n_1756),
.A3(n_1746),
.B(n_1748),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1745),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1738),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1745),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1736),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_SL g1776 ( 
.A(n_1746),
.B(n_1749),
.Y(n_1776)
);

NAND5xp2_ASAP7_75t_L g1777 ( 
.A(n_1757),
.B(n_1733),
.C(n_1749),
.D(n_1742),
.E(n_1751),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1747),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1733),
.A2(n_1716),
.B1(n_1729),
.B2(n_1722),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1742),
.B(n_1715),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1778),
.Y(n_1781)
);

AOI222xp33_ASAP7_75t_L g1782 ( 
.A1(n_1760),
.A2(n_1751),
.B1(n_1755),
.B2(n_1750),
.C1(n_1747),
.C2(n_1757),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1765),
.B(n_1755),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1763),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1761),
.B(n_1765),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1773),
.B(n_1779),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1773),
.B(n_1747),
.Y(n_1787)
);

NOR2x1_ASAP7_75t_L g1788 ( 
.A(n_1775),
.B(n_1750),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1762),
.B(n_1747),
.Y(n_1789)
);

INVxp67_ASAP7_75t_SL g1790 ( 
.A(n_1776),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1761),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1769),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1775),
.Y(n_1793)
);

AOI321xp33_ASAP7_75t_L g1794 ( 
.A1(n_1789),
.A2(n_1767),
.A3(n_1764),
.B1(n_1768),
.B2(n_1766),
.C(n_1777),
.Y(n_1794)
);

NAND2xp33_ASAP7_75t_L g1795 ( 
.A(n_1784),
.B(n_1740),
.Y(n_1795)
);

NAND4xp25_ASAP7_75t_SL g1796 ( 
.A(n_1782),
.B(n_1780),
.C(n_1770),
.D(n_1743),
.Y(n_1796)
);

AOI221x1_ASAP7_75t_L g1797 ( 
.A1(n_1781),
.A2(n_1774),
.B1(n_1772),
.B2(n_1768),
.C(n_1712),
.Y(n_1797)
);

OAI21xp33_ASAP7_75t_L g1798 ( 
.A1(n_1790),
.A2(n_1771),
.B(n_1743),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1788),
.A2(n_1700),
.B(n_1759),
.Y(n_1799)
);

AOI221xp5_ASAP7_75t_L g1800 ( 
.A1(n_1786),
.A2(n_1740),
.B1(n_1710),
.B2(n_1701),
.C(n_1731),
.Y(n_1800)
);

AOI211xp5_ASAP7_75t_L g1801 ( 
.A1(n_1786),
.A2(n_1758),
.B(n_1759),
.C(n_1726),
.Y(n_1801)
);

AOI221xp5_ASAP7_75t_L g1802 ( 
.A1(n_1793),
.A2(n_1758),
.B1(n_1722),
.B2(n_1727),
.C(n_1676),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1785),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1783),
.A2(n_1722),
.B(n_1685),
.Y(n_1804)
);

O2A1O1Ixp33_ASAP7_75t_SL g1805 ( 
.A1(n_1799),
.A2(n_1785),
.B(n_1791),
.C(n_1792),
.Y(n_1805)
);

OAI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1802),
.A2(n_1791),
.B1(n_1787),
.B2(n_1728),
.Y(n_1806)
);

OAI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1796),
.A2(n_1795),
.B(n_1798),
.Y(n_1807)
);

NAND2x1_ASAP7_75t_L g1808 ( 
.A(n_1803),
.B(n_1787),
.Y(n_1808)
);

AOI321xp33_ASAP7_75t_L g1809 ( 
.A1(n_1801),
.A2(n_1565),
.A3(n_1687),
.B1(n_1692),
.B2(n_1685),
.C(n_1684),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1797),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1808),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1805),
.Y(n_1812)
);

NOR2x1_ASAP7_75t_L g1813 ( 
.A(n_1810),
.B(n_1804),
.Y(n_1813)
);

OAI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1807),
.A2(n_1794),
.B1(n_1800),
.B2(n_1565),
.C(n_1687),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1809),
.B(n_1630),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1806),
.Y(n_1816)
);

INVxp67_ASAP7_75t_L g1817 ( 
.A(n_1808),
.Y(n_1817)
);

NAND2xp33_ASAP7_75t_R g1818 ( 
.A(n_1811),
.B(n_1439),
.Y(n_1818)
);

HB1xp67_ASAP7_75t_L g1819 ( 
.A(n_1817),
.Y(n_1819)
);

NOR2x1_ASAP7_75t_L g1820 ( 
.A(n_1812),
.B(n_1684),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1816),
.A2(n_1642),
.B1(n_1591),
.B2(n_1666),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1813),
.Y(n_1822)
);

NOR3x1_ASAP7_75t_L g1823 ( 
.A(n_1818),
.B(n_1814),
.C(n_1815),
.Y(n_1823)
);

OAI221xp5_ASAP7_75t_SL g1824 ( 
.A1(n_1822),
.A2(n_1692),
.B1(n_1681),
.B2(n_1666),
.C(n_1593),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1819),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1825),
.B(n_1823),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1826),
.A2(n_1824),
.B1(n_1820),
.B2(n_1821),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1827),
.Y(n_1828)
);

INVxp67_ASAP7_75t_SL g1829 ( 
.A(n_1827),
.Y(n_1829)
);

XNOR2xp5_ASAP7_75t_L g1830 ( 
.A(n_1828),
.B(n_1470),
.Y(n_1830)
);

BUFx2_ASAP7_75t_L g1831 ( 
.A(n_1829),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1831),
.B(n_1681),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1830),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1832),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1834),
.A2(n_1833),
.B(n_1620),
.Y(n_1835)
);

AOI222xp33_ASAP7_75t_L g1836 ( 
.A1(n_1835),
.A2(n_1647),
.B1(n_1646),
.B2(n_1637),
.C1(n_1634),
.C2(n_1638),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1836),
.A2(n_1630),
.B1(n_1635),
.B2(n_1636),
.Y(n_1837)
);

AOI221xp5_ASAP7_75t_L g1838 ( 
.A1(n_1837),
.A2(n_1647),
.B1(n_1646),
.B2(n_1634),
.C(n_1610),
.Y(n_1838)
);

AOI211xp5_ASAP7_75t_L g1839 ( 
.A1(n_1838),
.A2(n_1472),
.B(n_1439),
.C(n_1452),
.Y(n_1839)
);


endmodule