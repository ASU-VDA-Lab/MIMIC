module fake_jpeg_10236_n_118 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_118);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx10_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_8),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx8_ASAP7_75t_SL g58 ( 
.A(n_4),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_24),
.B(n_10),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_12),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_64),
.Y(n_85)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_69),
.Y(n_82)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_1),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_70),
.B(n_71),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_1),
.Y(n_71)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_65),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_72),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_52),
.B1(n_57),
.B2(n_50),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_74),
.A2(n_83),
.B1(n_84),
.B2(n_21),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_57),
.B1(n_61),
.B2(n_47),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_77),
.B(n_79),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_67),
.A2(n_49),
.B1(n_44),
.B2(n_54),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_56),
.B1(n_51),
.B2(n_23),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_25),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_59),
.B1(n_5),
.B2(n_2),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_7),
.Y(n_86)
);

AND2x4_ASAP7_75t_SL g90 ( 
.A(n_86),
.B(n_11),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_55),
.B1(n_45),
.B2(n_14),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_87),
.A2(n_45),
.B1(n_13),
.B2(n_16),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_92),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_26),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_27),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_94),
.B(n_97),
.C(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_104),
.B(n_98),
.Y(n_105)
);

FAx1_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_90),
.CI(n_96),
.CON(n_106),
.SN(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_102),
.C(n_100),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_99),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_109),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_112),
.Y(n_113)
);

AO21x2_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_89),
.B(n_95),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_114),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_28),
.C(n_30),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_34),
.C(n_36),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_91),
.B(n_38),
.Y(n_118)
);


endmodule