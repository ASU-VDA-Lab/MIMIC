module fake_jpeg_5306_n_44 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_44);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_17;
wire n_29;
wire n_37;
wire n_43;
wire n_32;
wire n_15;

INVx4_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_7),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_25),
.A2(n_10),
.B1(n_12),
.B2(n_2),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_21),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_30),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_5),
.B1(n_16),
.B2(n_18),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_23),
.B1(n_26),
.B2(n_19),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_13),
.B(n_18),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_17),
.C(n_20),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_34),
.B1(n_35),
.B2(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_39),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_37),
.A2(n_35),
.B(n_14),
.Y(n_39)
);

OA21x2_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_17),
.B(n_20),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_24),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_40),
.C(n_36),
.Y(n_43)
);

NOR5xp2_ASAP7_75t_SL g44 ( 
.A(n_43),
.B(n_24),
.C(n_27),
.D(n_15),
.E(n_22),
.Y(n_44)
);


endmodule