module real_aes_232_n_398 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_398);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_398;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_503;
wire n_635;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_1064;
wire n_540;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_948;
wire n_399;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_786;
wire n_512;
wire n_795;
wire n_816;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_1072;
wire n_994;
wire n_1078;
wire n_938;
wire n_744;
wire n_935;
wire n_1098;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_981;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_976;
wire n_872;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_517;
wire n_931;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_1081;
wire n_1084;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_754;
wire n_607;
wire n_449;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_1105;
wire n_902;
wire n_853;
wire n_1079;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1003;
wire n_1000;
wire n_1028;
wire n_1014;
wire n_727;
wire n_1083;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_1001;
wire n_494;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_1068;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_691;
wire n_481;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_922;
wire n_633;
wire n_482;
wire n_679;
wire n_926;
wire n_520;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_721;
wire n_446;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_1040;
wire n_652;
wire n_703;
wire n_601;
wire n_1101;
wire n_500;
wire n_661;
wire n_463;
wire n_1076;
wire n_804;
wire n_1102;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_1039;
wire n_424;
wire n_802;
wire n_868;
wire n_877;
wire n_574;
wire n_1069;
wire n_1024;
wire n_1104;
wire n_842;
wire n_849;
wire n_1061;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_0), .A2(n_346), .B1(n_597), .B2(n_598), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_1), .A2(n_238), .B1(n_605), .B2(n_763), .Y(n_762) );
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_2), .A2(n_294), .B1(n_451), .B2(n_496), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_3), .A2(n_128), .B1(n_438), .B2(n_442), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_4), .A2(n_140), .B1(n_512), .B2(n_694), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g879 ( .A(n_5), .Y(n_879) );
XOR2xp5_ASAP7_75t_L g1058 ( .A(n_6), .B(n_1059), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_7), .A2(n_93), .B1(n_517), .B2(n_737), .Y(n_935) );
AOI22xp5_ASAP7_75t_L g1006 ( .A1(n_8), .A2(n_209), .B1(n_734), .B2(n_847), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_9), .B(n_586), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_10), .A2(n_57), .B1(n_438), .B2(n_442), .Y(n_437) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_11), .A2(n_273), .B1(n_597), .B2(n_598), .Y(n_672) );
AOI22xp33_ASAP7_75t_SL g1066 ( .A1(n_12), .A2(n_344), .B1(n_474), .B2(n_533), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_13), .A2(n_201), .B1(n_468), .B2(n_471), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_14), .A2(n_385), .B1(n_648), .B2(n_868), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_15), .A2(n_219), .B1(n_607), .B2(n_608), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_16), .A2(n_89), .B1(n_469), .B2(n_471), .Y(n_535) );
AOI22xp33_ASAP7_75t_SL g903 ( .A1(n_17), .A2(n_92), .B1(n_527), .B2(n_593), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_18), .A2(n_111), .B1(n_465), .B2(n_468), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_19), .A2(n_342), .B1(n_476), .B2(n_531), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_20), .A2(n_204), .B1(n_438), .B2(n_702), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_21), .A2(n_261), .B1(n_633), .B2(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_22), .A2(n_94), .B1(n_803), .B2(n_847), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_23), .A2(n_239), .B1(n_591), .B2(n_667), .Y(n_904) );
AOI22xp33_ASAP7_75t_SL g676 ( .A1(n_24), .A2(n_193), .B1(n_605), .B2(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_25), .A2(n_367), .B1(n_618), .B2(n_863), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_26), .A2(n_161), .B1(n_428), .B2(n_498), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_27), .A2(n_71), .B1(n_496), .B2(n_524), .Y(n_523) );
AO222x2_ASAP7_75t_L g882 ( .A1(n_28), .A2(n_158), .B1(n_259), .B2(n_539), .C1(n_541), .C2(n_542), .Y(n_882) );
CKINVDCx20_ASAP7_75t_R g1074 ( .A(n_29), .Y(n_1074) );
CKINVDCx20_ASAP7_75t_R g1075 ( .A(n_30), .Y(n_1075) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_31), .A2(n_354), .B1(n_667), .B2(n_886), .Y(n_885) );
INVx1_ASAP7_75t_SL g416 ( .A(n_32), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g1045 ( .A(n_32), .B(n_49), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_33), .A2(n_361), .B1(n_476), .B2(n_480), .Y(n_644) );
CKINVDCx20_ASAP7_75t_R g899 ( .A(n_34), .Y(n_899) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_35), .A2(n_188), .B1(n_508), .B2(n_509), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_36), .A2(n_395), .B1(n_512), .B2(n_577), .Y(n_576) );
AOI22xp33_ASAP7_75t_SL g777 ( .A1(n_37), .A2(n_150), .B1(n_447), .B2(n_621), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_38), .B(n_630), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_39), .B(n_409), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_40), .A2(n_309), .B1(n_607), .B2(n_608), .Y(n_606) );
AOI22x1_ASAP7_75t_L g910 ( .A1(n_41), .A2(n_211), .B1(n_601), .B2(n_607), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_42), .A2(n_129), .B1(n_667), .B2(n_886), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_43), .A2(n_237), .B1(n_478), .B2(n_803), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_44), .A2(n_233), .B1(n_428), .B2(n_648), .Y(n_647) );
OA22x2_ASAP7_75t_L g956 ( .A1(n_45), .A2(n_957), .B1(n_958), .B2(n_984), .Y(n_956) );
CKINVDCx20_ASAP7_75t_R g984 ( .A(n_45), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_46), .A2(n_296), .B1(n_506), .B2(n_627), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_47), .A2(n_200), .B1(n_527), .B2(n_528), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_48), .A2(n_345), .B1(n_465), .B2(n_731), .Y(n_859) );
AO22x2_ASAP7_75t_L g418 ( .A1(n_49), .A2(n_376), .B1(n_415), .B2(n_419), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_50), .A2(n_186), .B1(n_600), .B2(n_788), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_51), .A2(n_230), .B1(n_457), .B2(n_518), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_52), .A2(n_378), .B1(n_468), .B2(n_618), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_53), .A2(n_62), .B1(n_451), .B2(n_496), .Y(n_495) );
AO21x1_ASAP7_75t_SL g1046 ( .A1(n_54), .A2(n_1047), .B(n_1055), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_55), .A2(n_163), .B1(n_730), .B2(n_731), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_56), .A2(n_299), .B1(n_460), .B2(n_465), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_58), .B(n_808), .Y(n_807) );
AO22x1_ASAP7_75t_L g1100 ( .A1(n_59), .A2(n_369), .B1(n_517), .B2(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g417 ( .A(n_60), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_61), .A2(n_328), .B1(n_604), .B2(n_608), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_63), .A2(n_255), .B1(n_478), .B2(n_733), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_64), .A2(n_313), .B1(n_428), .B2(n_433), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_65), .A2(n_311), .B1(n_476), .B2(n_478), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_66), .A2(n_325), .B1(n_607), .B2(n_674), .Y(n_673) );
AOI22xp33_ASAP7_75t_SL g1062 ( .A1(n_67), .A2(n_156), .B1(n_537), .B2(n_758), .Y(n_1062) );
CKINVDCx20_ASAP7_75t_R g835 ( .A(n_68), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_69), .A2(n_372), .B1(n_736), .B2(n_758), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_70), .A2(n_319), .B1(n_473), .B2(n_537), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_72), .A2(n_360), .B1(n_476), .B2(n_480), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_73), .B(n_409), .Y(n_408) );
AOI21xp5_ASAP7_75t_SL g1103 ( .A1(n_74), .A2(n_840), .B(n_1104), .Y(n_1103) );
AO22x2_ASAP7_75t_L g425 ( .A1(n_75), .A2(n_206), .B1(n_415), .B2(n_426), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_76), .A2(n_329), .B1(n_516), .B2(n_518), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_77), .A2(n_214), .B1(n_514), .B2(n_516), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_78), .A2(n_258), .B1(n_476), .B2(n_478), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_79), .A2(n_159), .B1(n_508), .B2(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_80), .A2(n_368), .B1(n_447), .B2(n_451), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_81), .A2(n_121), .B1(n_588), .B2(n_774), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_82), .A2(n_178), .B1(n_527), .B2(n_593), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_83), .A2(n_307), .B1(n_694), .B2(n_740), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_84), .A2(n_338), .B1(n_601), .B2(n_740), .Y(n_784) );
AOI22xp5_ASAP7_75t_L g911 ( .A1(n_85), .A2(n_182), .B1(n_608), .B2(n_674), .Y(n_911) );
AOI22xp33_ASAP7_75t_SL g1063 ( .A1(n_86), .A2(n_347), .B1(n_803), .B2(n_1064), .Y(n_1063) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_87), .A2(n_172), .B1(n_600), .B2(n_601), .Y(n_599) );
AOI22xp33_ASAP7_75t_SL g889 ( .A1(n_88), .A2(n_125), .B1(n_597), .B2(n_598), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_90), .A2(n_215), .B1(n_428), .B2(n_433), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_91), .A2(n_304), .B1(n_674), .B2(n_677), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_95), .A2(n_270), .B1(n_541), .B2(n_588), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g979 ( .A1(n_96), .A2(n_377), .B1(n_514), .B2(n_937), .C(n_980), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_97), .A2(n_116), .B1(n_736), .B2(n_737), .Y(n_735) );
AOI222xp33_ASAP7_75t_L g629 ( .A1(n_98), .A2(n_162), .B1(n_251), .B2(n_630), .C1(n_631), .C2(n_633), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_99), .B(n_630), .Y(n_994) );
AOI22xp33_ASAP7_75t_SL g839 ( .A1(n_100), .A2(n_207), .B1(n_524), .B2(n_840), .Y(n_839) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_101), .A2(n_257), .B1(n_457), .B2(n_473), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_102), .A2(n_249), .B1(n_480), .B2(n_803), .Y(n_939) );
AOI22xp5_ASAP7_75t_L g925 ( .A1(n_103), .A2(n_321), .B1(n_868), .B2(n_926), .Y(n_925) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_104), .A2(n_298), .B1(n_502), .B2(n_506), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_105), .A2(n_341), .B1(n_498), .B2(n_569), .Y(n_841) );
AO222x2_ASAP7_75t_L g664 ( .A1(n_106), .A2(n_229), .B1(n_381), .B2(n_539), .C1(n_591), .C2(n_593), .Y(n_664) );
AOI22xp33_ASAP7_75t_SL g686 ( .A1(n_107), .A2(n_141), .B1(n_687), .B2(n_688), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_108), .A2(n_252), .B1(n_562), .B2(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g962 ( .A(n_109), .Y(n_962) );
AOI22xp5_ASAP7_75t_L g993 ( .A1(n_110), .A2(n_254), .B1(n_650), .B2(n_749), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_112), .A2(n_272), .B1(n_471), .B2(n_473), .Y(n_470) );
AOI22xp33_ASAP7_75t_SL g669 ( .A1(n_113), .A2(n_275), .B1(n_541), .B2(n_588), .Y(n_669) );
AO22x1_ASAP7_75t_L g1099 ( .A1(n_114), .A2(n_375), .B1(n_468), .B2(n_922), .Y(n_1099) );
AOI222xp33_ASAP7_75t_L g927 ( .A1(n_115), .A2(n_190), .B1(n_359), .B2(n_442), .C1(n_491), .C2(n_631), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_117), .A2(n_174), .B1(n_593), .B2(n_668), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_118), .A2(n_149), .B1(n_1068), .B2(n_1069), .Y(n_1067) );
AOI22xp5_ASAP7_75t_L g936 ( .A1(n_119), .A2(n_208), .B1(n_937), .B2(n_938), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_120), .A2(n_231), .B1(n_840), .B2(n_1079), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_122), .A2(n_351), .B1(n_460), .B2(n_736), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_123), .B(n_719), .Y(n_718) );
AO22x2_ASAP7_75t_L g422 ( .A1(n_124), .A2(n_302), .B1(n_415), .B2(n_423), .Y(n_422) );
CKINVDCx20_ASAP7_75t_R g971 ( .A(n_126), .Y(n_971) );
OAI22x1_ASAP7_75t_L g520 ( .A1(n_127), .A2(n_521), .B1(n_543), .B2(n_544), .Y(n_520) );
CKINVDCx16_ASAP7_75t_R g544 ( .A(n_127), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_130), .A2(n_170), .B1(n_706), .B2(n_707), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_131), .A2(n_393), .B1(n_509), .B2(n_736), .Y(n_805) );
AO21x2_ASAP7_75t_L g930 ( .A1(n_132), .A2(n_931), .B(n_950), .Y(n_930) );
NOR2xp33_ASAP7_75t_L g950 ( .A(n_132), .B(n_933), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_133), .A2(n_137), .B1(n_816), .B2(n_946), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_134), .A2(n_245), .B1(n_460), .B2(n_625), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g1106 ( .A1(n_135), .A2(n_366), .B1(n_944), .B2(n_948), .Y(n_1106) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_136), .A2(n_157), .B1(n_509), .B2(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_138), .A2(n_263), .B1(n_621), .B2(n_866), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_139), .A2(n_286), .B1(n_726), .B2(n_727), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_142), .A2(n_266), .B1(n_731), .B2(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g928 ( .A(n_143), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_144), .A2(n_365), .B1(n_598), .B2(n_1023), .Y(n_1022) );
OA22x2_ASAP7_75t_L g987 ( .A1(n_145), .A2(n_988), .B1(n_989), .B2(n_990), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_145), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_146), .A2(n_320), .B1(n_531), .B2(n_1095), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_147), .A2(n_223), .B1(n_605), .B2(n_763), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_148), .B(n_409), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_151), .A2(n_256), .B1(n_469), .B2(n_618), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_152), .A2(n_184), .B1(n_625), .B2(n_1009), .Y(n_1008) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_153), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_154), .A2(n_247), .B1(n_512), .B2(n_642), .Y(n_641) );
OA22x2_ASAP7_75t_L g714 ( .A1(n_155), .A2(n_715), .B1(n_716), .B2(n_741), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_155), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g890 ( .A1(n_160), .A2(n_171), .B1(n_674), .B2(n_677), .Y(n_890) );
CKINVDCx20_ASAP7_75t_R g996 ( .A(n_164), .Y(n_996) );
CKINVDCx20_ASAP7_75t_R g974 ( .A(n_165), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_166), .A2(n_191), .B1(n_926), .B2(n_944), .Y(n_943) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_167), .A2(n_243), .B1(n_457), .B2(n_460), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g869 ( .A1(n_168), .A2(n_262), .B1(n_438), .B2(n_650), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_169), .B(n_702), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_173), .A2(n_240), .B1(n_460), .B2(n_533), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g1005 ( .A1(n_175), .A2(n_394), .B1(n_731), .B2(n_845), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_176), .B(n_630), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_177), .A2(n_305), .B1(n_480), .B2(n_734), .Y(n_759) );
AO22x1_ASAP7_75t_L g1097 ( .A1(n_179), .A2(n_253), .B1(n_845), .B2(n_1098), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_180), .A2(n_199), .B1(n_642), .B2(n_740), .Y(n_739) );
AOI22xp33_ASAP7_75t_SL g782 ( .A1(n_181), .A2(n_337), .B1(n_476), .B2(n_783), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_183), .A2(n_308), .B1(n_457), .B2(n_518), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_185), .A2(n_370), .B1(n_600), .B2(n_850), .Y(n_849) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_187), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_189), .A2(n_288), .B1(n_433), .B2(n_569), .Y(n_968) );
CKINVDCx20_ASAP7_75t_R g1001 ( .A(n_192), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_194), .B(n_491), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_195), .A2(n_396), .B1(n_633), .B2(n_816), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g964 ( .A(n_196), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_197), .A2(n_226), .B1(n_496), .B2(n_621), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_198), .A2(n_283), .B1(n_451), .B2(n_496), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g998 ( .A(n_202), .Y(n_998) );
AOI22xp33_ASAP7_75t_SL g690 ( .A1(n_203), .A2(n_331), .B1(n_516), .B2(n_691), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_205), .A2(n_271), .B1(n_754), .B2(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g1044 ( .A(n_206), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_210), .A2(n_250), .B1(n_607), .B2(n_608), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_212), .A2(n_278), .B1(n_597), .B2(n_598), .Y(n_907) );
CKINVDCx20_ASAP7_75t_R g978 ( .A(n_213), .Y(n_978) );
CKINVDCx20_ASAP7_75t_R g1105 ( .A(n_216), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_217), .A2(n_330), .B1(n_926), .B2(n_944), .Y(n_1081) );
XNOR2xp5_ASAP7_75t_L g894 ( .A(n_218), .B(n_895), .Y(n_894) );
XNOR2xp5_ASAP7_75t_L g913 ( .A(n_218), .B(n_895), .Y(n_913) );
CKINVDCx20_ASAP7_75t_R g976 ( .A(n_220), .Y(n_976) );
AOI22xp5_ASAP7_75t_L g1082 ( .A1(n_221), .A2(n_1083), .B1(n_1086), .B2(n_1088), .Y(n_1082) );
OA22x2_ASAP7_75t_L g1090 ( .A1(n_221), .A2(n_1091), .B1(n_1092), .B2(n_1110), .Y(n_1090) );
INVx1_ASAP7_75t_L g1110 ( .A(n_221), .Y(n_1110) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_222), .A2(n_379), .B1(n_496), .B2(n_524), .Y(n_752) );
INVx1_ASAP7_75t_L g697 ( .A(n_224), .Y(n_697) );
AOI22xp33_ASAP7_75t_SL g666 ( .A1(n_225), .A2(n_336), .B1(n_667), .B2(n_668), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_227), .A2(n_405), .B1(n_406), .B2(n_482), .Y(n_404) );
INVxp67_ASAP7_75t_L g482 ( .A(n_227), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g981 ( .A(n_228), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_232), .A2(n_297), .B1(n_798), .B2(n_799), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_234), .A2(n_333), .B1(n_642), .B2(n_740), .Y(n_800) );
OA22x2_ASAP7_75t_L g854 ( .A1(n_235), .A2(n_855), .B1(n_856), .B2(n_871), .Y(n_854) );
INVxp67_ASAP7_75t_L g871 ( .A(n_235), .Y(n_871) );
OA22x2_ASAP7_75t_L g873 ( .A1(n_235), .A2(n_855), .B1(n_856), .B2(n_871), .Y(n_873) );
XNOR2x1_ASAP7_75t_L g553 ( .A(n_236), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g1052 ( .A(n_241), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_242), .A2(n_389), .B1(n_604), .B2(n_605), .Y(n_892) );
AOI22xp33_ASAP7_75t_SL g511 ( .A1(n_244), .A2(n_291), .B1(n_512), .B2(n_514), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_246), .A2(n_264), .B1(n_788), .B2(n_922), .Y(n_921) );
CKINVDCx20_ASAP7_75t_R g1072 ( .A(n_248), .Y(n_1072) );
CKINVDCx20_ASAP7_75t_R g982 ( .A(n_260), .Y(n_982) );
CKINVDCx16_ASAP7_75t_R g1028 ( .A(n_265), .Y(n_1028) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_267), .A2(n_681), .B1(n_682), .B2(n_708), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_267), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_268), .A2(n_661), .B1(n_662), .B2(n_679), .Y(n_660) );
INVx1_ASAP7_75t_L g679 ( .A(n_268), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_269), .A2(n_358), .B1(n_721), .B2(n_779), .Y(n_778) );
AOI22xp5_ASAP7_75t_L g1016 ( .A1(n_274), .A2(n_356), .B1(n_541), .B2(n_542), .Y(n_1016) );
CKINVDCx20_ASAP7_75t_R g898 ( .A(n_276), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_277), .A2(n_318), .B1(n_496), .B2(n_524), .Y(n_967) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_279), .A2(n_289), .B1(n_438), .B2(n_442), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_280), .A2(n_334), .B1(n_648), .B2(n_721), .Y(n_720) );
AOI22xp33_ASAP7_75t_SL g884 ( .A1(n_281), .A2(n_300), .B1(n_593), .B2(n_668), .Y(n_884) );
AO22x2_ASAP7_75t_L g635 ( .A1(n_282), .A2(n_636), .B1(n_653), .B2(n_654), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_282), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_284), .A2(n_397), .B1(n_605), .B2(n_763), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_285), .B(n_630), .Y(n_942) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_287), .A2(n_316), .B1(n_442), .B2(n_749), .Y(n_748) );
AOI22x1_ASAP7_75t_L g485 ( .A1(n_290), .A2(n_486), .B1(n_487), .B2(n_519), .Y(n_485) );
INVx1_ASAP7_75t_L g519 ( .A(n_290), .Y(n_519) );
XNOR2x1_ASAP7_75t_L g547 ( .A(n_290), .B(n_487), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_292), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_293), .A2(n_374), .B1(n_473), .B2(n_537), .Y(n_761) );
OA22x2_ASAP7_75t_L g792 ( .A1(n_295), .A2(n_793), .B1(n_794), .B2(n_795), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_295), .Y(n_793) );
AOI22xp33_ASAP7_75t_SL g685 ( .A1(n_301), .A2(n_348), .B1(n_509), .B2(n_580), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g1042 ( .A(n_302), .B(n_1043), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_303), .A2(n_373), .B1(n_438), .B2(n_650), .Y(n_649) );
AOI222xp33_ASAP7_75t_L g538 ( .A1(n_306), .A2(n_317), .B1(n_355), .B2(n_539), .C1(n_540), .C2(n_542), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_310), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_312), .Y(n_837) );
CKINVDCx20_ASAP7_75t_R g900 ( .A(n_314), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_315), .A2(n_349), .B1(n_813), .B2(n_948), .Y(n_947) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_322), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g860 ( .A1(n_323), .A2(n_339), .B1(n_783), .B2(n_861), .Y(n_860) );
AOI22xp5_ASAP7_75t_L g1108 ( .A1(n_324), .A2(n_353), .B1(n_723), .B2(n_1109), .Y(n_1108) );
INVx1_ASAP7_75t_L g852 ( .A(n_326), .Y(n_852) );
INVx3_ASAP7_75t_L g415 ( .A(n_327), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_332), .A2(n_340), .B1(n_604), .B2(n_605), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_335), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_343), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g812 ( .A1(n_350), .A2(n_382), .B1(n_524), .B2(n_813), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_352), .A2(n_386), .B1(n_465), .B2(n_518), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_357), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g1002 ( .A(n_362), .Y(n_1002) );
INVx1_ASAP7_75t_L g767 ( .A(n_363), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_364), .A2(n_392), .B1(n_428), .B2(n_754), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_371), .A2(n_384), .B1(n_496), .B2(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g1039 ( .A(n_380), .Y(n_1039) );
AND2x4_ASAP7_75t_L g1054 ( .A(n_380), .B(n_1040), .Y(n_1054) );
AO21x1_ASAP7_75t_L g1084 ( .A1(n_380), .A2(n_1050), .B(n_1085), .Y(n_1084) );
INVx1_ASAP7_75t_L g1040 ( .A(n_383), .Y(n_1040) );
AND2x2_ASAP7_75t_R g1057 ( .A(n_383), .B(n_1039), .Y(n_1057) );
OA22x2_ASAP7_75t_L g612 ( .A1(n_387), .A2(n_613), .B1(n_614), .B2(n_634), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g613 ( .A(n_387), .Y(n_613) );
INVxp67_ASAP7_75t_L g1051 ( .A(n_388), .Y(n_1051) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_390), .B(n_539), .Y(n_1015) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_391), .Y(n_564) );
O2A1O1Ixp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_823), .B(n_1035), .C(n_1046), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g1035 ( .A1(n_399), .A2(n_823), .B(n_1036), .Y(n_1035) );
XNOR2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_711), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_550), .B1(n_709), .B2(n_710), .Y(n_400) );
INVx2_ASAP7_75t_L g709 ( .A(n_401), .Y(n_709) );
INVx2_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
OA22x2_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_483), .B1(n_548), .B2(n_549), .Y(n_402) );
HB1xp67_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g548 ( .A(n_404), .Y(n_548) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NOR2xp67_ASAP7_75t_L g406 ( .A(n_407), .B(n_455), .Y(n_406) );
NAND4xp25_ASAP7_75t_L g407 ( .A(n_408), .B(n_427), .C(n_437), .D(n_446), .Y(n_407) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_409), .Y(n_719) );
INVx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx4_ASAP7_75t_SL g491 ( .A(n_410), .Y(n_491) );
INVx4_ASAP7_75t_SL g586 ( .A(n_410), .Y(n_586) );
INVx3_ASAP7_75t_L g630 ( .A(n_410), .Y(n_630) );
INVx3_ASAP7_75t_SL g700 ( .A(n_410), .Y(n_700) );
BUFx2_ASAP7_75t_L g1073 ( .A(n_410), .Y(n_1073) );
INVx6_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_420), .Y(n_411) );
AND2x4_ASAP7_75t_L g435 ( .A(n_412), .B(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g452 ( .A(n_412), .B(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g528 ( .A(n_412), .B(n_436), .Y(n_528) );
AND2x4_ASAP7_75t_L g539 ( .A(n_412), .B(n_420), .Y(n_539) );
AND2x2_ASAP7_75t_L g591 ( .A(n_412), .B(n_453), .Y(n_591) );
AND2x2_ASAP7_75t_L g593 ( .A(n_412), .B(n_436), .Y(n_593) );
AND2x2_ASAP7_75t_L g886 ( .A(n_412), .B(n_453), .Y(n_886) );
AND2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_418), .Y(n_412) );
INVx2_ASAP7_75t_L g432 ( .A(n_413), .Y(n_432) );
AND2x2_ASAP7_75t_L g440 ( .A(n_413), .B(n_441), .Y(n_440) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_413), .Y(n_445) );
OAI22x1_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_415), .B1(n_416), .B2(n_417), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g419 ( .A(n_415), .Y(n_419) );
INVx2_ASAP7_75t_L g423 ( .A(n_415), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_415), .Y(n_426) );
AND2x2_ASAP7_75t_L g431 ( .A(n_418), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g441 ( .A(n_418), .Y(n_441) );
BUFx2_ASAP7_75t_L g481 ( .A(n_418), .Y(n_481) );
AND2x2_ASAP7_75t_L g459 ( .A(n_420), .B(n_431), .Y(n_459) );
AND2x4_ASAP7_75t_L g467 ( .A(n_420), .B(n_463), .Y(n_467) );
AND2x4_ASAP7_75t_L g472 ( .A(n_420), .B(n_440), .Y(n_472) );
AND2x2_ASAP7_75t_L g604 ( .A(n_420), .B(n_440), .Y(n_604) );
AND2x6_ASAP7_75t_L g607 ( .A(n_420), .B(n_431), .Y(n_607) );
AND2x2_ASAP7_75t_L g674 ( .A(n_420), .B(n_463), .Y(n_674) );
AND2x2_ASAP7_75t_L g763 ( .A(n_420), .B(n_440), .Y(n_763) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_424), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g430 ( .A(n_422), .B(n_424), .Y(n_430) );
AND2x2_ASAP7_75t_L g444 ( .A(n_422), .B(n_425), .Y(n_444) );
INVx1_ASAP7_75t_L g450 ( .A(n_422), .Y(n_450) );
INVxp67_ASAP7_75t_L g436 ( .A(n_424), .Y(n_436) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g449 ( .A(n_425), .B(n_450), .Y(n_449) );
BUFx3_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_429), .Y(n_569) );
BUFx2_ASAP7_75t_L g721 ( .A(n_429), .Y(n_721) );
BUFx2_ASAP7_75t_L g868 ( .A(n_429), .Y(n_868) );
AND2x4_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
AND2x2_ASAP7_75t_L g439 ( .A(n_430), .B(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g474 ( .A(n_430), .B(n_463), .Y(n_474) );
AND2x2_ASAP7_75t_L g527 ( .A(n_430), .B(n_431), .Y(n_527) );
AND2x4_ASAP7_75t_L g541 ( .A(n_430), .B(n_440), .Y(n_541) );
AND2x2_ASAP7_75t_L g668 ( .A(n_430), .B(n_431), .Y(n_668) );
AND2x2_ASAP7_75t_L g677 ( .A(n_430), .B(n_463), .Y(n_677) );
AND2x2_ASAP7_75t_L g477 ( .A(n_431), .B(n_449), .Y(n_477) );
AND2x2_ASAP7_75t_SL g597 ( .A(n_431), .B(n_449), .Y(n_597) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_431), .B(n_449), .Y(n_1023) );
AND2x4_ASAP7_75t_L g463 ( .A(n_432), .B(n_441), .Y(n_463) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_SL g498 ( .A(n_434), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_434), .A2(n_567), .B1(n_568), .B2(n_570), .Y(n_566) );
INVx1_ASAP7_75t_L g648 ( .A(n_434), .Y(n_648) );
INVx2_ASAP7_75t_SL g707 ( .A(n_434), .Y(n_707) );
INVx2_ASAP7_75t_L g754 ( .A(n_434), .Y(n_754) );
INVx2_ASAP7_75t_L g779 ( .A(n_434), .Y(n_779) );
INVx2_ASAP7_75t_L g926 ( .A(n_434), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g1000 ( .A1(n_434), .A2(n_568), .B1(n_1001), .B2(n_1002), .Y(n_1000) );
NOR2xp33_ASAP7_75t_L g1104 ( .A(n_434), .B(n_1105), .Y(n_1104) );
INVx6_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx5_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g632 ( .A(n_439), .Y(n_632) );
BUFx3_ASAP7_75t_L g724 ( .A(n_439), .Y(n_724) );
BUFx3_ASAP7_75t_L g817 ( .A(n_439), .Y(n_817) );
AND2x2_ASAP7_75t_L g448 ( .A(n_440), .B(n_449), .Y(n_448) );
AND2x4_ASAP7_75t_L g667 ( .A(n_440), .B(n_449), .Y(n_667) );
BUFx3_ASAP7_75t_L g633 ( .A(n_442), .Y(n_633) );
INVx2_ASAP7_75t_L g1076 ( .A(n_442), .Y(n_1076) );
BUFx12f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx3_ASAP7_75t_L g651 ( .A(n_443), .Y(n_651) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
AND2x4_ASAP7_75t_L g469 ( .A(n_444), .B(n_463), .Y(n_469) );
AND2x4_ASAP7_75t_L g480 ( .A(n_444), .B(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_SL g542 ( .A(n_444), .B(n_445), .Y(n_542) );
AND2x2_ASAP7_75t_SL g588 ( .A(n_444), .B(n_445), .Y(n_588) );
AND2x4_ASAP7_75t_L g598 ( .A(n_444), .B(n_481), .Y(n_598) );
AND2x4_ASAP7_75t_L g605 ( .A(n_444), .B(n_463), .Y(n_605) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_447), .Y(n_726) );
INVx1_ASAP7_75t_L g997 ( .A(n_447), .Y(n_997) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_448), .Y(n_496) );
INVx3_ASAP7_75t_L g563 ( .A(n_448), .Y(n_563) );
AND2x4_ASAP7_75t_L g462 ( .A(n_449), .B(n_463), .Y(n_462) );
AND2x6_ASAP7_75t_L g608 ( .A(n_449), .B(n_463), .Y(n_608) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_450), .Y(n_454) );
INVxp67_ASAP7_75t_L g565 ( .A(n_451), .Y(n_565) );
BUFx4f_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g525 ( .A(n_452), .Y(n_525) );
BUFx6f_ASAP7_75t_SL g621 ( .A(n_452), .Y(n_621) );
BUFx3_ASAP7_75t_L g949 ( .A(n_452), .Y(n_949) );
INVx1_ASAP7_75t_L g1080 ( .A(n_452), .Y(n_1080) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND4xp25_ASAP7_75t_L g455 ( .A(n_456), .B(n_464), .C(n_470), .D(n_475), .Y(n_455) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_SL g508 ( .A(n_458), .Y(n_508) );
INVx2_ASAP7_75t_SL g580 ( .A(n_458), .Y(n_580) );
INVx3_ASAP7_75t_L g736 ( .A(n_458), .Y(n_736) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx2_ASAP7_75t_L g533 ( .A(n_459), .Y(n_533) );
BUFx2_ASAP7_75t_L g845 ( .A(n_459), .Y(n_845) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_SL g509 ( .A(n_461), .Y(n_509) );
INVx1_ASAP7_75t_SL g640 ( .A(n_461), .Y(n_640) );
INVx2_ASAP7_75t_L g731 ( .A(n_461), .Y(n_731) );
INVx2_ASAP7_75t_SL g758 ( .A(n_461), .Y(n_758) );
INVx2_ASAP7_75t_L g938 ( .A(n_461), .Y(n_938) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_461), .Y(n_983) );
INVx2_ASAP7_75t_L g1098 ( .A(n_461), .Y(n_1098) );
INVx8_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx2_ASAP7_75t_L g798 ( .A(n_465), .Y(n_798) );
INVx2_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
INVx4_ASAP7_75t_L g517 ( .A(n_466), .Y(n_517) );
INVx2_ASAP7_75t_L g537 ( .A(n_466), .Y(n_537) );
INVx3_ASAP7_75t_SL g600 ( .A(n_466), .Y(n_600) );
INVx2_ASAP7_75t_SL g625 ( .A(n_466), .Y(n_625) );
INVx8_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx2_ASAP7_75t_SL g514 ( .A(n_469), .Y(n_514) );
INVx2_ASAP7_75t_L g643 ( .A(n_469), .Y(n_643) );
BUFx2_ASAP7_75t_SL g694 ( .A(n_469), .Y(n_694) );
BUFx3_ASAP7_75t_L g788 ( .A(n_469), .Y(n_788) );
BUFx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx6_ASAP7_75t_L g513 ( .A(n_472), .Y(n_513) );
BUFx3_ASAP7_75t_L g740 ( .A(n_472), .Y(n_740) );
INVx1_ASAP7_75t_L g578 ( .A(n_473), .Y(n_578) );
HB1xp67_ASAP7_75t_L g850 ( .A(n_473), .Y(n_850) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx3_ASAP7_75t_L g518 ( .A(n_474), .Y(n_518) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_474), .Y(n_601) );
INVx2_ASAP7_75t_L g692 ( .A(n_474), .Y(n_692) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g505 ( .A(n_477), .Y(n_505) );
BUFx3_ASAP7_75t_L g734 ( .A(n_477), .Y(n_734) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx3_ASAP7_75t_L g506 ( .A(n_479), .Y(n_506) );
INVx2_ASAP7_75t_L g688 ( .A(n_479), .Y(n_688) );
OAI22xp33_ASAP7_75t_L g970 ( .A1(n_479), .A2(n_971), .B1(n_972), .B2(n_974), .Y(n_970) );
INVx2_ASAP7_75t_L g1064 ( .A(n_479), .Y(n_1064) );
INVx5_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
BUFx2_ASAP7_75t_L g531 ( .A(n_480), .Y(n_531) );
BUFx2_ASAP7_75t_L g783 ( .A(n_480), .Y(n_783) );
BUFx3_ASAP7_75t_L g847 ( .A(n_480), .Y(n_847) );
INVx2_ASAP7_75t_L g549 ( .A(n_483), .Y(n_549) );
AO22x2_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_520), .B1(n_545), .B2(n_546), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_488), .B(n_499), .Y(n_487) );
NOR2xp67_ASAP7_75t_L g488 ( .A(n_489), .B(n_494), .Y(n_488) );
OAI21xp5_ASAP7_75t_SL g489 ( .A1(n_490), .A2(n_492), .B(n_493), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_497), .Y(n_494) );
BUFx6f_ASAP7_75t_SL g840 ( .A(n_496), .Y(n_840) );
NOR2x1_ASAP7_75t_L g499 ( .A(n_500), .B(n_510), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_507), .Y(n_500) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g973 ( .A(n_503), .Y(n_973) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g628 ( .A(n_504), .Y(n_628) );
BUFx6f_ASAP7_75t_L g861 ( .A(n_504), .Y(n_861) );
HB1xp67_ASAP7_75t_L g1095 ( .A(n_504), .Y(n_1095) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g804 ( .A(n_505), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_515), .Y(n_510) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx3_ASAP7_75t_L g618 ( .A(n_513), .Y(n_618) );
INVx2_ASAP7_75t_L g922 ( .A(n_513), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_513), .A2(n_981), .B1(n_982), .B2(n_983), .Y(n_980) );
INVx1_ASAP7_75t_SL g1068 ( .A(n_513), .Y(n_1068) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g977 ( .A(n_517), .Y(n_977) );
BUFx2_ASAP7_75t_L g799 ( .A(n_518), .Y(n_799) );
INVx2_ASAP7_75t_L g545 ( .A(n_520), .Y(n_545) );
NAND4xp25_ASAP7_75t_SL g521 ( .A(n_522), .B(n_529), .C(n_534), .D(n_538), .Y(n_521) );
AND4x1_ASAP7_75t_L g543 ( .A(n_522), .B(n_529), .C(n_534), .D(n_538), .Y(n_543) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_526), .Y(n_522) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .Y(n_529) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
INVx2_ASAP7_75t_SL g771 ( .A(n_539), .Y(n_771) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_SL g775 ( .A(n_541), .Y(n_775) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g710 ( .A(n_550), .Y(n_710) );
XOR2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_656), .Y(n_550) );
XNOR2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_610), .Y(n_551) );
XOR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_581), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_571), .Y(n_554) );
NOR3xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_559), .C(n_566), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_557), .B(n_558), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B1(n_564), .B2(n_565), .Y(n_559) );
INVx2_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
INVx4_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g814 ( .A(n_563), .Y(n_814) );
INVx2_ASAP7_75t_L g866 ( .A(n_563), .Y(n_866) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
BUFx4f_ASAP7_75t_SL g706 ( .A(n_569), .Y(n_706) );
BUFx2_ASAP7_75t_L g811 ( .A(n_569), .Y(n_811) );
BUFx2_ASAP7_75t_L g944 ( .A(n_569), .Y(n_944) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_575), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_579), .Y(n_575) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_581), .A2(n_765), .B1(n_766), .B2(n_820), .Y(n_819) );
INVx1_ASAP7_75t_SL g820 ( .A(n_581), .Y(n_820) );
XOR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_609), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_583), .B(n_594), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_584), .B(n_589), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
INVx1_ASAP7_75t_SL g961 ( .A(n_586), .Y(n_961) );
INVxp67_ASAP7_75t_L g901 ( .A(n_588), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_595), .B(n_602), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_599), .Y(n_595) );
INVx2_ASAP7_75t_L g738 ( .A(n_601), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_606), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B1(n_635), .B2(n_655), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_SL g634 ( .A(n_614), .Y(n_634) );
NAND4xp75_ASAP7_75t_L g614 ( .A(n_615), .B(n_619), .C(n_623), .D(n_629), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
BUFx2_ASAP7_75t_SL g727 ( .A(n_621), .Y(n_727) );
INVxp67_ASAP7_75t_L g999 ( .A(n_621), .Y(n_999) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
BUFx2_ASAP7_75t_L g730 ( .A(n_625), .Y(n_730) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g687 ( .A(n_628), .Y(n_687) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g749 ( .A(n_632), .Y(n_749) );
INVx1_ASAP7_75t_L g836 ( .A(n_633), .Y(n_836) );
INVx2_ASAP7_75t_L g655 ( .A(n_635), .Y(n_655) );
INVx1_ASAP7_75t_SL g654 ( .A(n_636), .Y(n_654) );
NOR2x1_ASAP7_75t_L g636 ( .A(n_637), .B(n_645), .Y(n_636) );
NAND4xp25_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .C(n_641), .D(n_644), .Y(n_637) );
INVx2_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_SL g863 ( .A(n_643), .Y(n_863) );
NAND4xp25_ASAP7_75t_SL g645 ( .A(n_646), .B(n_647), .C(n_649), .D(n_652), .Y(n_645) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx3_ASAP7_75t_L g702 ( .A(n_651), .Y(n_702) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
XNOR2x1_ASAP7_75t_L g657 ( .A(n_658), .B(n_680), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_663), .B(n_670), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_669), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_675), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
INVx1_ASAP7_75t_SL g708 ( .A(n_682), .Y(n_708) );
AND2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_695), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_689), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_693), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g1009 ( .A(n_692), .Y(n_1009) );
INVx2_ASAP7_75t_L g1101 ( .A(n_692), .Y(n_1101) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_703), .Y(n_695) );
OAI21xp33_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_698), .B(n_701), .Y(n_696) );
OAI222xp33_ASAP7_75t_L g831 ( .A1(n_698), .A2(n_832), .B1(n_834), .B2(n_835), .C1(n_836), .C2(n_837), .Y(n_831) );
INVx3_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
BUFx6f_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g809 ( .A(n_700), .Y(n_809) );
BUFx6f_ASAP7_75t_L g946 ( .A(n_702), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_790), .B1(n_821), .B2(n_822), .Y(n_711) );
INVx2_ASAP7_75t_L g821 ( .A(n_712), .Y(n_821) );
AOI22x1_ASAP7_75t_SL g712 ( .A1(n_713), .A2(n_714), .B1(n_742), .B2(n_789), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g741 ( .A(n_716), .Y(n_741) );
OR2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_728), .Y(n_716) );
NAND4xp25_ASAP7_75t_SL g717 ( .A(n_718), .B(n_720), .C(n_722), .D(n_725), .Y(n_717) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND4xp25_ASAP7_75t_L g728 ( .A(n_729), .B(n_732), .C(n_735), .D(n_739), .Y(n_728) );
BUFx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OAI22xp33_ASAP7_75t_L g975 ( .A1(n_738), .A2(n_976), .B1(n_977), .B2(n_978), .Y(n_975) );
INVx2_ASAP7_75t_L g789 ( .A(n_742), .Y(n_789) );
OA22x2_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_744), .B1(n_765), .B2(n_766), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
XOR2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_764), .Y(n_744) );
NAND2x1p5_ASAP7_75t_L g745 ( .A(n_746), .B(n_755), .Y(n_745) );
NOR2x1_ASAP7_75t_L g746 ( .A(n_747), .B(n_751), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_748), .B(n_750), .Y(n_747) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_749), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
NOR2x1_ASAP7_75t_L g755 ( .A(n_756), .B(n_760), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_759), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
INVx2_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
XNOR2x1_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
NAND2x1_ASAP7_75t_L g768 ( .A(n_769), .B(n_780), .Y(n_768) );
NOR2xp67_ASAP7_75t_L g769 ( .A(n_770), .B(n_776), .Y(n_769) );
OAI21xp5_ASAP7_75t_SL g770 ( .A1(n_771), .A2(n_772), .B(n_773), .Y(n_770) );
OAI222xp33_ASAP7_75t_L g897 ( .A1(n_771), .A2(n_775), .B1(n_898), .B2(n_899), .C1(n_900), .C2(n_901), .Y(n_897) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_785), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_784), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
BUFx6f_ASAP7_75t_L g1069 ( .A(n_788), .Y(n_1069) );
INVx3_ASAP7_75t_L g822 ( .A(n_790), .Y(n_822) );
OA22x2_ASAP7_75t_L g790 ( .A1(n_791), .A2(n_792), .B1(n_818), .B2(n_819), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NOR3x1_ASAP7_75t_SL g795 ( .A(n_796), .B(n_801), .C(n_806), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_797), .B(n_800), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_802), .B(n_805), .Y(n_801) );
BUFx6f_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
NAND4xp25_ASAP7_75t_SL g806 ( .A(n_807), .B(n_810), .C(n_812), .D(n_815), .Y(n_806) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
BUFx3_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g963 ( .A(n_816), .Y(n_963) );
BUFx6f_ASAP7_75t_SL g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
XNOR2x1_ASAP7_75t_L g825 ( .A(n_826), .B(n_953), .Y(n_825) );
OA22x2_ASAP7_75t_L g826 ( .A1(n_827), .A2(n_874), .B1(n_875), .B2(n_952), .Y(n_826) );
INVx1_ASAP7_75t_L g952 ( .A(n_827), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_853), .B1(n_872), .B2(n_873), .Y(n_827) );
INVx3_ASAP7_75t_L g872 ( .A(n_828), .Y(n_872) );
XOR2x2_ASAP7_75t_L g828 ( .A(n_829), .B(n_852), .Y(n_828) );
NAND2xp5_ASAP7_75t_SL g829 ( .A(n_830), .B(n_842), .Y(n_829) );
NOR2x1_ASAP7_75t_L g830 ( .A(n_831), .B(n_838), .Y(n_830) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_841), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g842 ( .A(n_843), .B(n_848), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_844), .B(n_846), .Y(n_843) );
BUFx3_ASAP7_75t_L g937 ( .A(n_845), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_849), .B(n_851), .Y(n_848) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx2_ASAP7_75t_SL g855 ( .A(n_856), .Y(n_855) );
NOR2x1_ASAP7_75t_L g856 ( .A(n_857), .B(n_864), .Y(n_856) );
NAND4xp25_ASAP7_75t_SL g857 ( .A(n_858), .B(n_859), .C(n_860), .D(n_862), .Y(n_857) );
NAND4xp25_ASAP7_75t_L g864 ( .A(n_865), .B(n_867), .C(n_869), .D(n_870), .Y(n_864) );
INVx2_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
AOI22x1_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_929), .B1(n_930), .B2(n_951), .Y(n_875) );
INVx2_ASAP7_75t_L g951 ( .A(n_876), .Y(n_951) );
XNOR2x1_ASAP7_75t_L g876 ( .A(n_877), .B(n_914), .Y(n_876) );
OAI21xp5_ASAP7_75t_L g877 ( .A1(n_878), .A2(n_894), .B(n_912), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_878), .B(n_913), .Y(n_912) );
XNOR2x1_ASAP7_75t_L g878 ( .A(n_879), .B(n_880), .Y(n_878) );
AND2x2_ASAP7_75t_L g880 ( .A(n_881), .B(n_887), .Y(n_880) );
NOR2xp33_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_884), .B(n_885), .Y(n_883) );
NOR2xp33_ASAP7_75t_L g887 ( .A(n_888), .B(n_891), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_889), .B(n_890), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_892), .B(n_893), .Y(n_891) );
NAND2x1p5_ASAP7_75t_L g895 ( .A(n_896), .B(n_905), .Y(n_895) );
NOR2x1_ASAP7_75t_L g896 ( .A(n_897), .B(n_902), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .Y(n_902) );
NOR2x1_ASAP7_75t_L g905 ( .A(n_906), .B(n_909), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_907), .B(n_908), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_910), .B(n_911), .Y(n_909) );
HB1xp67_ASAP7_75t_L g1033 ( .A(n_913), .Y(n_1033) );
XOR2x2_ASAP7_75t_L g914 ( .A(n_915), .B(n_928), .Y(n_914) );
NAND4xp75_ASAP7_75t_L g915 ( .A(n_916), .B(n_919), .C(n_923), .D(n_927), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_917), .B(n_918), .Y(n_916) );
AND2x2_ASAP7_75t_L g919 ( .A(n_920), .B(n_921), .Y(n_919) );
AND2x2_ASAP7_75t_L g923 ( .A(n_924), .B(n_925), .Y(n_923) );
INVx2_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
NOR2xp33_ASAP7_75t_L g933 ( .A(n_934), .B(n_941), .Y(n_933) );
NAND4xp25_ASAP7_75t_SL g934 ( .A(n_935), .B(n_936), .C(n_939), .D(n_940), .Y(n_934) );
NAND4xp25_ASAP7_75t_SL g941 ( .A(n_942), .B(n_943), .C(n_945), .D(n_947), .Y(n_941) );
BUFx6f_ASAP7_75t_SL g948 ( .A(n_949), .Y(n_948) );
OAI22xp5_ASAP7_75t_L g953 ( .A1(n_954), .A2(n_955), .B1(n_985), .B2(n_1034), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
INVx2_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
AND3x2_ASAP7_75t_L g958 ( .A(n_959), .B(n_969), .C(n_979), .Y(n_958) );
NOR2xp33_ASAP7_75t_L g959 ( .A(n_960), .B(n_966), .Y(n_959) );
OAI221xp5_ASAP7_75t_L g960 ( .A1(n_961), .A2(n_962), .B1(n_963), .B2(n_964), .C(n_965), .Y(n_960) );
OAI222xp33_ASAP7_75t_L g1071 ( .A1(n_963), .A2(n_1072), .B1(n_1073), .B2(n_1074), .C1(n_1075), .C2(n_1076), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_967), .B(n_968), .Y(n_966) );
NOR2xp33_ASAP7_75t_L g969 ( .A(n_970), .B(n_975), .Y(n_969) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
INVx2_ASAP7_75t_L g1034 ( .A(n_985), .Y(n_1034) );
XNOR2x1_ASAP7_75t_L g985 ( .A(n_986), .B(n_1031), .Y(n_985) );
AO22x2_ASAP7_75t_L g986 ( .A1(n_987), .A2(n_1011), .B1(n_1029), .B2(n_1030), .Y(n_986) );
INVx1_ASAP7_75t_L g1029 ( .A(n_987), .Y(n_1029) );
INVx2_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_991), .B(n_1003), .Y(n_990) );
NOR3xp33_ASAP7_75t_L g991 ( .A(n_992), .B(n_995), .C(n_1000), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_993), .B(n_994), .Y(n_992) );
OAI22xp5_ASAP7_75t_L g995 ( .A1(n_996), .A2(n_997), .B1(n_998), .B2(n_999), .Y(n_995) );
NOR2xp33_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1007), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1006), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1010), .Y(n_1007) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1011), .Y(n_1030) );
XOR2x2_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1028), .Y(n_1011) );
NAND2x1p5_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1020), .Y(n_1012) );
NOR2x1_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1017), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1016), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1019), .Y(n_1017) );
NOR2x1_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1025), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1024), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1027), .Y(n_1025) );
INVx2_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
INVx2_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1041), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1087 ( .A(n_1038), .B(n_1042), .Y(n_1087) );
NOR2xp33_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1040), .Y(n_1038) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1040), .Y(n_1085) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1045), .Y(n_1043) );
CKINVDCx20_ASAP7_75t_R g1047 ( .A(n_1048), .Y(n_1047) );
OR2x2_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1053), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
NOR2xp33_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1052), .Y(n_1050) );
INVxp67_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
OAI21xp33_ASAP7_75t_L g1055 ( .A1(n_1056), .A2(n_1058), .B(n_1082), .Y(n_1055) );
INVx1_ASAP7_75t_SL g1056 ( .A(n_1057), .Y(n_1056) );
AND2x4_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1070), .Y(n_1059) );
NOR2x1_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1065), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1063), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1067), .Y(n_1065) );
NOR2x1_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1077), .Y(n_1070) );
INVx2_ASAP7_75t_L g1109 ( .A(n_1076), .Y(n_1109) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1081), .Y(n_1077) );
INVx2_ASAP7_75t_SL g1079 ( .A(n_1080), .Y(n_1079) );
CKINVDCx20_ASAP7_75t_R g1083 ( .A(n_1084), .Y(n_1083) );
CKINVDCx6p67_ASAP7_75t_R g1086 ( .A(n_1087), .Y(n_1086) );
CKINVDCx5p33_ASAP7_75t_R g1088 ( .A(n_1089), .Y(n_1088) );
HB1xp67_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
NOR2xp67_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1102), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1096), .Y(n_1093) );
NOR3xp33_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1099), .C(n_1100), .Y(n_1096) );
NAND4xp25_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1106), .C(n_1107), .D(n_1108), .Y(n_1102) );
endmodule