module real_jpeg_11551_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_215;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

BUFx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_2),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_3),
.A2(n_76),
.B1(n_77),
.B2(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_3),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_3),
.A2(n_73),
.B(n_76),
.C(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_3),
.B(n_83),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_3),
.B(n_62),
.Y(n_201)
);

AOI21xp33_ASAP7_75t_SL g215 ( 
.A1(n_3),
.A2(n_62),
.B(n_201),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_3),
.B(n_30),
.C(n_50),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_145),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_3),
.B(n_89),
.Y(n_250)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_5),
.A2(n_76),
.B1(n_77),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_5),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_5),
.A2(n_62),
.B1(n_63),
.B2(n_134),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_134),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_5),
.A2(n_30),
.B1(n_34),
.B2(n_134),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_6),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_6),
.A2(n_47),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_6),
.A2(n_30),
.B1(n_34),
.B2(n_47),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_7),
.A2(n_56),
.B1(n_62),
.B2(n_63),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_7),
.A2(n_30),
.B1(n_34),
.B2(n_56),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_8),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_8),
.A2(n_33),
.B1(n_76),
.B2(n_77),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_8),
.A2(n_33),
.B1(n_44),
.B2(n_45),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_8),
.A2(n_33),
.B1(n_62),
.B2(n_63),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_11),
.A2(n_30),
.B1(n_34),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_11),
.A2(n_39),
.B1(n_62),
.B2(n_63),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_11),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_11),
.A2(n_39),
.B1(n_76),
.B2(n_77),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_12),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_13),
.A2(n_76),
.B1(n_77),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_13),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_13),
.A2(n_62),
.B1(n_63),
.B2(n_148),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_148),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_13),
.A2(n_30),
.B1(n_34),
.B2(n_148),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_14),
.A2(n_76),
.B1(n_77),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_14),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_14),
.A2(n_62),
.B1(n_63),
.B2(n_81),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_81),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_14),
.A2(n_30),
.B1(n_34),
.B2(n_81),
.Y(n_232)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_137),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_135),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_113),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_19),
.B(n_113),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_85),
.B2(n_112),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_57),
.C(n_70),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_22),
.A2(n_23),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_41),
.Y(n_267)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_35),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_27),
.A2(n_36),
.B(n_232),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_28),
.A2(n_123),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_28),
.A2(n_35),
.B(n_163),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_28),
.A2(n_162),
.B1(n_229),
.B2(n_231),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_29),
.A2(n_125),
.B(n_162),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_30),
.A2(n_34),
.B1(n_50),
.B2(n_51),
.Y(n_53)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_34),
.B(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_36),
.A2(n_37),
.B(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_36),
.A2(n_122),
.B(n_124),
.Y(n_121)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_36),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_36),
.A2(n_37),
.B1(n_230),
.B2(n_238),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_37),
.B(n_38),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_37),
.B(n_145),
.Y(n_236)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_48),
.B1(n_54),
.B2(n_55),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_43),
.A2(n_53),
.B(n_94),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_45),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_45),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_SL g202 ( 
.A(n_44),
.B(n_59),
.C(n_63),
.Y(n_202)
);

INVx5_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_45),
.A2(n_60),
.B(n_200),
.C(n_202),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_45),
.B(n_224),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_48),
.A2(n_55),
.B(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_48),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_48),
.A2(n_54),
.B1(n_196),
.B2(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_48),
.A2(n_54),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_48),
.A2(n_54),
.B1(n_217),
.B2(n_227),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_53),
.B(n_145),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_54),
.B(n_95),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_57),
.B(n_70),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_61),
.B(n_65),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_58),
.A2(n_67),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_58),
.A2(n_67),
.B1(n_151),
.B2(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_58),
.A2(n_67),
.B1(n_173),
.B2(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_68)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_61),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_63),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_62),
.A2(n_74),
.B(n_145),
.Y(n_166)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_87)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_67),
.A2(n_129),
.B(n_130),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_67),
.A2(n_152),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_69),
.B(n_89),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_80),
.B(n_82),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_109),
.B(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_71),
.A2(n_72),
.B1(n_80),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_71),
.A2(n_72),
.B1(n_133),
.B2(n_147),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_73),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_73),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_83),
.A2(n_143),
.B1(n_144),
.B2(n_146),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_97),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_91),
.B(n_96),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_87),
.B(n_91),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_89),
.B(n_180),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_92),
.A2(n_155),
.B(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_105),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_99),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_101),
.B1(n_102),
.B2(n_106),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_104),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.C(n_119),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_114),
.A2(n_115),
.B1(n_118),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_118),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_119),
.B(n_275),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_127),
.C(n_131),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_120),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_121),
.B(n_126),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_127),
.A2(n_128),
.B1(n_131),
.B2(n_132),
.Y(n_269)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_272),
.B(n_277),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_185),
.B(n_263),
.C(n_271),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_174),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_140),
.B(n_174),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_158),
.C(n_167),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_141),
.B(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_149),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_153),
.C(n_157),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_153),
.B1(n_154),
.B2(n_157),
.Y(n_149)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_159),
.B1(n_167),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_164),
.B2(n_165),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.C(n_172),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_193)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_172),
.B(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_182),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_175),
.B(n_183),
.C(n_184),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_181),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_177),
.B(n_178),
.C(n_181),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_261),
.B(n_262),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_205),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_188),
.B(n_191),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.C(n_197),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_194),
.A2(n_197),
.B1(n_198),
.B2(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_203),
.B1(n_204),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_218),
.B(n_260),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_207),
.B(n_210),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.C(n_216),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_211),
.B(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_216),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_254),
.B(n_259),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_244),
.B(n_253),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_233),
.B(n_243),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_228),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_228),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_225),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_239),
.B(n_242),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_241),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_246),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_249),
.C(n_252),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_251),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_258),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_270),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_270),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_267),
.C(n_268),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_274),
.Y(n_277)
);


endmodule