module fake_jpeg_4097_n_229 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_41),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_1),
.Y(n_39)
);

INVx2_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_31),
.Y(n_52)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx5_ASAP7_75t_SL g42 ( 
.A(n_37),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_41),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_49),
.Y(n_64)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_18),
.Y(n_49)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_54),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_30),
.Y(n_74)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_26),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_35),
.A2(n_32),
.B1(n_31),
.B2(n_23),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_23),
.B1(n_21),
.B2(n_18),
.Y(n_68)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_59),
.Y(n_91)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_61),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_63),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_48),
.A2(n_33),
.B1(n_35),
.B2(n_32),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_69),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_68),
.B(n_77),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_36),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_29),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_72),
.B(n_41),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_34),
.B(n_36),
.C(n_27),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_34),
.B1(n_38),
.B2(n_36),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_82),
.B1(n_20),
.B2(n_28),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_52),
.A2(n_32),
.B1(n_38),
.B2(n_29),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_20),
.B(n_26),
.C(n_24),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_38),
.B(n_41),
.C(n_30),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_78),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_50),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_44),
.A2(n_24),
.B1(n_21),
.B2(n_26),
.Y(n_82)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_85),
.A2(n_28),
.B1(n_25),
.B2(n_22),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_86),
.B(n_57),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_64),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_88),
.A2(n_89),
.B(n_94),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_26),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_73),
.B1(n_78),
.B2(n_57),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_20),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_72),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_76),
.Y(n_112)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_102),
.Y(n_117)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_80),
.B(n_47),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_108),
.A2(n_22),
.B(n_25),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_130),
.B(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_113),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_108),
.B(n_104),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_SL g151 ( 
.A1(n_111),
.A2(n_121),
.B(n_128),
.C(n_127),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_94),
.Y(n_139)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_71),
.Y(n_114)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_67),
.Y(n_115)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_118),
.A2(n_85),
.B1(n_84),
.B2(n_106),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_73),
.C(n_74),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_99),
.C(n_101),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_62),
.Y(n_121)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_122),
.B(n_123),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_58),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_128),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_1),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_125),
.B(n_131),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_28),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_92),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_69),
.B1(n_25),
.B2(n_22),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_129),
.A2(n_118),
.B1(n_130),
.B2(n_101),
.Y(n_138)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_2),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_2),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_133),
.A2(n_138),
.B1(n_144),
.B2(n_149),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_119),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_152),
.Y(n_161)
);

OAI321xp33_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_87),
.A3(n_97),
.B1(n_100),
.B2(n_92),
.C(n_108),
.Y(n_136)
);

OA21x2_ASAP7_75t_SL g156 ( 
.A1(n_136),
.A2(n_147),
.B(n_125),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_148),
.C(n_131),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_145),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_111),
.A2(n_84),
.B1(n_106),
.B2(n_102),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_115),
.A2(n_97),
.B1(n_86),
.B2(n_94),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_105),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_112),
.A2(n_116),
.B1(n_120),
.B2(n_111),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_109),
.B(n_117),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_122),
.B(n_110),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_151),
.A2(n_126),
.B(n_4),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_129),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_154)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_156),
.B(n_168),
.Y(n_176)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_159),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_172),
.C(n_143),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_113),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_163),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_147),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_126),
.B1(n_3),
.B2(n_4),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_164),
.A2(n_154),
.B1(n_138),
.B2(n_145),
.Y(n_188)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_169),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_135),
.B(n_140),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_171),
.A2(n_174),
.B(n_139),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_126),
.C(n_4),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_2),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_180),
.C(n_157),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_161),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_177),
.B(n_165),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_148),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_187),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_157),
.C(n_166),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_166),
.A2(n_151),
.B1(n_141),
.B2(n_143),
.Y(n_184)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_188),
.B(n_171),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_150),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_192),
.B1(n_196),
.B2(n_174),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_193),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_173),
.B(n_155),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_155),
.C(n_172),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_179),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_181),
.A2(n_173),
.B1(n_151),
.B2(n_165),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_197),
.B(n_199),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_183),
.B(n_174),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_204),
.Y(n_209)
);

NAND4xp25_ASAP7_75t_SL g202 ( 
.A(n_198),
.B(n_184),
.C(n_188),
.D(n_7),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_203),
.Y(n_211)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_191),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_192),
.B(n_193),
.Y(n_215)
);

BUFx24_ASAP7_75t_SL g206 ( 
.A(n_191),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_206),
.B(n_208),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_194),
.A2(n_176),
.B1(n_175),
.B2(n_178),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_207),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_187),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_210),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_189),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_214),
.A2(n_185),
.B(n_14),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_215),
.A2(n_190),
.B(n_196),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_216),
.A2(n_219),
.B(n_220),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_185),
.C(n_15),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_211),
.C(n_6),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_13),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g226 ( 
.A(n_222),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_213),
.B(n_8),
.C(n_9),
.Y(n_223)
);

AOI322xp5_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_224),
.A3(n_5),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_216),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_225),
.B(n_221),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_228),
.Y(n_229)
);

O2A1O1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_226),
.A2(n_11),
.B(n_5),
.C(n_9),
.Y(n_228)
);


endmodule