module real_jpeg_6600_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx5_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_0),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_0),
.Y(n_133)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_0),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_1),
.A2(n_27),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_1),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_1),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_1),
.A2(n_41),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_1),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_1),
.A2(n_154),
.B1(n_217),
.B2(n_220),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_1),
.A2(n_256),
.B(n_259),
.C(n_262),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_1),
.B(n_270),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_1),
.B(n_60),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_1),
.B(n_80),
.C(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_1),
.B(n_117),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_1),
.B(n_113),
.C(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_1),
.B(n_34),
.Y(n_330)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_2),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_3),
.A2(n_83),
.B1(n_86),
.B2(n_88),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_3),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_3),
.A2(n_88),
.B1(n_119),
.B2(n_123),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_3),
.A2(n_31),
.B1(n_88),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_3),
.A2(n_88),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_4),
.A2(n_15),
.B1(n_18),
.B2(n_20),
.Y(n_14)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_5),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_5),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_5),
.A2(n_94),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_5),
.A2(n_94),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_5),
.A2(n_94),
.B1(n_197),
.B2(n_201),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_6),
.Y(n_173)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_7),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_8),
.Y(n_169)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_8),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_8),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_8),
.Y(n_270)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_9),
.Y(n_258)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_12),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_12),
.A2(n_29),
.B1(n_146),
.B2(n_149),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_12),
.A2(n_29),
.B1(n_186),
.B2(n_190),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_12),
.A2(n_29),
.B1(n_167),
.B2(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_13),
.Y(n_80)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_13),
.Y(n_82)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_406),
.B(n_408),
.Y(n_20)
);

AO21x2_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_134),
.B(n_405),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_131),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_23),
.B(n_131),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_125),
.C(n_129),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_24),
.B(n_402),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_57),
.C(n_89),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_25),
.A2(n_180),
.B1(n_181),
.B2(n_192),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_25),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_25),
.B(n_141),
.C(n_181),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_25),
.B(n_237),
.C(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_25),
.A2(n_192),
.B1(n_237),
.B2(n_331),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_25),
.A2(n_192),
.B1(n_377),
.B2(n_378),
.Y(n_376)
);

OA22x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_33),
.B1(n_53),
.B2(n_56),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g225 ( 
.A1(n_26),
.A2(n_33),
.B1(n_53),
.B2(n_56),
.Y(n_225)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_33),
.A2(n_53),
.B1(n_56),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_33),
.A2(n_56),
.B1(n_126),
.B2(n_132),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_33),
.A2(n_53),
.B(n_56),
.Y(n_232)
);

AO21x1_ASAP7_75t_L g407 ( 
.A1(n_33),
.A2(n_56),
.B(n_132),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_43),
.Y(n_33)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_35),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_36),
.Y(n_184)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_37),
.Y(n_122)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_41),
.Y(n_261)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_49),
.B2(n_51),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_50),
.Y(n_127)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_57),
.A2(n_89),
.B1(n_379),
.B2(n_380),
.Y(n_378)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_57),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_57),
.B(n_225),
.C(n_382),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_57),
.A2(n_380),
.B1(n_382),
.B2(n_389),
.Y(n_388)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_85),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_58),
.B(n_151),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_73),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_59),
.A2(n_73),
.B1(n_144),
.B2(n_150),
.Y(n_143)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_60),
.A2(n_196),
.B(n_202),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_60),
.B(n_145),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_60),
.A2(n_74),
.B1(n_85),
.B2(n_196),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_64),
.B1(n_67),
.B2(n_71),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_65),
.Y(n_168)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx8_ASAP7_75t_L g163 ( 
.A(n_66),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_66),
.Y(n_219)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_70),
.Y(n_175)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_74),
.B(n_151),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_79),
.B1(n_81),
.B2(n_83),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_77),
.Y(n_153)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_77),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_77),
.Y(n_294)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_87),
.Y(n_201)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_89),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_96),
.B1(n_117),
.B2(n_118),
.Y(n_89)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_90),
.Y(n_383)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_93),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_96),
.B(n_224),
.Y(n_384)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_97),
.B(n_108),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g181 ( 
.A1(n_97),
.A2(n_108),
.B1(n_182),
.B2(n_185),
.Y(n_181)
);

OA22x2_ASAP7_75t_L g237 ( 
.A1(n_97),
.A2(n_108),
.B1(n_182),
.B2(n_185),
.Y(n_237)
);

NAND2x1_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_108),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_103),
.B1(n_105),
.B2(n_107),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_104),
.Y(n_313)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_108),
.A2(n_383),
.B(n_384),
.Y(n_382)
);

AOI22x1_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_113),
.B2(n_115),
.Y(n_108)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx8_ASAP7_75t_L g315 ( 
.A(n_111),
.Y(n_315)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_122),
.Y(n_189)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_125),
.B(n_129),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_130),
.B(n_224),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_131),
.B(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_131),
.B(n_407),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_400),
.B(n_404),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_371),
.B(n_397),
.Y(n_135)
);

OAI211xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_271),
.B(n_365),
.C(n_370),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_242),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g365 ( 
.A1(n_138),
.A2(n_242),
.B(n_366),
.C(n_369),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_226),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g370 ( 
.A(n_139),
.B(n_226),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_193),
.C(n_209),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_140),
.B(n_193),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_179),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_159),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_142),
.A2(n_143),
.B1(n_159),
.B2(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_142),
.A2(n_143),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_142),
.A2(n_143),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_143),
.B(n_266),
.C(n_303),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_143),
.B(n_323),
.C(n_325),
.Y(n_336)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx5_ASAP7_75t_SL g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_159),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_165),
.B1(n_170),
.B2(n_176),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_161),
.A2(n_213),
.B(n_214),
.Y(n_212)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_162),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_165),
.B(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_166),
.A2(n_216),
.B1(n_267),
.B2(n_270),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_166),
.A2(n_216),
.B1(n_267),
.B2(n_285),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_167),
.Y(n_282)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_205),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_173),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_173),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_178),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_180),
.A2(n_181),
.B1(n_221),
.B2(n_292),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_180),
.B(n_292),
.C(n_310),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_180),
.A2(n_181),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_181),
.B(n_225),
.C(n_341),
.Y(n_358)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_183),
.A2(n_257),
.B(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_204),
.B2(n_208),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_204),
.Y(n_233)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_SL g221 ( 
.A(n_203),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_204),
.A2(n_208),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_204),
.A2(n_232),
.B(n_233),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_205),
.B(n_216),
.Y(n_316)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_206),
.Y(n_285)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_223),
.C(n_225),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_221),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_212),
.A2(n_221),
.B1(n_292),
.B2(n_357),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_212),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_219),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_221),
.A2(n_292),
.B1(n_293),
.B2(n_297),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_221),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_223),
.A2(n_225),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_225),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_225),
.A2(n_249),
.B1(n_339),
.B2(n_340),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_225),
.A2(n_249),
.B1(n_375),
.B2(n_376),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_225),
.A2(n_249),
.B1(n_387),
.B2(n_388),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_225),
.B(n_376),
.C(n_381),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_240),
.B2(n_241),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_234),
.B1(n_235),
.B2(n_239),
.Y(n_228)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_229),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_234),
.B(n_239),
.C(n_241),
.Y(n_396)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B(n_238),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_237),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_237),
.A2(n_327),
.B1(n_328),
.B2(n_331),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_237),
.Y(n_331)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_238),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_238),
.A2(n_386),
.B1(n_390),
.B2(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_240),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_243),
.B(n_245),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_251),
.C(n_253),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_247),
.B(n_251),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_253),
.B(n_364),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_254),
.B(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_265),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_255),
.A2(n_265),
.B1(n_266),
.B2(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_255),
.Y(n_348)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_265),
.A2(n_266),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_266),
.B(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_287),
.Y(n_288)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_350),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_335),
.B(n_349),
.Y(n_272)
);

AOI21x1_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_320),
.B(n_334),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_307),
.B(n_319),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_299),
.B(n_306),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_289),
.B(n_298),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_286),
.B(n_288),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_284),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_284),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_284),
.A2(n_290),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_291),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_290),
.B(n_329),
.C(n_331),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_297),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_293),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_305),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_305),
.Y(n_306)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_303),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_309),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_318),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_316),
.B2(n_317),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_317),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_316),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_333),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_333),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_325),
.B1(n_326),
.B2(n_332),
.Y(n_321)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_322),
.Y(n_332)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_330),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_336),
.B(n_337),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_343),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_345),
.C(n_346),
.Y(n_359)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_341),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_344),
.A2(n_345),
.B1(n_346),
.B2(n_347),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

NOR2x1_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_360),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_352),
.B(n_359),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_359),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_355),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_353),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_358),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_356),
.B(n_358),
.C(n_362),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_360),
.A2(n_367),
.B(n_368),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_361),
.B(n_363),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_392),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_372),
.A2(n_398),
.B(n_399),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_385),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_373),
.B(n_385),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_381),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_382),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_390),
.C(n_391),
.Y(n_385)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_386),
.Y(n_395)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_391),
.B(n_394),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_393),
.B(n_396),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_393),
.B(n_396),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_403),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_401),
.B(n_403),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_409),
.Y(n_408)
);


endmodule