module fake_jpeg_10199_n_327 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_20),
.B(n_33),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_32),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_42),
.B(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_0),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_51),
.Y(n_74)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_27),
.B1(n_34),
.B2(n_19),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_22),
.B1(n_57),
.B2(n_31),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_28),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_66),
.Y(n_102)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_39),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_27),
.B1(n_34),
.B2(n_17),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_57),
.A2(n_61),
.B1(n_70),
.B2(n_23),
.Y(n_105)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_27),
.B1(n_34),
.B2(n_17),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_62),
.B1(n_21),
.B2(n_39),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_17),
.B1(n_26),
.B2(n_32),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_32),
.B1(n_18),
.B2(n_21),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_65),
.B(n_31),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_31),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_72),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_29),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_41),
.A2(n_33),
.B1(n_20),
.B2(n_18),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_69),
.B(n_41),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_73),
.B(n_106),
.C(n_46),
.Y(n_122)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_75),
.A2(n_81),
.B1(n_91),
.B2(n_108),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_21),
.B1(n_19),
.B2(n_22),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_77),
.A2(n_96),
.B1(n_99),
.B2(n_23),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_29),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_84),
.Y(n_114)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_16),
.C(n_15),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_SL g117 ( 
.A(n_85),
.B(n_101),
.C(n_107),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_87),
.Y(n_118)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_89),
.B(n_105),
.Y(n_123)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_60),
.Y(n_93)
);

AO22x2_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_46),
.B1(n_44),
.B2(n_43),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_94),
.A2(n_46),
.B1(n_43),
.B2(n_47),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_28),
.B1(n_25),
.B2(n_23),
.Y(n_96)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_98),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_72),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_61),
.A2(n_30),
.B1(n_20),
.B2(n_33),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_103),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_54),
.B(n_15),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_104),
.B(n_25),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_46),
.C(n_40),
.Y(n_106)
);

AND2x4_ASAP7_75t_L g107 ( 
.A(n_52),
.B(n_46),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_54),
.B(n_0),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_0),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_111),
.B(n_89),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_54),
.B1(n_50),
.B2(n_47),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_128),
.B1(n_50),
.B2(n_75),
.Y(n_141)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_130),
.Y(n_158)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_16),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_121),
.A2(n_104),
.B(n_82),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_106),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_102),
.B(n_44),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_131),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_SL g155 ( 
.A1(n_126),
.A2(n_117),
.B(n_135),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_46),
.C(n_43),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_71),
.C(n_49),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_94),
.A2(n_50),
.B1(n_47),
.B2(n_44),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_84),
.A2(n_94),
.B1(n_107),
.B2(n_86),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_88),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_44),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_25),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_133),
.B(n_134),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_73),
.B(n_1),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_135),
.A2(n_109),
.B(n_101),
.Y(n_143)
);

OR2x2_ASAP7_75t_SL g136 ( 
.A(n_80),
.B(n_35),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_136),
.A2(n_28),
.B(n_35),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_114),
.B(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_140),
.B(n_151),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_141),
.A2(n_144),
.B1(n_157),
.B2(n_138),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_107),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_152),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_136),
.B(n_126),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_145),
.B(n_161),
.C(n_162),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_105),
.B1(n_101),
.B2(n_107),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_146),
.A2(n_149),
.B1(n_154),
.B2(n_111),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_153),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_148),
.A2(n_156),
.B(n_126),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_123),
.A2(n_99),
.B1(n_107),
.B2(n_80),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_109),
.B(n_100),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_150),
.A2(n_155),
.B(n_167),
.Y(n_172)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_131),
.B(n_87),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_114),
.A2(n_40),
.B(n_92),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_137),
.B1(n_121),
.B2(n_112),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_75),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_160),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_97),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_92),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_97),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_165),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_113),
.B(n_76),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_91),
.C(n_90),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_171),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_119),
.B(n_35),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_132),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_76),
.Y(n_170)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_135),
.B(n_30),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_158),
.B(n_133),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_173),
.B(n_180),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g174 ( 
.A(n_164),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_179),
.Y(n_206)
);

O2A1O1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_121),
.B(n_119),
.C(n_137),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_175),
.A2(n_151),
.B1(n_148),
.B2(n_154),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_177),
.B(n_182),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_178),
.A2(n_141),
.B1(n_144),
.B2(n_176),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_147),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_165),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_168),
.A2(n_137),
.B1(n_120),
.B2(n_117),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_181),
.A2(n_193),
.B1(n_196),
.B2(n_149),
.Y(n_216)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_189),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_150),
.A2(n_132),
.B(n_137),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_186),
.B(n_192),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_194),
.Y(n_209)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_140),
.A2(n_138),
.B(n_134),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_116),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_198),
.C(n_201),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_SL g196 ( 
.A1(n_154),
.A2(n_116),
.B(n_110),
.C(n_30),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_158),
.B(n_164),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_202),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_143),
.A2(n_30),
.B(n_20),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_33),
.B(n_2),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_153),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_204),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_217),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_190),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_208),
.B(n_211),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_200),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_212),
.B(n_215),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_213),
.A2(n_221),
.B1(n_226),
.B2(n_182),
.Y(n_239)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_214),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_200),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_196),
.B1(n_198),
.B2(n_183),
.Y(n_238)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_145),
.C(n_139),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_222),
.C(n_185),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_175),
.A2(n_181),
.B1(n_196),
.B2(n_204),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_145),
.C(n_139),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_142),
.Y(n_223)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_224),
.A2(n_228),
.B1(n_171),
.B2(n_172),
.Y(n_244)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_187),
.Y(n_225)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_196),
.A2(n_145),
.B1(n_142),
.B2(n_171),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_178),
.A2(n_161),
.B1(n_167),
.B2(n_95),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_231),
.B(n_183),
.Y(n_232)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

NOR3xp33_ASAP7_75t_SL g234 ( 
.A(n_213),
.B(n_188),
.C(n_211),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_239),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_221),
.A2(n_216),
.B1(n_209),
.B2(n_219),
.Y(n_235)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_235),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_185),
.Y(n_236)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_236),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_218),
.Y(n_237)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_237),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_238),
.A2(n_240),
.B1(n_244),
.B2(n_246),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_226),
.A2(n_196),
.B1(n_186),
.B2(n_203),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_243),
.B(n_250),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_172),
.B1(n_195),
.B2(n_192),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_223),
.A2(n_201),
.B(n_177),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_205),
.B(n_229),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_227),
.B1(n_217),
.B2(n_225),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_249),
.A2(n_253),
.B1(n_214),
.B2(n_230),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_169),
.C(n_71),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_210),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_207),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_219),
.A2(n_210),
.B1(n_222),
.B2(n_205),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_256),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_265),
.B(n_268),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_258),
.A2(n_264),
.B1(n_272),
.B2(n_240),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_261),
.Y(n_274)
);

AOI31xp67_ASAP7_75t_L g261 ( 
.A1(n_234),
.A2(n_230),
.A3(n_212),
.B(n_206),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_235),
.A2(n_108),
.B(n_2),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_12),
.Y(n_284)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_246),
.B(n_1),
.CI(n_2),
.CON(n_263),
.SN(n_263)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_263),
.B(n_267),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_249),
.A2(n_95),
.B1(n_78),
.B2(n_49),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_3),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_242),
.A2(n_78),
.B1(n_10),
.B2(n_11),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_14),
.B(n_9),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_244),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_253),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_282),
.C(n_283),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_284),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_259),
.B(n_232),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_285),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_269),
.A2(n_247),
.B(n_245),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_280),
.A2(n_262),
.B(n_264),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_270),
.A2(n_233),
.B1(n_254),
.B2(n_241),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_281),
.A2(n_255),
.B1(n_272),
.B2(n_241),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_243),
.C(n_250),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_236),
.C(n_247),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_271),
.B(n_251),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g287 ( 
.A(n_261),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_263),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_255),
.B(n_239),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_248),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_290),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_274),
.A2(n_260),
.B(n_257),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_282),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_295),
.B(n_301),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_276),
.A2(n_254),
.B(n_277),
.Y(n_296)
);

OAI21x1_ASAP7_75t_SL g305 ( 
.A1(n_296),
.A2(n_297),
.B(n_300),
.Y(n_305)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_273),
.C(n_263),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_281),
.A2(n_256),
.B1(n_268),
.B2(n_265),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_303)
);

NOR2xp67_ASAP7_75t_SL g300 ( 
.A(n_283),
.B(n_10),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_278),
.A2(n_286),
.B(n_288),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_303),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_301),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_306),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_3),
.Y(n_307)
);

A2O1A1Ixp33_ASAP7_75t_L g318 ( 
.A1(n_307),
.A2(n_309),
.B(n_311),
.C(n_5),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_4),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_296),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_4),
.Y(n_309)
);

OAI21x1_ASAP7_75t_L g311 ( 
.A1(n_297),
.A2(n_5),
.B(n_6),
.Y(n_311)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_312),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_289),
.C(n_293),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_6),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_317),
.A3(n_304),
.B1(n_293),
.B2(n_316),
.C1(n_308),
.C2(n_314),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_310),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_6),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_321),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_317),
.C(n_7),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_324),
.A2(n_322),
.B(n_7),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_323),
.B(n_7),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_7),
.Y(n_327)
);


endmodule