module fake_jpeg_27562_n_80 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_80);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_80;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_4),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_11),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_2),
.B(n_10),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_0),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_24),
.A2(n_14),
.B1(n_6),
.B2(n_8),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_35),
.A2(n_36),
.B1(n_44),
.B2(n_28),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_2),
.B1(n_8),
.B2(n_9),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_39),
.Y(n_50)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_9),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_10),
.C(n_13),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

OR2x2_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_45),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_16),
.A2(n_13),
.B1(n_20),
.B2(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_20),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_57),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_44),
.B1(n_38),
.B2(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_22),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_54),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_48),
.B1(n_39),
.B2(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_32),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_62),
.C(n_51),
.Y(n_66)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_68),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_51),
.C(n_50),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_70),
.B(n_65),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_73),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_66),
.A2(n_64),
.B(n_63),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_68),
.C(n_59),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_58),
.C(n_49),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_62),
.B(n_58),
.Y(n_76)
);

AOI322xp5_ASAP7_75t_L g78 ( 
.A1(n_76),
.A2(n_77),
.A3(n_49),
.B1(n_61),
.B2(n_53),
.C1(n_23),
.C2(n_67),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_67),
.B1(n_61),
.B2(n_46),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_23),
.Y(n_80)
);


endmodule