module real_jpeg_6341_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g77 ( 
.A(n_0),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_1),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_1),
.Y(n_160)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_1),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_2),
.A2(n_175),
.B1(n_179),
.B2(n_180),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_2),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_3),
.A2(n_190),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_3),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_4),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_4),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_4),
.A2(n_93),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_4),
.A2(n_93),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_6),
.Y(n_157)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_6),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_6),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_6),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_7),
.A2(n_163),
.B1(n_168),
.B2(n_170),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_7),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_7),
.A2(n_170),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_8),
.Y(n_146)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_10),
.A2(n_46),
.B1(n_204),
.B2(n_205),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_10),
.B(n_246),
.C(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_10),
.B(n_71),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_10),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_10),
.B(n_240),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_10),
.B(n_139),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_12),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_12),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_12),
.A2(n_55),
.B1(n_117),
.B2(n_120),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_12),
.A2(n_55),
.B1(n_84),
.B2(n_90),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_12),
.A2(n_55),
.B1(n_168),
.B2(n_258),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_13),
.A2(n_108),
.B1(n_111),
.B2(n_114),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_13),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_13),
.A2(n_114),
.B1(n_189),
.B2(n_192),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_14),
.A2(n_41),
.B1(n_84),
.B2(n_87),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_14),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_87),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_14),
.A2(n_76),
.B1(n_87),
.B2(n_205),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_14),
.A2(n_87),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_15),
.Y(n_99)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_15),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_15),
.Y(n_246)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_230),
.B1(n_231),
.B2(n_342),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_18),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_229),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_197),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_20),
.B(n_197),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_134),
.C(n_181),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_21),
.B(n_339),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_59),
.B2(n_133),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_22),
.B(n_60),
.C(n_95),
.Y(n_214)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_43),
.B(n_52),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_24),
.B(n_54),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_25)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_29),
.Y(n_143)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_34),
.B(n_46),
.Y(n_196)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_36),
.Y(n_308)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_39),
.Y(n_142)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_46),
.B(n_47),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_48),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_46),
.A2(n_154),
.B(n_255),
.Y(n_274)
);

OAI21xp33_ASAP7_75t_SL g307 ( 
.A1(n_46),
.A2(n_308),
.B(n_309),
.Y(n_307)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_47),
.A2(n_138),
.A3(n_143),
.B1(n_144),
.B2(n_147),
.Y(n_137)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_58),
.Y(n_53)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_58),
.Y(n_227)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_95),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_83),
.B1(n_88),
.B2(n_89),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_61),
.Y(n_186)
);

OR2x2_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_71),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_65),
.B1(n_68),
.B2(n_69),
.Y(n_62)
);

INVx6_ASAP7_75t_L g323 ( 
.A(n_63),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_70),
.Y(n_151)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

AO22x2_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_75),
.B1(n_78),
.B2(n_80),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_74),
.Y(n_321)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g322 ( 
.A(n_76),
.B(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_77),
.Y(n_205)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_77),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g304 ( 
.A(n_77),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_79),
.Y(n_204)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_83),
.A2(n_88),
.B(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_86),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_88),
.B(n_185),
.Y(n_223)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_89),
.Y(n_222)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_107),
.B(n_115),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_96),
.A2(n_107),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_96),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_96),
.A2(n_115),
.B(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_96),
.A2(n_201),
.B1(n_265),
.B2(n_301),
.Y(n_300)
);

AOI22x1_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_100),
.B1(n_103),
.B2(n_104),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_101),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_102),
.Y(n_281)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_103),
.Y(n_248)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_123),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_116),
.B(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_117),
.Y(n_302)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_123),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_127),
.B1(n_130),
.B2(n_132),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_SL g320 ( 
.A(n_132),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_134),
.A2(n_135),
.B1(n_181),
.B2(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_152),
.B2(n_153),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_137),
.B(n_152),
.Y(n_218)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_145),
.B(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_149),
.Y(n_148)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_161),
.B1(n_171),
.B2(n_173),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_154),
.A2(n_251),
.B(n_255),
.Y(n_250)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_155),
.A2(n_162),
.B1(n_188),
.B2(n_194),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_155),
.A2(n_174),
.B1(n_207),
.B2(n_212),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_155),
.B(n_257),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_155),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_157),
.Y(n_273)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_157),
.Y(n_290)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx8_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_160),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_165),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_171),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_171),
.A2(n_277),
.B(n_282),
.Y(n_276)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_175),
.Y(n_278)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_180),
.B(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_181),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_187),
.C(n_196),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_182),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_186),
.A2(n_222),
.B(n_223),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_186),
.A2(n_223),
.B(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_187),
.B(n_196),
.Y(n_333)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_188),
.Y(n_313)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx8_ASAP7_75t_L g254 ( 
.A(n_191),
.Y(n_254)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_217),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_198)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_206),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_201),
.A2(n_238),
.B(n_239),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_201),
.A2(n_239),
.B(n_301),
.Y(n_330)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_224),
.B2(n_225),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B(n_228),
.Y(n_225)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

AOI21x1_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_336),
.B(n_341),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_325),
.B(n_335),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_295),
.B(n_324),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_268),
.B(n_294),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_249),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_236),
.B(n_249),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_241),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_237),
.A2(n_241),
.B1(n_242),
.B2(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_237),
.Y(n_292)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_262),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_250),
.B(n_263),
.C(n_267),
.Y(n_296)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_251),
.Y(n_288)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_285),
.B(n_293),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_275),
.B(n_284),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_274),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_283),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_283),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_277),
.Y(n_287)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_282),
.A2(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_291),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_291),
.Y(n_293)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_296),
.B(n_297),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_311),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_305),
.B2(n_306),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_305),
.C(n_311),
.Y(n_326)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

AOI32xp33_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_318),
.A3(n_320),
.B1(n_321),
.B2(n_322),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_317),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_312),
.B(n_317),
.Y(n_331)
);

INVx3_ASAP7_75t_SL g314 ( 
.A(n_315),
.Y(n_314)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx4_ASAP7_75t_SL g318 ( 
.A(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_326),
.B(n_327),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_332),
.B2(n_334),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_331),
.C(n_334),
.Y(n_337)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_332),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_337),
.B(n_338),
.Y(n_341)
);


endmodule