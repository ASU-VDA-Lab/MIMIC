module fake_jpeg_29216_n_543 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_543);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_543;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_378;
wire n_133;
wire n_419;
wire n_132;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_4),
.B(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_56),
.Y(n_136)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_57),
.Y(n_150)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_59),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_63),
.Y(n_151)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_65),
.Y(n_169)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_69),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_8),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_104),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_71),
.Y(n_157)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_76),
.Y(n_165)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_32),
.B(n_8),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_96),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_97),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_98),
.Y(n_172)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_100),
.Y(n_176)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

BUFx10_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_16),
.B(n_8),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_107),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_106),
.Y(n_116)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_33),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_109),
.Y(n_134)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_35),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_110),
.B(n_28),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_72),
.A2(n_47),
.B1(n_35),
.B2(n_51),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_114),
.A2(n_125),
.B1(n_137),
.B2(n_144),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_19),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_123),
.B(n_129),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_47),
.B1(n_35),
.B2(n_51),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_19),
.Y(n_129)
);

OR2x2_ASAP7_75t_SL g135 ( 
.A(n_91),
.B(n_51),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_135),
.B(n_174),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_56),
.A2(n_24),
.B1(n_50),
.B2(n_23),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_106),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_138),
.B(n_60),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_110),
.B(n_24),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_141),
.B(n_41),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_75),
.A2(n_47),
.B1(n_51),
.B2(n_35),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_59),
.A2(n_50),
.B1(n_18),
.B2(n_40),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_145),
.A2(n_146),
.B1(n_155),
.B2(n_171),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_107),
.A2(n_41),
.B1(n_38),
.B2(n_23),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_65),
.A2(n_16),
.B1(n_18),
.B2(n_40),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_69),
.A2(n_34),
.B1(n_29),
.B2(n_39),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_78),
.A2(n_34),
.B1(n_29),
.B2(n_39),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_175),
.B(n_45),
.Y(n_224)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_177),
.Y(n_252)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_112),
.Y(n_179)
);

INVx11_ASAP7_75t_L g263 ( 
.A(n_179),
.Y(n_263)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_180),
.Y(n_251)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_119),
.A2(n_86),
.B1(n_62),
.B2(n_68),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_183),
.A2(n_201),
.B1(n_204),
.B2(n_209),
.Y(n_240)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_127),
.Y(n_184)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_185),
.B(n_186),
.Y(n_233)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_128),
.Y(n_187)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_187),
.Y(n_253)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_130),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_188),
.B(n_196),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_71),
.B1(n_74),
.B2(n_98),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_189),
.A2(n_206),
.B1(n_217),
.B2(n_229),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_190),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_191),
.Y(n_243)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_192),
.Y(n_258)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_112),
.Y(n_193)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_193),
.Y(n_261)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_115),
.B(n_38),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_203),
.Y(n_241)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_131),
.Y(n_200)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_156),
.A2(n_57),
.B1(n_87),
.B2(n_95),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_133),
.Y(n_202)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_165),
.A2(n_87),
.B1(n_60),
.B2(n_97),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_111),
.B(n_26),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_208),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_L g206 ( 
.A1(n_121),
.A2(n_103),
.B1(n_100),
.B2(n_93),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_207),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_134),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_120),
.A2(n_27),
.B1(n_26),
.B2(n_28),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_124),
.B(n_36),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_215),
.Y(n_247)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_150),
.Y(n_211)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_211),
.Y(n_264)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_122),
.Y(n_212)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_212),
.Y(n_271)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_213),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_136),
.Y(n_214)
);

CKINVDCx6p67_ASAP7_75t_R g269 ( 
.A(n_214),
.Y(n_269)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_154),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_150),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_218),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_157),
.A2(n_36),
.B1(n_27),
.B2(n_45),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_133),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_113),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_219),
.B(n_220),
.Y(n_254)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_152),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_221),
.B(n_222),
.Y(n_267)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_172),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_223),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_225),
.Y(n_255)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_176),
.Y(n_225)
);

AND2x2_ASAP7_75t_SL g226 ( 
.A(n_139),
.B(n_164),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_228),
.C(n_31),
.Y(n_257)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_121),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_143),
.Y(n_238)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_139),
.B(n_0),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_157),
.A2(n_45),
.B1(n_31),
.B2(n_30),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_143),
.B(n_48),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_230),
.B(n_48),
.Y(n_245)
);

O2A1O1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_194),
.A2(n_146),
.B(n_171),
.C(n_161),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_231),
.A2(n_183),
.B(n_209),
.Y(n_274)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_238),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_194),
.A2(n_120),
.B1(n_159),
.B2(n_118),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_239),
.A2(n_180),
.B(n_211),
.Y(n_297)
);

XNOR2x1_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_257),
.Y(n_278)
);

AND2x2_ASAP7_75t_SL g248 ( 
.A(n_178),
.B(n_164),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_248),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_143),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_226),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_199),
.B(n_151),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_262),
.B(n_265),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_228),
.A2(n_31),
.B(n_30),
.C(n_114),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_195),
.B(n_10),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_268),
.B(n_14),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_262),
.A2(n_181),
.B1(n_189),
.B2(n_125),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_272),
.A2(n_276),
.B1(n_279),
.B2(n_292),
.Y(n_313)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_273),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_274),
.A2(n_284),
.B(n_297),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_275),
.B(n_277),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_240),
.A2(n_144),
.B1(n_229),
.B2(n_217),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_233),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_248),
.A2(n_201),
.B1(n_204),
.B2(n_228),
.Y(n_279)
);

OAI21xp33_ASAP7_75t_L g330 ( 
.A1(n_281),
.A2(n_299),
.B(n_267),
.Y(n_330)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_243),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_282),
.Y(n_312)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_243),
.Y(n_283)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_283),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_232),
.A2(n_190),
.B1(n_231),
.B2(n_167),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_254),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_254),
.Y(n_308)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_243),
.Y(n_287)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_287),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_248),
.B(n_226),
.C(n_198),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_290),
.C(n_256),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_245),
.B(n_207),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_291),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_218),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_255),
.B(n_202),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_248),
.A2(n_158),
.B1(n_152),
.B2(n_170),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_259),
.A2(n_206),
.B1(n_158),
.B2(n_126),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_293),
.A2(n_296),
.B1(n_269),
.B2(n_238),
.Y(n_310)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_294),
.Y(n_328)
);

OAI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_231),
.A2(n_167),
.B1(n_126),
.B2(n_220),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_295),
.A2(n_298),
.B1(n_302),
.B2(n_250),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_255),
.A2(n_170),
.B1(n_169),
.B2(n_214),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_241),
.A2(n_169),
.B1(n_191),
.B2(n_179),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_255),
.B(n_216),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_301),
.B(n_303),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_265),
.A2(n_163),
.B1(n_149),
.B2(n_147),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_255),
.B(n_30),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_241),
.B(n_48),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_304),
.B(n_265),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_305),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_274),
.A2(n_232),
.B1(n_270),
.B2(n_269),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_306),
.A2(n_264),
.B(n_283),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_308),
.B(n_316),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_309),
.B(n_315),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_310),
.A2(n_323),
.B1(n_333),
.B2(n_292),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_301),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_311),
.B(n_317),
.Y(n_347)
);

MAJx2_ASAP7_75t_L g315 ( 
.A(n_278),
.B(n_288),
.C(n_290),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_277),
.B(n_247),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_291),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_300),
.B(n_235),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_320),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_247),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_321),
.A2(n_284),
.B1(n_297),
.B2(n_286),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_280),
.A2(n_235),
.B1(n_246),
.B2(n_233),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_246),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_324),
.B(n_316),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_299),
.B(n_268),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_325),
.B(n_270),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_267),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_326),
.B(n_334),
.C(n_278),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_330),
.B(n_242),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_280),
.A2(n_250),
.B(n_271),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_332),
.A2(n_244),
.B(n_242),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_293),
.A2(n_252),
.B1(n_269),
.B2(n_244),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_290),
.B(n_237),
.C(n_266),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_335),
.A2(n_321),
.B1(n_317),
.B2(n_318),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_338),
.A2(n_339),
.B1(n_346),
.B2(n_358),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_313),
.A2(n_286),
.B1(n_272),
.B2(n_295),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_322),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_340),
.B(n_343),
.Y(n_371)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_342),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_319),
.B(n_289),
.Y(n_343)
);

AO21x2_ASAP7_75t_L g344 ( 
.A1(n_329),
.A2(n_269),
.B(n_302),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_344),
.A2(n_359),
.B1(n_306),
.B2(n_321),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_345),
.B(n_326),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_313),
.A2(n_279),
.B1(n_296),
.B2(n_281),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_315),
.B(n_303),
.C(n_298),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_348),
.B(n_309),
.C(n_334),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_324),
.B(n_276),
.Y(n_349)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_349),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_307),
.A2(n_269),
.B(n_271),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_350),
.A2(n_351),
.B(n_356),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_353),
.A2(n_327),
.B(n_314),
.Y(n_387)
);

XNOR2x1_ASAP7_75t_L g395 ( 
.A(n_354),
.B(n_270),
.Y(n_395)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_322),
.Y(n_355)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_355),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_305),
.A2(n_236),
.B(n_264),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_315),
.B(n_237),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_357),
.B(n_334),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_313),
.A2(n_252),
.B1(n_283),
.B2(n_282),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_310),
.A2(n_282),
.B1(n_287),
.B2(n_294),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_328),
.Y(n_360)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_360),
.Y(n_391)
);

A2O1A1Ixp33_ASAP7_75t_L g361 ( 
.A1(n_332),
.A2(n_260),
.B(n_236),
.C(n_266),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_361),
.B(n_362),
.Y(n_385)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_328),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_363),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_322),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_364),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_365),
.B(n_372),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_341),
.B(n_320),
.Y(n_367)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_367),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_326),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_373),
.B(n_381),
.C(n_344),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_374),
.A2(n_380),
.B1(n_393),
.B2(n_358),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_338),
.A2(n_333),
.B1(n_323),
.B2(n_311),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_377),
.A2(n_384),
.B1(n_390),
.B2(n_359),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_341),
.B(n_308),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_378),
.B(n_379),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_362),
.B(n_307),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_337),
.B(n_309),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_382),
.B(n_383),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_331),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_339),
.A2(n_329),
.B1(n_318),
.B2(n_327),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_387),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_357),
.B(n_331),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_388),
.B(n_392),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_342),
.B(n_325),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_389),
.B(n_352),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_346),
.A2(n_312),
.B1(n_314),
.B2(n_287),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_354),
.B(n_253),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_335),
.A2(n_312),
.B1(n_263),
.B2(n_273),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_253),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_394),
.B(n_395),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_397),
.A2(n_422),
.B1(n_376),
.B2(n_390),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_366),
.B(n_347),
.Y(n_398)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_398),
.Y(n_427)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_371),
.Y(n_399)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_399),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_368),
.B(n_336),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_401),
.B(n_406),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_402),
.B(n_410),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_366),
.B(n_347),
.Y(n_403)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_403),
.Y(n_434)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_391),
.Y(n_405)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_405),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_369),
.B(n_336),
.Y(n_406)
);

NOR3xp33_ASAP7_75t_L g407 ( 
.A(n_385),
.B(n_375),
.C(n_349),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_407),
.B(n_408),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_377),
.B(n_343),
.Y(n_408)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_409),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_388),
.B(n_351),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_370),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_411),
.B(n_413),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_394),
.B(n_383),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_384),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_414),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_387),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_415),
.A2(n_419),
.B1(n_355),
.B2(n_251),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_386),
.A2(n_356),
.B(n_350),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_417),
.B(n_421),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_373),
.B(n_361),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_393),
.B(n_360),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_374),
.A2(n_344),
.B1(n_353),
.B2(n_363),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_423),
.B(n_312),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_381),
.B(n_344),
.C(n_251),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_424),
.B(n_395),
.C(n_382),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_386),
.B(n_364),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_425),
.B(n_344),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_426),
.B(n_441),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_423),
.B(n_372),
.C(n_365),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_429),
.B(n_432),
.C(n_439),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_412),
.B(n_396),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_431),
.B(n_446),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_392),
.C(n_376),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_437),
.A2(n_447),
.B1(n_430),
.B2(n_438),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_438),
.B(n_400),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_396),
.B(n_344),
.C(n_340),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_416),
.B(n_312),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_440),
.B(n_403),
.Y(n_464)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_444),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_420),
.B(n_251),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_397),
.A2(n_263),
.B1(n_249),
.B2(n_234),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_420),
.B(n_263),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_448),
.B(n_416),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_441),
.B(n_424),
.C(n_414),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_451),
.B(n_460),
.C(n_464),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_436),
.A2(n_422),
.B1(n_400),
.B2(n_399),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_452),
.A2(n_464),
.B1(n_462),
.B2(n_456),
.Y(n_483)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_442),
.Y(n_453)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_453),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_435),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_454),
.B(n_455),
.Y(n_474)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_428),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_443),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_457),
.B(n_461),
.Y(n_485)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_427),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_SL g478 ( 
.A1(n_458),
.A2(n_467),
.B1(n_411),
.B2(n_418),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_462),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_429),
.B(n_432),
.C(n_426),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_449),
.B(n_404),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_434),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_463),
.B(n_405),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_431),
.B(n_402),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_448),
.C(n_446),
.Y(n_476)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_445),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_468),
.A2(n_439),
.B1(n_433),
.B2(n_425),
.Y(n_473)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_470),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_473),
.B(n_476),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_452),
.A2(n_430),
.B(n_437),
.Y(n_475)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_475),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_456),
.B(n_440),
.C(n_398),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_472),
.C(n_483),
.Y(n_494)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_478),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_466),
.A2(n_421),
.B1(n_417),
.B2(n_447),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_479),
.A2(n_481),
.B1(n_13),
.B2(n_12),
.Y(n_502)
);

NAND2x1p5_ASAP7_75t_L g480 ( 
.A(n_459),
.B(n_468),
.Y(n_480)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_480),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_451),
.A2(n_258),
.B1(n_249),
.B2(n_234),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_465),
.A2(n_213),
.B1(n_212),
.B2(n_132),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_483),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_450),
.A2(n_258),
.B(n_10),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_486),
.B(n_487),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_450),
.A2(n_9),
.B(n_13),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_487),
.B(n_460),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_488),
.B(n_492),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_485),
.B(n_469),
.Y(n_490)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_490),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_469),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_494),
.B(n_489),
.C(n_497),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_472),
.B(n_9),
.Y(n_496)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_496),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_471),
.B(n_122),
.C(n_48),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_476),
.C(n_471),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_473),
.B(n_13),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_498),
.B(n_502),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_474),
.B(n_48),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_503),
.B(n_484),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_494),
.A2(n_495),
.B(n_492),
.Y(n_505)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_505),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_499),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_508),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_501),
.Y(n_507)
);

NAND3xp33_ASAP7_75t_SL g525 ( 
.A(n_507),
.B(n_1),
.C(n_3),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_509),
.B(n_510),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_499),
.B(n_475),
.C(n_486),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_489),
.B(n_482),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_511),
.A2(n_493),
.B(n_1),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_500),
.A2(n_481),
.B1(n_480),
.B2(n_48),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_514),
.C(n_7),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_491),
.B(n_480),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_515),
.B(n_61),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_518),
.B(n_516),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_SL g521 ( 
.A1(n_507),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_521)
);

AOI21xp33_ASAP7_75t_L g531 ( 
.A1(n_521),
.A2(n_504),
.B(n_5),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_522),
.B(n_523),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_525),
.B(n_526),
.Y(n_530)
);

NOR2x1_ASAP7_75t_L g526 ( 
.A(n_512),
.B(n_1),
.Y(n_526)
);

AOI21xp33_ASAP7_75t_L g533 ( 
.A1(n_528),
.A2(n_531),
.B(n_525),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_520),
.B(n_517),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_529),
.A2(n_3),
.B(n_5),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_519),
.B(n_506),
.C(n_510),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_532),
.A2(n_524),
.B(n_508),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_533),
.B(n_536),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_534),
.B(n_535),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_527),
.A2(n_521),
.B(n_511),
.Y(n_535)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_538),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_539),
.A2(n_537),
.B(n_530),
.Y(n_540)
);

OAI211xp5_ASAP7_75t_L g541 ( 
.A1(n_540),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_3),
.C(n_5),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_542),
.A2(n_6),
.B1(n_7),
.B2(n_539),
.Y(n_543)
);


endmodule