module fake_jpeg_23222_n_236 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_30),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_33),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_1),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_28),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_49),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_18),
.B1(n_17),
.B2(n_16),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_41),
.A2(n_16),
.B1(n_21),
.B2(n_25),
.Y(n_76)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_30),
.B(n_24),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_30),
.Y(n_65)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_64),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_72),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_49),
.A2(n_18),
.B1(n_23),
.B2(n_17),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_67),
.B1(n_68),
.B2(n_76),
.Y(n_91)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_37),
.Y(n_85)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_69),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_18),
.B1(n_23),
.B2(n_17),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_50),
.A2(n_16),
.B1(n_23),
.B2(n_34),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_50),
.Y(n_69)
);

NAND2x1_ASAP7_75t_SL g70 ( 
.A(n_55),
.B(n_36),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_72),
.B(n_77),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_34),
.B1(n_31),
.B2(n_36),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_54),
.B1(n_52),
.B2(n_47),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_40),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_60),
.B(n_44),
.Y(n_78)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_65),
.B(n_44),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_84),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_SL g116 ( 
.A1(n_82),
.A2(n_75),
.B(n_58),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_46),
.B1(n_42),
.B2(n_45),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_87),
.B1(n_88),
.B2(n_90),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_59),
.B(n_32),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_89),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_33),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_33),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_37),
.B1(n_30),
.B2(n_32),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_37),
.B1(n_21),
.B2(n_25),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_48),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_56),
.A2(n_32),
.B1(n_14),
.B2(n_19),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_32),
.B1(n_15),
.B2(n_20),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_99),
.B1(n_64),
.B2(n_57),
.Y(n_106)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_97),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_96),
.A2(n_77),
.B(n_14),
.Y(n_111)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_56),
.A2(n_32),
.B1(n_14),
.B2(n_19),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_101),
.B(n_108),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_74),
.B(n_66),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_106),
.B1(n_122),
.B2(n_93),
.Y(n_130)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_104),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_100),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_107),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_111),
.A2(n_19),
.B(n_27),
.Y(n_126)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_81),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_58),
.B1(n_94),
.B2(n_97),
.Y(n_138)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_85),
.B1(n_91),
.B2(n_79),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_33),
.C(n_28),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_118),
.B(n_33),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_84),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_27),
.C(n_26),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_58),
.B1(n_75),
.B2(n_21),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_121),
.A2(n_89),
.B1(n_83),
.B2(n_87),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_123),
.A2(n_130),
.B1(n_101),
.B2(n_104),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_127),
.Y(n_145)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_121),
.B(n_85),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_142),
.C(n_115),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_141),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_138),
.B1(n_139),
.B2(n_122),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_79),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_111),
.A2(n_28),
.B(n_20),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_105),
.B(n_103),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_118),
.Y(n_155)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_144),
.B(n_149),
.Y(n_172)
);

AOI22x1_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_142),
.B1(n_141),
.B2(n_138),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_146),
.A2(n_162),
.B1(n_163),
.B2(n_135),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_147),
.A2(n_148),
.B(n_150),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_123),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_152),
.A2(n_156),
.B1(n_160),
.B2(n_161),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_124),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_153),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_142),
.Y(n_154)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_28),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_102),
.B1(n_109),
.B2(n_108),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_102),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_143),
.C(n_132),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_125),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_128),
.A2(n_114),
.B1(n_92),
.B2(n_62),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_173),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_167),
.C(n_174),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_140),
.C(n_92),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_146),
.B(n_126),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_171),
.B(n_175),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_151),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_155),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_62),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_178),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_20),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_20),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_175),
.A2(n_158),
.B1(n_145),
.B2(n_147),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_181),
.A2(n_190),
.B1(n_192),
.B2(n_6),
.Y(n_201)
);

NAND2xp33_ASAP7_75t_SL g183 ( 
.A(n_168),
.B(n_145),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_183),
.A2(n_174),
.B(n_176),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_171),
.A2(n_163),
.B1(n_161),
.B2(n_15),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_177),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_6),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_179),
.A2(n_15),
.B1(n_3),
.B2(n_4),
.Y(n_188)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_188),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_2),
.Y(n_189)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_169),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_170),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_192)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_167),
.C(n_166),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_184),
.C(n_180),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_172),
.Y(n_195)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_185),
.Y(n_196)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_203),
.B(n_180),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_182),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_200),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_5),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_8),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_199),
.A2(n_184),
.B1(n_187),
.B2(n_191),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_204),
.A2(n_196),
.B(n_201),
.Y(n_214)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_210),
.C(n_202),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_198),
.C(n_197),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_8),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_217),
.C(n_208),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_210),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_209),
.B(n_206),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_216),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_193),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_8),
.C(n_9),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_218),
.B(n_9),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_220),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_204),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_221),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_223),
.A2(n_224),
.B1(n_9),
.B2(n_10),
.Y(n_228)
);

OAI21x1_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_219),
.B(n_10),
.Y(n_225)
);

AOI21xp33_ASAP7_75t_L g230 ( 
.A1(n_225),
.A2(n_10),
.B(n_11),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_222),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_229),
.A2(n_230),
.B(n_226),
.Y(n_231)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_231),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_227),
.C(n_11),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_232),
.C(n_11),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_234),
.A2(n_13),
.B(n_203),
.Y(n_235)
);

BUFx24_ASAP7_75t_SL g236 ( 
.A(n_235),
.Y(n_236)
);


endmodule