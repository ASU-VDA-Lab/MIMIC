module fake_jpeg_15340_n_63 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_24;
wire n_38;
wire n_26;
wire n_28;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_0),
.B(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_42),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_21),
.A2(n_2),
.B(n_9),
.C(n_20),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_41),
.B(n_45),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_2),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_37),
.B1(n_32),
.B2(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_44),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_38),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_24),
.A2(n_27),
.B(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_23),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_22),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_46),
.B(n_49),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_54),
.A2(n_48),
.B1(n_50),
.B2(n_49),
.Y(n_55)
);

FAx1_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_48),
.CI(n_25),
.CON(n_58),
.SN(n_58)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_47),
.B1(n_28),
.B2(n_30),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_33),
.B(n_58),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_57),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

NOR3xp33_ASAP7_75t_SL g62 ( 
.A(n_61),
.B(n_58),
.C(n_60),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);


endmodule