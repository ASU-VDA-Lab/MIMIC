module fake_jpeg_4734_n_179 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_0),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_33),
.Y(n_41)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_27),
.B1(n_23),
.B2(n_26),
.Y(n_44)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_29),
.B(n_28),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_26),
.B1(n_24),
.B2(n_27),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_32),
.B1(n_22),
.B2(n_16),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_27),
.B1(n_15),
.B2(n_29),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_14),
.B1(n_20),
.B2(n_28),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_15),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_30),
.B(n_32),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_31),
.C(n_22),
.Y(n_57)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_50),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_38),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_58),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_61),
.Y(n_98)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_62),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_64),
.B1(n_21),
.B2(n_35),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_66),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_32),
.B1(n_35),
.B2(n_33),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_25),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_65),
.A2(n_73),
.B(n_21),
.Y(n_95)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_17),
.B1(n_19),
.B2(n_32),
.Y(n_82)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_72),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_14),
.C(n_20),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_12),
.B(n_2),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_17),
.Y(n_71)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_21),
.B(n_25),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_80),
.B(n_90),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_57),
.A2(n_37),
.B1(n_35),
.B2(n_33),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_37),
.B1(n_33),
.B2(n_36),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_37),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_94),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_95),
.B(n_61),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_51),
.A2(n_36),
.B1(n_2),
.B2(n_3),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_92),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_99),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_110),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_98),
.B(n_80),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_96),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_115),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_59),
.C(n_58),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_114),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_108),
.B(n_112),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_93),
.A2(n_90),
.B(n_78),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_109),
.A2(n_98),
.B(n_86),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_54),
.Y(n_111)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_70),
.C(n_67),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

HAxp5_ASAP7_75t_SL g127 ( 
.A(n_116),
.B(n_88),
.CON(n_127),
.SN(n_127)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_86),
.A2(n_52),
.B1(n_56),
.B2(n_75),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

NOR3xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_78),
.C(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_130),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_109),
.B(n_114),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_123),
.B(n_129),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_77),
.B1(n_68),
.B2(n_88),
.Y(n_126)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_127),
.A2(n_108),
.B1(n_100),
.B2(n_117),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_77),
.B1(n_79),
.B2(n_65),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_112),
.A2(n_72),
.B1(n_79),
.B2(n_89),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_116),
.A2(n_36),
.B1(n_89),
.B2(n_94),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_105),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_104),
.C(n_107),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_120),
.C(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_110),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_135),
.B(n_137),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_118),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_118),
.B(n_115),
.Y(n_138)
);

OA21x2_ASAP7_75t_SL g146 ( 
.A1(n_138),
.A2(n_140),
.B(n_129),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_103),
.B(n_105),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_145),
.B1(n_124),
.B2(n_132),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_128),
.B(n_99),
.Y(n_144)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_131),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_148),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_124),
.B1(n_125),
.B2(n_132),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_150),
.B1(n_1),
.B2(n_4),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_136),
.A2(n_125),
.B1(n_126),
.B2(n_120),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_152),
.C(n_141),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_81),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_157),
.B(n_161),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_142),
.Y(n_156)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_140),
.C(n_36),
.Y(n_157)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_1),
.C(n_4),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_1),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_162),
.A2(n_150),
.B(n_6),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_154),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_163),
.A2(n_164),
.B(n_168),
.Y(n_170)
);

NAND4xp25_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_146),
.C(n_154),
.D(n_152),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_160),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_171),
.C(n_172),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_167),
.B1(n_148),
.B2(n_155),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_5),
.C(n_6),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_5),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_173),
.A2(n_175),
.B(n_5),
.Y(n_176)
);

BUFx24_ASAP7_75t_SL g175 ( 
.A(n_171),
.Y(n_175)
);

AOI221xp5_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_177),
.B1(n_7),
.B2(n_9),
.C(n_10),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_174),
.A2(n_7),
.B(n_9),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_7),
.Y(n_179)
);


endmodule