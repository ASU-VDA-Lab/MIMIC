module fake_jpeg_4270_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_23),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_21),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_23),
.A2(n_9),
.B(n_10),
.C(n_16),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_0),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_10),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_25),
.A2(n_20),
.B1(n_19),
.B2(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_15),
.B1(n_17),
.B2(n_22),
.Y(n_36)
);

OAI22x1_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_29),
.B1(n_17),
.B2(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_19),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_35),
.B1(n_22),
.B2(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_26),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_30),
.B(n_29),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_30),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_21),
.C(n_1),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_51),
.B(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_24),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_1),
.Y(n_59)
);

XOR2x2_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_21),
.Y(n_54)
);

MAJx2_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_42),
.C(n_41),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_60),
.C(n_49),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_51),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_56),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_59),
.B1(n_52),
.B2(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_62),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_47),
.C(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_65),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_4),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_69),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_1),
.B1(n_5),
.B2(n_7),
.Y(n_69)
);

NOR2x1_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_66),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_71),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_7),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_8),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_73),
.Y(n_75)
);

AOI21x1_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_70),
.B(n_74),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_8),
.Y(n_77)
);


endmodule