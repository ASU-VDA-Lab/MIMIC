module fake_jpeg_22991_n_341 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_40),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_18),
.B(n_7),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_46),
.Y(n_51)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_54),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_36),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_59),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_36),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_38),
.Y(n_90)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_63),
.Y(n_73)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

CKINVDCx12_ASAP7_75t_R g66 ( 
.A(n_38),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_66),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_33),
.B1(n_34),
.B2(n_25),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_30),
.B1(n_32),
.B2(n_22),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_38),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_70),
.Y(n_99)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_56),
.B(n_30),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_87),
.Y(n_118)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_77),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_51),
.B(n_26),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_79),
.B(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_83),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_33),
.B1(n_34),
.B2(n_25),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_57),
.B1(n_58),
.B2(n_53),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_20),
.Y(n_85)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_31),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_93),
.Y(n_117)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_57),
.A2(n_19),
.B1(n_30),
.B2(n_22),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_45),
.B1(n_25),
.B2(n_24),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_96),
.B1(n_65),
.B2(n_53),
.Y(n_125)
);

AND2x4_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_39),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_39),
.B(n_61),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_57),
.A2(n_22),
.B1(n_32),
.B2(n_24),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_98),
.A2(n_32),
.B1(n_62),
.B2(n_39),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_51),
.B(n_50),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_55),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_54),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_65),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

NOR2x1_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_97),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_90),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_58),
.B1(n_24),
.B2(n_43),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_107),
.A2(n_112),
.B1(n_122),
.B2(n_125),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_115),
.B1(n_128),
.B2(n_130),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_39),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_84),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_96),
.B(n_97),
.C(n_87),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_116),
.B(n_120),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_72),
.B(n_61),
.Y(n_141)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_97),
.A2(n_58),
.B1(n_62),
.B2(n_26),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_75),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_124),
.B(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_81),
.A2(n_65),
.B1(n_70),
.B2(n_63),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_76),
.B(n_21),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_129),
.B(n_131),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_80),
.B(n_29),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_132),
.B(n_138),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_99),
.C(n_100),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_139),
.C(n_110),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_125),
.A2(n_72),
.B1(n_80),
.B2(n_88),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_135),
.A2(n_150),
.B1(n_151),
.B2(n_106),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_137),
.A2(n_141),
.B(n_146),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_99),
.C(n_93),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_84),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_131),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_142),
.B(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_92),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_147),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_92),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_153),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_120),
.A2(n_76),
.B1(n_78),
.B2(n_101),
.Y(n_151)
);

AO22x2_ASAP7_75t_L g152 ( 
.A1(n_115),
.A2(n_49),
.B1(n_47),
.B2(n_43),
.Y(n_152)
);

AO22x1_ASAP7_75t_SL g166 ( 
.A1(n_152),
.A2(n_49),
.B1(n_114),
.B2(n_107),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_104),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_154),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_78),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_157),
.Y(n_173)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_126),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_77),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_94),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_116),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_114),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_161),
.Y(n_196)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_162),
.A2(n_108),
.B1(n_121),
.B2(n_89),
.Y(n_168)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_167),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g209 ( 
.A1(n_166),
.A2(n_142),
.B(n_162),
.Y(n_209)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_152),
.A2(n_115),
.B1(n_128),
.B2(n_119),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_169),
.A2(n_31),
.B1(n_28),
.B2(n_133),
.Y(n_225)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_176),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_178),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_110),
.C(n_117),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_172),
.B(n_29),
.C(n_102),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_111),
.B1(n_117),
.B2(n_121),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_182),
.B1(n_188),
.B2(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_187),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_189),
.Y(n_218)
);

OAI22x1_ASAP7_75t_SL g182 ( 
.A1(n_152),
.A2(n_102),
.B1(n_47),
.B2(n_28),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_129),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_137),
.Y(n_203)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_132),
.B(n_106),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_190),
.B(n_192),
.Y(n_220)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_191),
.A2(n_193),
.B(n_195),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_83),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_143),
.A2(n_148),
.B1(n_149),
.B2(n_161),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_146),
.A2(n_23),
.B(n_21),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_163),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_200),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_180),
.A2(n_159),
.B1(n_137),
.B2(n_153),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_202),
.A2(n_213),
.B(n_224),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_214),
.C(n_222),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_165),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_205),
.B(n_206),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_163),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_174),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_207),
.B(n_211),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_212),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_177),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_183),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_SL g213 ( 
.A(n_185),
.B(n_173),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_158),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_173),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_221),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_181),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_219),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_178),
.B(n_171),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_35),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_195),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_184),
.B1(n_31),
.B2(n_28),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_35),
.C(n_31),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_196),
.C(n_169),
.Y(n_230)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_227),
.B(n_231),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_241),
.C(n_245),
.Y(n_264)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_218),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_208),
.A2(n_196),
.B(n_193),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_232),
.A2(n_249),
.B(n_250),
.Y(n_271)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_233),
.B(n_240),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_213),
.A2(n_189),
.B1(n_187),
.B2(n_166),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_225),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_221),
.A2(n_166),
.B1(n_167),
.B2(n_164),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_202),
.A2(n_172),
.B1(n_176),
.B2(n_184),
.Y(n_236)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_220),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_203),
.B(n_186),
.C(n_35),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_210),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_243)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_35),
.C(n_20),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_226),
.C(n_201),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_35),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_209),
.A2(n_0),
.B(n_1),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_199),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_222),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_251),
.B(n_198),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_234),
.B(n_223),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_255),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_197),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_256),
.A2(n_259),
.B1(n_273),
.B2(n_238),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_197),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_262),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_246),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_258),
.B(n_260),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_215),
.B1(n_209),
.B2(n_224),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_240),
.B(n_207),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_198),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_263),
.A2(n_266),
.B(n_271),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_242),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_265),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_SL g266 ( 
.A(n_239),
.B(n_215),
.C(n_206),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_268),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_201),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_233),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_261),
.A2(n_244),
.B1(n_236),
.B2(n_230),
.Y(n_276)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_272),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_278),
.Y(n_302)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_269),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_254),
.A2(n_242),
.B1(n_227),
.B2(n_250),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_281),
.A2(n_286),
.B1(n_289),
.B2(n_290),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_267),
.A2(n_235),
.B1(n_251),
.B2(n_229),
.Y(n_282)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_282),
.Y(n_296)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_273),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_284),
.A2(n_285),
.B(n_8),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_229),
.B1(n_232),
.B2(n_237),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_268),
.B(n_248),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_20),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_288),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_256),
.A2(n_259),
.B1(n_271),
.B2(n_264),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_262),
.A2(n_249),
.B1(n_243),
.B2(n_247),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_253),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_300),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_264),
.B1(n_252),
.B2(n_255),
.Y(n_293)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_293),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_257),
.C(n_241),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_305),
.C(n_279),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_297),
.Y(n_308)
);

INVx4_ASAP7_75t_SL g298 ( 
.A(n_280),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_298),
.A2(n_290),
.B1(n_279),
.B2(n_274),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_20),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_301),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_20),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_2),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_281),
.A2(n_7),
.B(n_15),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_304),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_1),
.C(n_2),
.Y(n_305)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_306),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_307),
.B(n_310),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_309),
.A2(n_12),
.B(n_14),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_294),
.A2(n_11),
.B1(n_15),
.B2(n_5),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_291),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_316),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_7),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_314),
.A2(n_318),
.B(n_302),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_295),
.B(n_11),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_11),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_319),
.B(n_323),
.Y(n_331)
);

OAI321xp33_ASAP7_75t_L g322 ( 
.A1(n_312),
.A2(n_299),
.A3(n_305),
.B1(n_293),
.B2(n_300),
.C(n_292),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_327),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_317),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_299),
.C(n_317),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_326),
.C(n_320),
.Y(n_334)
);

AOI31xp33_ASAP7_75t_L g327 ( 
.A1(n_312),
.A2(n_12),
.A3(n_14),
.B(n_16),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_325),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_329),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_324),
.A2(n_311),
.B(n_308),
.Y(n_329)
);

AOI21x1_ASAP7_75t_L g332 ( 
.A1(n_323),
.A2(n_14),
.B(n_16),
.Y(n_332)
);

O2A1O1Ixp33_ASAP7_75t_SL g336 ( 
.A1(n_332),
.A2(n_3),
.B(n_4),
.C(n_330),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_321),
.B(n_16),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_333),
.A2(n_334),
.B(n_3),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_336),
.A2(n_337),
.B(n_331),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_328),
.B1(n_335),
.B2(n_4),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_4),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_4),
.Y(n_341)
);


endmodule