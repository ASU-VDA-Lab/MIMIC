module fake_jpeg_2840_n_599 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_599);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_599;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_7),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_56),
.B(n_57),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_22),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_58),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_29),
.B(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_60),
.B(n_61),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_20),
.B(n_7),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_24),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_64),
.B(n_68),
.Y(n_141)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_24),
.B(n_51),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_73),
.Y(n_186)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_74),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_75),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_76),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_8),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_77),
.B(n_89),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_79),
.Y(n_172)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_82),
.Y(n_163)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_8),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_85),
.B(n_98),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_86),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_6),
.B1(n_15),
.B2(n_14),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_87),
.A2(n_19),
.B1(n_44),
.B2(n_40),
.Y(n_190)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_42),
.B(n_6),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_90),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_91),
.Y(n_145)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_92),
.Y(n_178)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_6),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_99),
.Y(n_189)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_46),
.Y(n_100)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g132 ( 
.A(n_102),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_103),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_48),
.B(n_6),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_29),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

INVx5_ASAP7_75t_SL g133 ( 
.A(n_107),
.Y(n_133)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_25),
.Y(n_109)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_110),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_38),
.Y(n_111)
);

NAND2xp33_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_38),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx5_ASAP7_75t_SL g140 ( 
.A(n_113),
.Y(n_140)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_114),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g115 ( 
.A(n_26),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_115),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_56),
.A2(n_85),
.B1(n_79),
.B2(n_96),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_116),
.A2(n_118),
.B1(n_160),
.B2(n_190),
.Y(n_222)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_117),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_63),
.A2(n_53),
.B1(n_50),
.B2(n_52),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_119),
.Y(n_200)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_120),
.Y(n_204)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_123),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_67),
.A2(n_51),
.B1(n_36),
.B2(n_44),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_129),
.A2(n_32),
.B1(n_30),
.B2(n_55),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_136),
.B(n_32),
.Y(n_216)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_147),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_153),
.B(n_188),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_69),
.A2(n_53),
.B1(n_50),
.B2(n_52),
.Y(n_160)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_72),
.Y(n_168)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_92),
.Y(n_169)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_169),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_99),
.B(n_109),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_171),
.B(n_52),
.Y(n_231)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_173),
.Y(n_242)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_86),
.Y(n_174)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_174),
.Y(n_251)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_179),
.Y(n_253)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_104),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_180),
.Y(n_246)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_59),
.B(n_36),
.Y(n_188)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_121),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_191),
.Y(n_263)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_121),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_193),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_130),
.A2(n_58),
.B1(n_113),
.B2(n_65),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_194),
.A2(n_230),
.B1(n_241),
.B2(n_257),
.Y(n_266)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_195),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_40),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_196),
.B(n_201),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_171),
.A2(n_19),
.B(n_115),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_197),
.Y(n_264)
);

AND2x2_ASAP7_75t_SL g199 ( 
.A(n_131),
.B(n_66),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g269 ( 
.A(n_199),
.B(n_232),
.C(n_235),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_141),
.B(n_73),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_143),
.A2(n_78),
.B1(n_76),
.B2(n_70),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_202),
.A2(n_249),
.B1(n_252),
.B2(n_30),
.Y(n_285)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_127),
.Y(n_206)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_206),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_124),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_207),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_134),
.B(n_33),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_208),
.B(n_227),
.Y(n_261)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_138),
.Y(n_209)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_209),
.Y(n_293)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_149),
.Y(n_210)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_210),
.Y(n_273)
);

INVx5_ASAP7_75t_SL g211 ( 
.A(n_133),
.Y(n_211)
);

INVx13_ASAP7_75t_L g289 ( 
.A(n_211),
.Y(n_289)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_146),
.Y(n_212)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_212),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_133),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_213),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_125),
.A2(n_75),
.B1(n_106),
.B2(n_32),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_215),
.B(n_216),
.Y(n_280)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_152),
.Y(n_219)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_219),
.Y(n_283)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_157),
.Y(n_220)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_220),
.Y(n_307)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_149),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_221),
.Y(n_284)
);

O2A1O1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_140),
.A2(n_107),
.B(n_80),
.C(n_115),
.Y(n_223)
);

OA22x2_ASAP7_75t_L g308 ( 
.A1(n_223),
.A2(n_236),
.B1(n_26),
.B2(n_140),
.Y(n_308)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_162),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_224),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_183),
.Y(n_225)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_225),
.Y(n_282)
);

AO22x1_ASAP7_75t_SL g226 ( 
.A1(n_184),
.A2(n_90),
.B1(n_102),
.B2(n_101),
.Y(n_226)
);

AO22x1_ASAP7_75t_L g305 ( 
.A1(n_226),
.A2(n_182),
.B1(n_37),
.B2(n_28),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_145),
.B(n_151),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_156),
.B(n_27),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_228),
.B(n_238),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_132),
.A2(n_97),
.B1(n_108),
.B2(n_74),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_229),
.A2(n_139),
.B1(n_159),
.B2(n_176),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_126),
.A2(n_46),
.B1(n_50),
.B2(n_52),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_231),
.B(n_235),
.Y(n_310)
);

AND2x2_ASAP7_75t_SL g232 ( 
.A(n_177),
.B(n_66),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_178),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_233),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_122),
.Y(n_234)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_234),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_152),
.B(n_59),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_132),
.A2(n_17),
.B1(n_55),
.B2(n_41),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_163),
.B(n_33),
.Y(n_238)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_167),
.Y(n_240)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_240),
.Y(n_295)
);

INVx11_ASAP7_75t_L g241 ( 
.A(n_149),
.Y(n_241)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_178),
.Y(n_243)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_243),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_122),
.Y(n_244)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_244),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_135),
.Y(n_245)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_245),
.Y(n_317)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_247),
.Y(n_318)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_189),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_250),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_183),
.B(n_27),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_158),
.A2(n_52),
.B1(n_50),
.B2(n_46),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_166),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_254),
.Y(n_291)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_164),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_258),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_150),
.B(n_41),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_256),
.B(n_139),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_166),
.A2(n_114),
.B1(n_30),
.B2(n_26),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_167),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_186),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_128),
.Y(n_268)
);

INVx8_ASAP7_75t_L g260 ( 
.A(n_135),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_260),
.A2(n_225),
.B1(n_241),
.B2(n_259),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_268),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_269),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_216),
.B(n_172),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_270),
.B(n_298),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_271),
.A2(n_285),
.B1(n_297),
.B2(n_305),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_203),
.B(n_186),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_275),
.B(n_299),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_192),
.B(n_199),
.C(n_237),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_277),
.B(n_232),
.C(n_200),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_279),
.B(n_296),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_197),
.A2(n_172),
.B1(n_154),
.B2(n_175),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_281),
.A2(n_304),
.B1(n_243),
.B2(n_248),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_290),
.A2(n_292),
.B1(n_303),
.B2(n_315),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_226),
.A2(n_175),
.B1(n_170),
.B2(n_165),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_213),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_222),
.A2(n_159),
.B1(n_176),
.B2(n_158),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_199),
.B(n_170),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_251),
.B(n_128),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_242),
.B(n_142),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_300),
.B(n_301),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_217),
.B(n_142),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_202),
.B(n_154),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_302),
.B(n_309),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_246),
.A2(n_155),
.B1(n_144),
.B2(n_182),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_222),
.A2(n_165),
.B1(n_155),
.B2(n_144),
.Y(n_304)
);

OA21x2_ASAP7_75t_L g335 ( 
.A1(n_308),
.A2(n_223),
.B(n_229),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_218),
.B(n_14),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_232),
.B(n_0),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_312),
.B(n_240),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_239),
.B(n_204),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_313),
.B(n_211),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_246),
.A2(n_148),
.B1(n_18),
.B2(n_28),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_230),
.A2(n_37),
.B1(n_28),
.B2(n_18),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_316),
.A2(n_260),
.B1(n_234),
.B2(n_245),
.Y(n_344)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_282),
.Y(n_320)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_320),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_272),
.B(n_261),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_321),
.B(n_323),
.C(n_326),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_265),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_324),
.B(n_318),
.Y(n_390)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_282),
.Y(n_325)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_325),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_277),
.B(n_214),
.C(n_255),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_272),
.B(n_253),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_327),
.B(n_348),
.Y(n_389)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_276),
.Y(n_330)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_330),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_331),
.B(n_351),
.Y(n_381)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_276),
.Y(n_332)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_332),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_302),
.A2(n_215),
.B1(n_226),
.B2(n_194),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_334),
.A2(n_344),
.B1(n_347),
.B2(n_316),
.Y(n_370)
);

OAI31xp33_ASAP7_75t_L g410 ( 
.A1(n_335),
.A2(n_289),
.A3(n_273),
.B(n_284),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_285),
.A2(n_264),
.B1(n_280),
.B2(n_297),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_336),
.A2(n_341),
.B1(n_342),
.B2(n_352),
.Y(n_387)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_295),
.Y(n_338)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_338),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_264),
.A2(n_236),
.B1(n_191),
.B2(n_193),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_286),
.Y(n_345)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_345),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_286),
.Y(n_346)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_346),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_280),
.A2(n_195),
.B1(n_257),
.B2(n_198),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_274),
.B(n_205),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_349),
.B(n_350),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_274),
.B(n_224),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_261),
.B(n_219),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_305),
.A2(n_244),
.B1(n_254),
.B2(n_221),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_305),
.A2(n_210),
.B1(n_37),
.B2(n_28),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_353),
.A2(n_362),
.B1(n_266),
.B2(n_291),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_287),
.A2(n_37),
.B1(n_28),
.B2(n_18),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_354),
.A2(n_271),
.B1(n_334),
.B2(n_347),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_279),
.B(n_0),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_355),
.B(n_365),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_295),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_356),
.Y(n_379)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_314),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_357),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_269),
.B(n_37),
.C(n_28),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_361),
.C(n_269),
.Y(n_378)
);

AND2x2_ASAP7_75t_SL g360 ( 
.A(n_310),
.B(n_312),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_364),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_SL g361 ( 
.A(n_280),
.B(n_37),
.C(n_34),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_298),
.A2(n_34),
.B1(n_31),
.B2(n_10),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_262),
.B(n_10),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_363),
.B(n_291),
.Y(n_397)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_311),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_287),
.B(n_0),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_311),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_366),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_296),
.B(n_1),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_367),
.B(n_368),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_309),
.B(n_1),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_369),
.A2(n_337),
.B1(n_341),
.B2(n_359),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_370),
.A2(n_335),
.B1(n_410),
.B2(n_387),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_310),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_372),
.B(n_391),
.C(n_405),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_329),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_373),
.B(n_377),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_321),
.B(n_310),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_374),
.B(n_368),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_327),
.B(n_278),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_378),
.B(n_406),
.Y(n_418)
);

INVxp33_ASAP7_75t_L g433 ( 
.A(n_383),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_322),
.A2(n_270),
.B1(n_308),
.B2(n_317),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_384),
.B(n_394),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_390),
.B(n_404),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_360),
.B(n_318),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_328),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_393),
.B(n_397),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_322),
.A2(n_308),
.B1(n_317),
.B2(n_314),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_339),
.A2(n_308),
.B(n_278),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_396),
.A2(n_402),
.B(n_355),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_336),
.A2(n_267),
.B1(n_263),
.B2(n_283),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_400),
.A2(n_401),
.B1(n_352),
.B2(n_344),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_335),
.A2(n_267),
.B1(n_263),
.B2(n_283),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_333),
.A2(n_289),
.B(n_319),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_324),
.B(n_359),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_339),
.B(n_319),
.C(n_307),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_326),
.B(n_307),
.C(n_294),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_342),
.A2(n_263),
.B1(n_267),
.B2(n_293),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_407),
.B(n_353),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_323),
.B(n_294),
.C(n_293),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_408),
.B(n_358),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_410),
.A2(n_396),
.B(n_402),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_411),
.A2(n_422),
.B1(n_434),
.B2(n_388),
.Y(n_450)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_385),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_412),
.B(n_413),
.Y(n_462)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_385),
.Y(n_413)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_371),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_415),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_416),
.A2(n_429),
.B1(n_432),
.B2(n_439),
.Y(n_466)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_382),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_419),
.B(n_424),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_421),
.B(n_443),
.C(n_378),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_394),
.A2(n_367),
.B1(n_365),
.B2(n_350),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_425),
.A2(n_431),
.B(n_436),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_395),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_426),
.B(n_427),
.Y(n_470)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_382),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_381),
.B(n_338),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_428),
.B(n_437),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_389),
.B(n_343),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_430),
.Y(n_448)
);

NAND2x1_ASAP7_75t_L g431 ( 
.A(n_375),
.B(n_343),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_370),
.A2(n_340),
.B1(n_348),
.B2(n_349),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_384),
.A2(n_320),
.B1(n_325),
.B2(n_345),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_406),
.B(n_306),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_438),
.B(n_372),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_401),
.A2(n_362),
.B1(n_346),
.B2(n_345),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_389),
.B(n_366),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_440),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_409),
.B(n_364),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_441),
.Y(n_469)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_399),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_442),
.B(n_446),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_374),
.B(n_330),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_400),
.A2(n_375),
.B1(n_409),
.B2(n_398),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_444),
.A2(n_445),
.B1(n_447),
.B2(n_386),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_375),
.A2(n_346),
.B1(n_357),
.B2(n_332),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_403),
.B(n_361),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_398),
.A2(n_403),
.B1(n_376),
.B2(n_391),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_450),
.A2(n_416),
.B1(n_439),
.B2(n_411),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_418),
.B(n_376),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_451),
.B(n_452),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_417),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_454),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_435),
.B(n_408),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_455),
.B(n_456),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_418),
.B(n_405),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_443),
.B(n_369),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_457),
.B(n_459),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_421),
.B(n_395),
.C(n_379),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_472),
.C(n_476),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_447),
.B(n_379),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_420),
.B(n_392),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_461),
.B(n_465),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_420),
.B(n_392),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_417),
.B(n_306),
.Y(n_467)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_467),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_438),
.B(n_388),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_471),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_431),
.B(n_430),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_431),
.B(n_386),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_474),
.A2(n_413),
.B1(n_415),
.B2(n_442),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_446),
.B(n_380),
.C(n_273),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_441),
.B(n_380),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_477),
.B(n_479),
.C(n_480),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_423),
.B(n_288),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_478),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_426),
.B(n_288),
.C(n_284),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_440),
.B(n_444),
.C(n_436),
.Y(n_480)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_470),
.Y(n_483)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_483),
.Y(n_510)
);

BUFx24_ASAP7_75t_SL g485 ( 
.A(n_475),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_485),
.B(n_465),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_469),
.B(n_428),
.Y(n_488)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_488),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_466),
.A2(n_474),
.B1(n_463),
.B2(n_414),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_491),
.B(n_500),
.Y(n_520)
);

XNOR2x2_ASAP7_75t_SL g492 ( 
.A(n_472),
.B(n_459),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_492),
.B(n_501),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_451),
.B(n_445),
.C(n_434),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_493),
.B(n_498),
.C(n_505),
.Y(n_517)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_470),
.Y(n_495)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_495),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_479),
.Y(n_496)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_496),
.Y(n_513)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_462),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_497),
.B(n_499),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_461),
.B(n_432),
.C(n_414),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_473),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_466),
.A2(n_429),
.B1(n_425),
.B2(n_433),
.Y(n_500)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_473),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_502),
.B(n_504),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_448),
.A2(n_422),
.B1(n_424),
.B2(n_412),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_456),
.B(n_427),
.C(n_419),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_507),
.B(n_477),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_488),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_508),
.B(n_516),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_SL g509 ( 
.A(n_494),
.B(n_457),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_509),
.B(n_521),
.Y(n_540)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_514),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_484),
.B(n_458),
.C(n_452),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_518),
.B(n_519),
.C(n_522),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_484),
.B(n_476),
.C(n_468),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_490),
.B(n_480),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_503),
.B(n_460),
.C(n_455),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_490),
.B(n_460),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_523),
.B(n_489),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_503),
.B(n_464),
.C(n_471),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_525),
.B(n_527),
.C(n_505),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_SL g526 ( 
.A(n_494),
.B(n_450),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_526),
.B(n_528),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_487),
.B(n_449),
.C(n_407),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_SL g528 ( 
.A(n_489),
.B(n_449),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_500),
.A2(n_289),
.B(n_13),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_530),
.A2(n_481),
.B(n_504),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g531 ( 
.A(n_524),
.Y(n_531)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_531),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_511),
.A2(n_501),
.B1(n_506),
.B2(n_482),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_533),
.A2(n_538),
.B1(n_539),
.B2(n_543),
.Y(n_562)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_534),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_536),
.B(n_547),
.Y(n_551)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_510),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_537),
.B(n_542),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_512),
.A2(n_493),
.B1(n_498),
.B2(n_491),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_520),
.A2(n_529),
.B1(n_530),
.B2(n_527),
.Y(n_539)
);

BUFx24_ASAP7_75t_SL g541 ( 
.A(n_521),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_541),
.B(n_532),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_520),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_515),
.A2(n_496),
.B1(n_487),
.B2(n_486),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_544),
.B(n_522),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_519),
.B(n_486),
.C(n_492),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_545),
.B(n_546),
.Y(n_561)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_525),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_514),
.B(n_10),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_534),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_550),
.B(n_556),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_552),
.B(n_557),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_536),
.B(n_517),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_554),
.B(n_555),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_532),
.B(n_517),
.C(n_518),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_549),
.B(n_523),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_535),
.B(n_513),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_558),
.B(n_540),
.Y(n_573)
);

AOI211xp5_ASAP7_75t_L g559 ( 
.A1(n_549),
.A2(n_515),
.B(n_526),
.C(n_528),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_559),
.A2(n_565),
.B1(n_562),
.B2(n_556),
.Y(n_568)
);

AO21x1_ASAP7_75t_L g560 ( 
.A1(n_547),
.A2(n_509),
.B(n_13),
.Y(n_560)
);

AO21x1_ASAP7_75t_L g576 ( 
.A1(n_560),
.A2(n_3),
.B(n_4),
.Y(n_576)
);

NOR2x1_ASAP7_75t_L g563 ( 
.A(n_548),
.B(n_16),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_563),
.A2(n_547),
.B(n_548),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_555),
.B(n_544),
.C(n_545),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_566),
.B(n_574),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_567),
.A2(n_570),
.B1(n_577),
.B2(n_3),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_SL g578 ( 
.A(n_568),
.B(n_573),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_553),
.A2(n_540),
.B1(n_16),
.B2(n_31),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_554),
.B(n_1),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_SL g575 ( 
.A1(n_561),
.A2(n_31),
.B(n_34),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_SL g585 ( 
.A1(n_575),
.A2(n_34),
.B(n_4),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_576),
.B(n_560),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_564),
.A2(n_34),
.B1(n_4),
.B2(n_5),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_571),
.B(n_551),
.C(n_558),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_579),
.B(n_581),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_566),
.B(n_551),
.C(n_563),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_569),
.Y(n_582)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_582),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_583),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_584),
.B(n_585),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_578),
.B(n_568),
.Y(n_590)
);

MAJx2_ASAP7_75t_L g592 ( 
.A(n_590),
.B(n_573),
.C(n_567),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_587),
.A2(n_580),
.B(n_572),
.Y(n_591)
);

OAI321xp33_ASAP7_75t_L g595 ( 
.A1(n_591),
.A2(n_588),
.A3(n_586),
.B1(n_583),
.B2(n_570),
.C(n_576),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_592),
.A2(n_593),
.B(n_590),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_589),
.Y(n_593)
);

OAI21x1_ASAP7_75t_L g596 ( 
.A1(n_594),
.A2(n_595),
.B(n_577),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_SL g597 ( 
.A1(n_596),
.A2(n_4),
.B(n_5),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_597),
.B(n_5),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_598),
.B(n_5),
.Y(n_599)
);


endmodule