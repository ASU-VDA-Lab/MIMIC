module real_jpeg_18364_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_524),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_0),
.B(n_525),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_1),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_1),
.B(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_1),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_1),
.B(n_126),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_1),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_1),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_1),
.B(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_2),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_3),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g412 ( 
.A(n_3),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_3),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_4),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_4),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_4),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_4),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_4),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_4),
.B(n_73),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_4),
.B(n_93),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_4),
.B(n_220),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_5),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_5),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_5),
.B(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_5),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_5),
.B(n_460),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_5),
.B(n_467),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_5),
.B(n_471),
.Y(n_470)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_6),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_6),
.Y(n_222)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_6),
.Y(n_270)
);

BUFx5_ASAP7_75t_L g474 ( 
.A(n_6),
.Y(n_474)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_7),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_7),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_7),
.B(n_124),
.Y(n_123)
);

NAND2x1_ASAP7_75t_SL g159 ( 
.A(n_7),
.B(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_7),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_7),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_8),
.B(n_224),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_8),
.B(n_257),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_8),
.B(n_309),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_8),
.B(n_64),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_8),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_8),
.B(n_448),
.Y(n_447)
);

AND2x2_ASAP7_75t_SL g456 ( 
.A(n_8),
.B(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_9),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_9),
.Y(n_126)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_9),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_10),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_11),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_11),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_12),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_12),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_12),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_SL g298 ( 
.A(n_12),
.B(n_299),
.Y(n_298)
);

AND2x2_ASAP7_75t_SL g358 ( 
.A(n_12),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_12),
.B(n_410),
.Y(n_409)
);

AND2x2_ASAP7_75t_SL g414 ( 
.A(n_12),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_12),
.B(n_220),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_14),
.B(n_142),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_14),
.B(n_179),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_14),
.Y(n_259)
);

AND2x2_ASAP7_75t_SL g274 ( 
.A(n_14),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_14),
.B(n_287),
.Y(n_286)
);

AND2x2_ASAP7_75t_SL g418 ( 
.A(n_14),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_14),
.B(n_423),
.Y(n_422)
);

BUFx4f_ASAP7_75t_L g94 ( 
.A(n_15),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_15),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_15),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_63),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_16),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_16),
.B(n_93),
.Y(n_92)
);

AND2x4_ASAP7_75t_SL g137 ( 
.A(n_16),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_16),
.B(n_142),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_16),
.B(n_145),
.Y(n_144)
);

NAND2x2_ASAP7_75t_SL g154 ( 
.A(n_16),
.B(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g162 ( 
.A(n_17),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_17),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_509),
.Y(n_19)
);

AO21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_244),
.B(n_503),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND3xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_166),
.C(n_239),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_23),
.A2(n_505),
.B(n_508),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_146),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_24),
.B(n_146),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_79),
.C(n_110),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_25),
.B(n_79),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_55),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_26),
.B(n_56),
.C(n_71),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_45),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_27),
.B(n_49),
.C(n_53),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_36),
.C(n_40),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_29),
.B(n_40),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_30),
.B(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_33),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_35),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g357 ( 
.A(n_35),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_36),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_36),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_36),
.A2(n_131),
.B1(n_517),
.B2(n_518),
.Y(n_516)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_38),
.Y(n_179)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_38),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_40),
.B(n_187),
.C(n_188),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_40),
.A2(n_41),
.B1(n_188),
.B2(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_43),
.Y(n_120)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_43),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_49),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_49),
.A2(n_54),
.B1(n_144),
.B2(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_49),
.A2(n_54),
.B1(n_189),
.B2(n_190),
.Y(n_212)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_52),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_52),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_54),
.B(n_135),
.C(n_144),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_54),
.B(n_186),
.C(n_189),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_71),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_61),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_57),
.B(n_62),
.C(n_67),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_61)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_62),
.A2(n_70),
.B1(n_154),
.B2(n_157),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_62),
.B(n_102),
.C(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_62),
.A2(n_70),
.B1(n_202),
.B2(n_203),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_62),
.B(n_97),
.C(n_154),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_65),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_67),
.B1(n_72),
.B2(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_66),
.B(n_121),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_72),
.C(n_76),
.Y(n_71)
);

MAJx2_ASAP7_75t_L g281 ( 
.A(n_67),
.B(n_122),
.C(n_282),
.Y(n_281)
);

OR2x2_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_68),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_72),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_SL g83 ( 
.A(n_72),
.B(n_84),
.C(n_91),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_72),
.A2(n_82),
.B1(n_91),
.B2(n_92),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_72),
.B(n_272),
.C(n_274),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_72),
.A2(n_82),
.B1(n_272),
.B2(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_75),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_76),
.B(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.C(n_95),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_80),
.B(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_83),
.B(n_95),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_90),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_137),
.C(n_141),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_91),
.A2(n_92),
.B1(n_137),
.B2(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_92),
.B(n_219),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_94),
.Y(n_417)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_94),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.C(n_105),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_96),
.A2(n_97),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

INVxp33_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_105),
.B1(n_106),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_102),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_102),
.A2(n_115),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx6_ASAP7_75t_L g401 ( 
.A(n_104),
.Y(n_401)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_111),
.B(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_129),
.C(n_134),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_112),
.B(n_236),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.C(n_127),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_113),
.B(n_116),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_123),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_117),
.A2(n_118),
.B1(n_123),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_125),
.Y(n_275)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2x2_ASAP7_75t_SL g194 ( 
.A(n_127),
.B(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_129),
.A2(n_130),
.B1(n_134),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_134),
.Y(n_237)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2x1_ASAP7_75t_L g191 ( 
.A(n_136),
.B(n_192),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_175),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_137),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_137),
.A2(n_175),
.B1(n_183),
.B2(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_137),
.B(n_422),
.Y(n_421)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_141),
.A2(n_154),
.B(n_519),
.Y(n_518)
);

NAND2xp33_ASAP7_75t_SL g519 ( 
.A(n_141),
.B(n_154),
.Y(n_519)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_143),
.Y(n_206)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_143),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_144),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_147),
.B(n_149),
.C(n_150),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_158),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_151),
.B(n_163),
.C(n_164),
.Y(n_513)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_154),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g214 ( 
.A(n_154),
.B(n_215),
.C(n_225),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_154),
.A2(n_157),
.B1(n_225),
.B2(n_332),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_159),
.Y(n_164)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_229),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_167),
.B(n_229),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_194),
.C(n_196),
.Y(n_167)
);

XNOR2x1_ASAP7_75t_L g385 ( 
.A(n_168),
.B(n_194),
.Y(n_385)
);

XOR2x1_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_184),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_169),
.B(n_185),
.C(n_191),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.C(n_181),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_170),
.B(n_173),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_180),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_175),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_175),
.B(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_175),
.A2(n_200),
.B1(n_264),
.B2(n_265),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_180),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_180),
.A2(n_307),
.B1(n_488),
.B2(n_489),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_181),
.B(n_373),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_183),
.B(n_422),
.Y(n_429)
);

XNOR2x1_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_191),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_196),
.B(n_385),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_210),
.C(n_213),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_197),
.B(n_371),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.C(n_207),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_198),
.B(n_201),
.Y(n_326)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2x2_ASAP7_75t_L g325 ( 
.A(n_207),
.B(n_326),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_371)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_215),
.B(n_331),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.C(n_223),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_216),
.B(n_219),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx5_ASAP7_75t_L g419 ( 
.A(n_221),
.Y(n_419)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_223),
.B(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_225),
.Y(n_332)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_227),
.Y(n_457)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_238),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_234),
.C(n_238),
.Y(n_243)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_240),
.A2(n_506),
.B(n_507),
.Y(n_505)
);

NOR2x1_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_241),
.B(n_243),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_387),
.Y(n_244)
);

A2O1A1O1Ixp25_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_364),
.B(n_378),
.C(n_379),
.D(n_386),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_336),
.B(n_363),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_322),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_248),
.B(n_322),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_294),
.C(n_315),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_249),
.B(n_338),
.Y(n_337)
);

XOR2x2_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_276),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_250),
.B(n_277),
.C(n_280),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_262),
.C(n_271),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_251),
.B(n_345),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_258),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.Y(n_252)
);

MAJx3_ASAP7_75t_L g321 ( 
.A(n_253),
.B(n_256),
.C(n_258),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_255),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_259),
.B(n_433),
.Y(n_432)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_262),
.A2(n_263),
.B1(n_271),
.B2(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_269),
.Y(n_304)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_271),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_272),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_274),
.B(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_285),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_281),
.B(n_286),
.C(n_291),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_282),
.B(n_296),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_291),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_294),
.B(n_315),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_297),
.C(n_306),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_295),
.B(n_297),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_302),
.B(n_305),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_302),
.Y(n_305)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_305),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_306),
.B(n_342),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.C(n_310),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_308),
.A2(n_310),
.B1(n_311),
.B2(n_490),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_308),
.Y(n_490)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_318),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_319),
.C(n_321),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_323),
.B(n_325),
.C(n_377),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_327),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g377 ( 
.A(n_327),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_328),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_330),
.A2(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_329)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_330),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_333),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_333),
.B(n_334),
.C(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_339),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_337),
.B(n_339),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_343),
.C(n_347),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_340),
.A2(n_341),
.B1(n_499),
.B2(n_500),
.Y(n_498)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_343),
.A2(n_344),
.B1(n_347),
.B2(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_347),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_351),
.C(n_352),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_348),
.B(n_493),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_351),
.B(n_352),
.Y(n_493)
);

MAJx2_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_358),
.C(n_362),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_353),
.A2(n_354),
.B1(n_362),
.B2(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_357),
.Y(n_356)
);

XNOR2x2_ASAP7_75t_L g440 ( 
.A(n_358),
.B(n_441),
.Y(n_440)
);

INVx5_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_362),
.Y(n_442)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_363),
.Y(n_390)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_365),
.B(n_380),
.Y(n_389)
);

AND2x2_ASAP7_75t_SL g365 ( 
.A(n_366),
.B(n_376),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_366),
.B(n_376),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_369),
.Y(n_366)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_367),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_370),
.A2(n_372),
.B1(n_374),
.B2(n_375),
.Y(n_369)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_370),
.Y(n_375)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_372),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_372),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_375),
.B(n_382),
.C(n_383),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_384),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_381),
.B(n_384),
.Y(n_386)
);

NAND4xp25_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_389),
.C(n_390),
.D(n_391),
.Y(n_387)
);

OAI21x1_ASAP7_75t_SL g391 ( 
.A1(n_392),
.A2(n_496),
.B(n_502),
.Y(n_391)
);

AOI21x1_ASAP7_75t_SL g392 ( 
.A1(n_393),
.A2(n_484),
.B(n_495),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_394),
.A2(n_443),
.B(n_483),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_427),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_395),
.B(n_427),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_413),
.C(n_420),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_396),
.B(n_480),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_402),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_397),
.B(n_409),
.C(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_409),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_403),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_413),
.A2(n_420),
.B1(n_421),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_413),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_418),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_414),
.B(n_418),
.Y(n_453)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_437),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_428),
.B(n_438),
.C(n_440),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_429),
.B(n_432),
.C(n_435),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_431),
.A2(n_432),
.B1(n_435),
.B2(n_436),
.Y(n_430)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_431),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_432),
.Y(n_436)
);

INVx6_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_440),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_477),
.B(n_482),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_445),
.A2(n_464),
.B(n_476),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_452),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_446),
.B(n_452),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_451),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_447),
.B(n_451),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_447),
.B(n_470),
.Y(n_469)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_454),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_453),
.B(n_456),
.C(n_458),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_455),
.A2(n_456),
.B1(n_458),
.B2(n_459),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_456),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_457),
.Y(n_467)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_465),
.A2(n_469),
.B(n_475),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_468),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_466),
.B(n_468),
.Y(n_475)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx6_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

BUFx12f_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_478),
.B(n_479),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_485),
.B(n_494),
.Y(n_484)
);

NOR2xp67_ASAP7_75t_SL g495 ( 
.A(n_485),
.B(n_494),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_492),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_491),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_487),
.B(n_491),
.C(n_492),
.Y(n_497)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_497),
.B(n_498),
.Y(n_502)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_523),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_522),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_512),
.B(n_522),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_514),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_515),
.A2(n_516),
.B1(n_520),
.B2(n_521),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_515),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_516),
.Y(n_521)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_518),
.Y(n_517)
);


endmodule