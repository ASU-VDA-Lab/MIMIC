module fake_jpeg_23763_n_327 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_1),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_17),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_38),
.A2(n_31),
.B1(n_20),
.B2(n_32),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_8),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_43),
.B(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx6p67_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_8),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_50),
.B(n_57),
.Y(n_106)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_58),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_49),
.A2(n_17),
.B1(n_26),
.B2(n_21),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_22),
.B1(n_25),
.B2(n_29),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_35),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_39),
.B(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_59),
.B(n_62),
.Y(n_113)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_72),
.Y(n_92)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_34),
.B(n_37),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_69),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_31),
.B1(n_20),
.B2(n_32),
.Y(n_83)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_26),
.B1(n_21),
.B2(n_22),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_73),
.A2(n_30),
.B1(n_27),
.B2(n_18),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_74),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_35),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_34),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_78),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_35),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_22),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_80),
.B(n_84),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_83),
.A2(n_67),
.B1(n_76),
.B2(n_77),
.Y(n_121)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_50),
.A2(n_21),
.B1(n_26),
.B2(n_25),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_85),
.A2(n_86),
.B1(n_71),
.B2(n_61),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_25),
.B1(n_35),
.B2(n_29),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_55),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_88),
.B(n_94),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_103),
.B1(n_114),
.B2(n_74),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_91),
.B(n_98),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_95),
.B(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g97 ( 
.A(n_63),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_97),
.A2(n_104),
.B1(n_105),
.B2(n_110),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_22),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_29),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_99),
.A2(n_19),
.B(n_9),
.Y(n_150)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_36),
.B1(n_33),
.B2(n_30),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_60),
.A2(n_36),
.B1(n_33),
.B2(n_18),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_77),
.A2(n_18),
.B1(n_30),
.B2(n_27),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_64),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_109),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_63),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_54),
.B(n_75),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_115),
.A2(n_37),
.B1(n_19),
.B2(n_2),
.Y(n_147)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_SL g118 ( 
.A(n_75),
.B(n_37),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_118),
.A2(n_37),
.B1(n_19),
.B2(n_9),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_125),
.B1(n_131),
.B2(n_142),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_122),
.A2(n_135),
.B1(n_138),
.B2(n_151),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_72),
.B(n_65),
.C(n_57),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_124),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_71),
.B1(n_61),
.B2(n_30),
.Y(n_125)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_132),
.B(n_141),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

INVxp67_ASAP7_75t_SL g176 ( 
.A(n_133),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_108),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_139),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_27),
.B1(n_18),
.B2(n_19),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_99),
.A2(n_27),
.B1(n_37),
.B2(n_19),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_92),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_85),
.A2(n_86),
.B1(n_98),
.B2(n_81),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_95),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_80),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_81),
.A2(n_37),
.B1(n_19),
.B2(n_2),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_152),
.B1(n_84),
.B2(n_110),
.Y(n_167)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_146),
.B(n_153),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

NAND2xp33_ASAP7_75t_SL g183 ( 
.A(n_148),
.B(n_10),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_13),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_L g151 ( 
.A1(n_109),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_81),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_83),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_129),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_165),
.Y(n_190)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_166),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_122),
.A2(n_91),
.B1(n_96),
.B2(n_100),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_158),
.A2(n_168),
.B1(n_175),
.B2(n_177),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_91),
.C(n_88),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_164),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_82),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_170),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_163),
.B(n_127),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_117),
.C(n_107),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_167),
.B(n_169),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_153),
.A2(n_142),
.B1(n_135),
.B2(n_138),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_90),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_82),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_0),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_179),
.B(n_183),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_124),
.A2(n_90),
.B(n_94),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_130),
.B(n_119),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_150),
.C(n_125),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_174),
.B(n_185),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_140),
.A2(n_115),
.B1(n_116),
.B2(n_111),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_131),
.A2(n_97),
.B1(n_93),
.B2(n_87),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_178),
.A2(n_148),
.B1(n_141),
.B2(n_120),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_4),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_133),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_181),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_11),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_10),
.Y(n_182)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_4),
.C(n_5),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_152),
.Y(n_197)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_176),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_187),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_188),
.A2(n_208),
.B(n_217),
.Y(n_223)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_191),
.B(n_198),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_124),
.B1(n_144),
.B2(n_120),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_173),
.B1(n_168),
.B2(n_158),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_199),
.Y(n_219)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_154),
.B(n_121),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_130),
.Y(n_200)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_172),
.B(n_167),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_119),
.Y(n_202)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_203),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_204),
.Y(n_228)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_205),
.Y(n_231)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_210),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_157),
.B(n_136),
.Y(n_207)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_207),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_173),
.A2(n_133),
.B(n_136),
.C(n_127),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_157),
.B(n_136),
.Y(n_209)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_165),
.B(n_123),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_178),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_212),
.Y(n_240)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_218),
.B(n_243),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_220),
.A2(n_230),
.B1(n_242),
.B2(n_212),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_160),
.B(n_177),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g254 ( 
.A1(n_221),
.A2(n_228),
.B1(n_235),
.B2(n_218),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_213),
.A2(n_161),
.B1(n_160),
.B2(n_174),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_226),
.A2(n_235),
.B1(n_217),
.B2(n_215),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_159),
.C(n_186),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_238),
.C(n_239),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_191),
.A2(n_183),
.B(n_179),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_175),
.B1(n_171),
.B2(n_179),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_185),
.C(n_171),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_123),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_193),
.B(n_126),
.C(n_5),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_197),
.C(n_211),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_213),
.A2(n_126),
.B1(n_4),
.B2(n_7),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_210),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_234),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_244),
.B(n_250),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_248),
.B1(n_260),
.B2(n_240),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_190),
.Y(n_246)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_226),
.B(n_195),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_256),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_228),
.B(n_189),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_261),
.C(n_238),
.Y(n_275)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_253),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_234),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_254),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_194),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_258),
.Y(n_266)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_259),
.A2(n_222),
.B1(n_229),
.B2(n_207),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_220),
.A2(n_194),
.B1(n_198),
.B2(n_199),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_206),
.C(n_209),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_224),
.B(n_216),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_196),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_225),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_263),
.A2(n_231),
.B1(n_225),
.B2(n_187),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_257),
.Y(n_265)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_L g268 ( 
.A1(n_263),
.A2(n_221),
.B1(n_240),
.B2(n_243),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_268),
.A2(n_271),
.B1(n_278),
.B2(n_237),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_277),
.Y(n_288)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_259),
.A2(n_221),
.B1(n_219),
.B2(n_229),
.Y(n_271)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

A2O1A1Ixp33_ASAP7_75t_L g274 ( 
.A1(n_254),
.A2(n_219),
.B(n_223),
.C(n_196),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_274),
.A2(n_202),
.B(n_200),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_247),
.C(n_261),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_268),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_241),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_258),
.A2(n_237),
.B1(n_233),
.B2(n_242),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_255),
.A2(n_249),
.B1(n_254),
.B2(n_252),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_279),
.A2(n_248),
.B1(n_260),
.B2(n_254),
.Y(n_286)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_264),
.B(n_189),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_283),
.B(n_284),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_286),
.A2(n_270),
.B1(n_281),
.B2(n_230),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_273),
.C(n_251),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_266),
.A2(n_231),
.B(n_233),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_292),
.B(n_232),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_290),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_247),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_275),
.Y(n_298)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_267),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_257),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_298),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_291),
.A2(n_274),
.B1(n_271),
.B2(n_278),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_300),
.A2(n_304),
.B1(n_285),
.B2(n_286),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_301),
.A2(n_287),
.B(n_289),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_305),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_303),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_244),
.B1(n_203),
.B2(n_187),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_277),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_310),
.Y(n_315)
);

OR2x2_ASAP7_75t_SL g307 ( 
.A(n_296),
.B(n_292),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_298),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_290),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_312),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_203),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_297),
.A3(n_282),
.B1(n_288),
.B2(n_304),
.C1(n_305),
.C2(n_204),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_307),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_316),
.A2(n_318),
.B(n_313),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_309),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_320),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_313),
.B(n_301),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_293),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_317),
.Y(n_324)
);

AOI221xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_322),
.B1(n_310),
.B2(n_188),
.C(n_192),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_6),
.C(n_13),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_6),
.Y(n_327)
);


endmodule