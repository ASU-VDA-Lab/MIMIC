module fake_jpeg_2001_n_131 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_21),
.B(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_40),
.Y(n_48)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_33),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_34),
.A2(n_22),
.B1(n_16),
.B2(n_23),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_12),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_4),
.Y(n_39)
);

NAND3xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_10),
.C(n_6),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVxp33_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_6),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_46),
.Y(n_57)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_25),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_22),
.B1(n_16),
.B2(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_12),
.B(n_7),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_54),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_18),
.C(n_15),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_45),
.C(n_28),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_14),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_53),
.B(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_14),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_15),
.Y(n_55)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_49),
.B1(n_64),
.B2(n_60),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_67),
.B(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_36),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_29),
.B1(n_32),
.B2(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_83),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_50),
.C(n_47),
.Y(n_74)
);

OAI32xp33_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_82),
.A3(n_73),
.B1(n_85),
.B2(n_84),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_65),
.B1(n_48),
.B2(n_55),
.Y(n_75)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_61),
.B(n_59),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_86),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_58),
.A2(n_64),
.B(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_81),
.Y(n_96)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_91),
.B1(n_90),
.B2(n_87),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_97),
.Y(n_99)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_71),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_71),
.B(n_98),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_80),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_98),
.B(n_70),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_77),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_99),
.C(n_104),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_86),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_102),
.B(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_103),
.B(n_105),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_87),
.B(n_90),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_92),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_106),
.B(n_107),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_110),
.C(n_114),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_88),
.C(n_89),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_101),
.Y(n_111)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_112),
.A2(n_114),
.B(n_108),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_118),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_113),
.A2(n_89),
.B1(n_93),
.B2(n_92),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_109),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_119),
.B(n_115),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_115),
.C(n_119),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_116),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_116),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_117),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_117),
.C(n_118),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_126),
.A2(n_127),
.B(n_124),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_123),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_117),
.Y(n_131)
);


endmodule