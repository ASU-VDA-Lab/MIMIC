module fake_jpeg_28437_n_167 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_47),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_17),
.B(n_48),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_15),
.B(n_11),
.Y(n_63)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_7),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_9),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

BUFx8_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_78),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_0),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_82),
.Y(n_87)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_1),
.B(n_2),
.Y(n_82)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_62),
.B1(n_60),
.B2(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_64),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_81),
.B1(n_56),
.B2(n_58),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_73),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_60),
.B1(n_57),
.B2(n_62),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

OA22x2_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_60),
.B1(n_73),
.B2(n_64),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_68),
.B(n_77),
.C(n_73),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_61),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_96),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_68),
.B1(n_72),
.B2(n_71),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_8),
.B(n_9),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_63),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_100),
.Y(n_133)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_103),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_67),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_107),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_69),
.B(n_59),
.C(n_55),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_112),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_98),
.B(n_51),
.Y(n_107)
);

NAND3xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_52),
.C(n_23),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_32),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_1),
.B(n_3),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_118),
.B(n_19),
.Y(n_136)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_3),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_113),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_24),
.C(n_46),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_115),
.C(n_119),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_20),
.C(n_42),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_117),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_4),
.B(n_5),
.C(n_7),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_30),
.C(n_40),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_100),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_137),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_97),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_127),
.B(n_136),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_49),
.B1(n_36),
.B2(n_37),
.Y(n_147)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_10),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_131),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_16),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_18),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_134),
.A2(n_38),
.B1(n_140),
.B2(n_124),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_105),
.B(n_25),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_27),
.Y(n_138)
);

XOR2x1_ASAP7_75t_SL g151 ( 
.A(n_138),
.B(n_35),
.Y(n_151)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_146),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_153),
.B1(n_133),
.B2(n_140),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_125),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_149),
.Y(n_154)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_150),
.B(n_152),
.Y(n_155)
);

NAND2x1p5_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_137),
.Y(n_156)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_156),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_139),
.C(n_145),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_161),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_143),
.C(n_138),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_159),
.B1(n_155),
.B2(n_154),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_132),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_151),
.A3(n_155),
.B1(n_143),
.B2(n_121),
.C1(n_141),
.C2(n_133),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_142),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_142),
.Y(n_167)
);


endmodule