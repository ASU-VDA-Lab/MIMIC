module fake_jpeg_28603_n_23 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_23);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_23;

wire n_13;
wire n_21;
wire n_10;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

AOI22xp33_ASAP7_75t_SL g7 ( 
.A1(n_4),
.A2(n_5),
.B1(n_1),
.B2(n_2),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_1),
.B(n_5),
.Y(n_8)
);

INVx13_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_3),
.B(n_1),
.Y(n_11)
);

AOI22xp33_ASAP7_75t_SL g12 ( 
.A1(n_2),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_0),
.B(n_3),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_8),
.B(n_2),
.C(n_11),
.Y(n_15)
);

AND2x6_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_16),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_14),
.B(n_8),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_14),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_17),
.A2(n_18),
.B1(n_10),
.B2(n_12),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_10),
.B(n_9),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_15),
.C(n_7),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_7),
.C(n_12),
.Y(n_22)
);

AOI322xp5_ASAP7_75t_L g23 ( 
.A1(n_22),
.A2(n_9),
.A3(n_13),
.B1(n_20),
.B2(n_21),
.C1(n_7),
.C2(n_19),
.Y(n_23)
);


endmodule