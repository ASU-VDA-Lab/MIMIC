module fake_jpeg_26654_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_7),
.B(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_SL g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_39),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_30),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_31),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_31),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_31),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_54),
.B(n_56),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_22),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_21),
.B1(n_28),
.B2(n_23),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_21),
.B1(n_34),
.B2(n_24),
.Y(n_67)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_21),
.B1(n_28),
.B2(n_18),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_63),
.A2(n_67),
.B1(n_29),
.B2(n_57),
.Y(n_98)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_22),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_68),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_70),
.B(n_72),
.Y(n_120)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_71),
.Y(n_102)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_75),
.Y(n_119)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_23),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_79),
.Y(n_116)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_58),
.A2(n_20),
.B1(n_26),
.B2(n_24),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_20),
.B1(n_26),
.B2(n_34),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_91),
.B1(n_93),
.B2(n_36),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_30),
.Y(n_90)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_58),
.A2(n_29),
.B1(n_55),
.B2(n_19),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_107),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_99),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_77),
.B1(n_80),
.B2(n_70),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_53),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_43),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_69),
.B(n_64),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_32),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_111),
.B(n_122),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_92),
.C(n_76),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_121),
.C(n_88),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_74),
.B(n_42),
.C(n_35),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_25),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_136),
.Y(n_157)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_146),
.Y(n_161)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_112),
.A2(n_72),
.B1(n_71),
.B2(n_67),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_143),
.B1(n_144),
.B2(n_148),
.Y(n_156)
);

OAI32xp33_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_84),
.A3(n_89),
.B1(n_82),
.B2(n_18),
.Y(n_129)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_132),
.B1(n_102),
.B2(n_119),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_17),
.B(n_93),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_131),
.A2(n_145),
.B(n_151),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_104),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_133),
.Y(n_169)
);

NOR3xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_17),
.C(n_11),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_14),
.Y(n_155)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_75),
.C(n_66),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_138),
.C(n_149),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_25),
.C(n_16),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_84),
.B1(n_62),
.B2(n_78),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_19),
.B1(n_18),
.B2(n_25),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_99),
.A2(n_19),
.B1(n_25),
.B2(n_32),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_115),
.B1(n_111),
.B2(n_105),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_121),
.A2(n_19),
.B1(n_32),
.B2(n_16),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_32),
.B1(n_16),
.B2(n_27),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_17),
.B(n_2),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_150),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_97),
.A2(n_16),
.B1(n_27),
.B2(n_4),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_95),
.B(n_27),
.C(n_10),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_9),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_102),
.A2(n_0),
.B(n_3),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_152),
.B(n_170),
.Y(n_204)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_155),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_140),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_123),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_168),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_113),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_167),
.B(n_174),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_110),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_172),
.B(n_176),
.Y(n_208)
);

CKINVDCx12_ASAP7_75t_R g173 ( 
.A(n_146),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_125),
.B(n_113),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_131),
.A2(n_103),
.B(n_119),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_183),
.B(n_151),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_101),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_124),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_0),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_148),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_179),
.Y(n_214)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_182),
.Y(n_202)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_132),
.Y(n_182)
);

XNOR2x2_ASAP7_75t_L g183 ( 
.A(n_125),
.B(n_12),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_135),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_184),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_144),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_180),
.B1(n_171),
.B2(n_182),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_186),
.A2(n_195),
.B1(n_200),
.B2(n_212),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_166),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_189),
.B(n_3),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_191),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_156),
.A2(n_145),
.B1(n_141),
.B2(n_138),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_193),
.A2(n_207),
.B1(n_211),
.B2(n_204),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_143),
.C(n_110),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_201),
.C(n_162),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_94),
.B1(n_108),
.B2(n_103),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_94),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_203),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_171),
.A2(n_108),
.B1(n_101),
.B2(n_117),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_101),
.C(n_117),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_9),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_174),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_205),
.B(n_210),
.Y(n_229)
);

NAND4xp25_ASAP7_75t_SL g206 ( 
.A(n_153),
.B(n_154),
.C(n_175),
.D(n_169),
.Y(n_206)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_156),
.A2(n_161),
.B1(n_177),
.B2(n_183),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_161),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_212)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_168),
.Y(n_217)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_221),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_165),
.Y(n_220)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_162),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_154),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_226),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_163),
.C(n_8),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_237),
.C(n_194),
.Y(n_242)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_227),
.Y(n_245)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_163),
.Y(n_228)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_232),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_211),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_241),
.B1(n_212),
.B2(n_216),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_0),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_233),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_262)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_235),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_195),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_201),
.C(n_209),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_240),
.Y(n_248)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_255),
.C(n_256),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_230),
.A2(n_210),
.B1(n_213),
.B2(n_186),
.Y(n_244)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_238),
.A2(n_236),
.B1(n_239),
.B2(n_219),
.Y(n_247)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_249),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_213),
.B1(n_191),
.B2(n_192),
.Y(n_253)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_203),
.C(n_192),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_190),
.C(n_206),
.Y(n_256)
);

FAx1_ASAP7_75t_SL g257 ( 
.A(n_229),
.B(n_196),
.CI(n_198),
.CON(n_257),
.SN(n_257)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_236),
.A2(n_198),
.B(n_10),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_259),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_10),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_231),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_228),
.A2(n_4),
.B(n_5),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_223),
.C(n_224),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_270),
.C(n_259),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_226),
.C(n_221),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_277),
.Y(n_280)
);

XOR2x2_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_222),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_276),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_232),
.Y(n_273)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

OA21x2_ASAP7_75t_SL g277 ( 
.A1(n_257),
.A2(n_222),
.B(n_220),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_243),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_279),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_217),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_256),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_285),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_251),
.B1(n_250),
.B2(n_246),
.Y(n_282)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_282),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_247),
.Y(n_284)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_272),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_263),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_286),
.B(n_288),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_289),
.C(n_270),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_278),
.B(n_248),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_254),
.C(n_253),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_254),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_294),
.B(n_4),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_266),
.A2(n_248),
.B1(n_262),
.B2(n_244),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_293),
.A2(n_8),
.B1(n_11),
.B2(n_15),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_258),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_287),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_291),
.A2(n_267),
.B1(n_266),
.B2(n_264),
.Y(n_296)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_276),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_297),
.B(n_300),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_267),
.C(n_264),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_301),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_274),
.B(n_260),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_281),
.A2(n_15),
.B(n_5),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_303),
.A2(n_5),
.B(n_7),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_283),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_307),
.A2(n_310),
.B(n_309),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_305),
.B(n_283),
.Y(n_308)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_308),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_314),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_315),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_292),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_298),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_317),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_297),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_319),
.A2(n_299),
.B1(n_300),
.B2(n_302),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_295),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_321),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_322),
.A2(n_319),
.B(n_316),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

AOI21x1_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_323),
.B(n_320),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_324),
.B(n_318),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_301),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_296),
.B(n_7),
.Y(n_330)
);


endmodule