module fake_jpeg_23498_n_178 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_32),
.Y(n_48)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_31),
.A2(n_36),
.B1(n_16),
.B2(n_19),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_13),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_24),
.B1(n_21),
.B2(n_17),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_40),
.B1(n_43),
.B2(n_49),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_38),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_42),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_35),
.B1(n_27),
.B2(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_14),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_28),
.A2(n_24),
.B1(n_21),
.B2(n_17),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_21),
.B1(n_17),
.B2(n_22),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_27),
.A2(n_21),
.B1(n_17),
.B2(n_22),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_31),
.B1(n_36),
.B2(n_27),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_19),
.B1(n_16),
.B2(n_14),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_30),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_54),
.B(n_65),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_59),
.B1(n_37),
.B2(n_43),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_52),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_36),
.B1(n_33),
.B2(n_29),
.Y(n_59)
);

OR2x2_ASAP7_75t_SL g60 ( 
.A(n_38),
.B(n_32),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_66),
.B(n_49),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_63),
.A2(n_46),
.B1(n_44),
.B2(n_19),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_42),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_20),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_14),
.C(n_18),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_68),
.B(n_69),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_47),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_70),
.A2(n_65),
.B1(n_61),
.B2(n_60),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_40),
.B1(n_45),
.B2(n_51),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_73),
.B1(n_74),
.B2(n_78),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_47),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_76),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_64),
.A2(n_40),
.B1(n_45),
.B2(n_51),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_29),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_82),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_54),
.A2(n_46),
.B1(n_29),
.B2(n_44),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_44),
.B1(n_22),
.B2(n_18),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_61),
.B1(n_62),
.B2(n_60),
.Y(n_95)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_87),
.Y(n_103)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_94),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_68),
.B(n_62),
.Y(n_101)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_91),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_90),
.A2(n_95),
.B1(n_70),
.B2(n_56),
.Y(n_115)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_99),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_81),
.B(n_58),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_62),
.C(n_63),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_82),
.C(n_73),
.Y(n_106)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_91),
.A2(n_80),
.B1(n_63),
.B2(n_76),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_113),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_75),
.B(n_81),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_107),
.B(n_115),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_85),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_104),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_113),
.C(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_84),
.B(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_108),
.B(n_111),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_58),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_56),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_71),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_0),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_102),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_118),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_89),
.B1(n_70),
.B2(n_93),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_121),
.C(n_115),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_93),
.C(n_98),
.Y(n_121)
);

NOR2xp67_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_89),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_105),
.B(n_112),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_55),
.C(n_20),
.Y(n_125)
);

FAx1_ASAP7_75t_SL g133 ( 
.A(n_125),
.B(n_101),
.CI(n_105),
.CON(n_133),
.SN(n_133)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_110),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_131),
.C(n_134),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_109),
.C(n_103),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_133),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_112),
.C(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_132),
.B(n_126),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_55),
.C(n_26),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_140),
.C(n_120),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_20),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_127),
.B(n_10),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

NAND4xp25_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_150),
.C(n_11),
.D(n_12),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_135),
.A2(n_129),
.B1(n_117),
.B2(n_127),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_147),
.B1(n_149),
.B2(n_143),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_129),
.B1(n_118),
.B2(n_123),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_149),
.B(n_7),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_125),
.B(n_10),
.Y(n_150)
);

OAI322xp33_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_13),
.A3(n_20),
.B1(n_15),
.B2(n_8),
.C1(n_4),
.C2(n_5),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_8),
.Y(n_154)
);

XNOR2x1_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_133),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_155),
.B(n_159),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_144),
.A2(n_137),
.B1(n_139),
.B2(n_11),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_154),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_26),
.C(n_23),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_157),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_145),
.B(n_7),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_4),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_147),
.A3(n_148),
.B1(n_15),
.B2(n_13),
.C1(n_26),
.C2(n_7),
.Y(n_160)
);

OAI321xp33_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_15),
.A3(n_26),
.B1(n_4),
.B2(n_11),
.C(n_12),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_148),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_165),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_154),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_155),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_163),
.B1(n_160),
.B2(n_168),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_12),
.Y(n_170)
);

AOI21xp33_ASAP7_75t_L g173 ( 
.A1(n_170),
.A2(n_171),
.B(n_0),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_164),
.A2(n_0),
.B(n_1),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_172),
.A2(n_173),
.A3(n_2),
.B1(n_3),
.B2(n_15),
.C1(n_167),
.C2(n_124),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

NOR2xp67_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_2),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_176),
.Y(n_178)
);


endmodule