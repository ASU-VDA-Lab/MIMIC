module fake_jpeg_30133_n_90 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_90);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_90;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_27),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_28),
.B(n_17),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_41),
.Y(n_47)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_29),
.Y(n_50)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_1),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_35),
.B1(n_34),
.B2(n_36),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_13),
.B(n_22),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_51),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_30),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_2),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_14),
.C(n_23),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_61),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_54),
.B(n_2),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_64),
.B(n_11),
.Y(n_69)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_12),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_68),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_16),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp67_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_21),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_4),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_74),
.A2(n_75),
.B1(n_18),
.B2(n_20),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_78),
.A2(n_79),
.B(n_68),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_67),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_73),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_77),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_84),
.B(n_77),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_85),
.B(n_71),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_81),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_80),
.C(n_72),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_25),
.Y(n_90)
);


endmodule