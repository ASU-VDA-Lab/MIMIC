module fake_jpeg_26103_n_296 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_296);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_33),
.B(n_37),
.Y(n_50)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx2_ASAP7_75t_SL g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_15),
.B1(n_30),
.B2(n_19),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_19),
.B1(n_30),
.B2(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_31),
.B1(n_29),
.B2(n_23),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_53),
.B1(n_55),
.B2(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_31),
.B1(n_25),
.B2(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_21),
.B1(n_18),
.B2(n_25),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_39),
.B1(n_32),
.B2(n_26),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_58),
.A2(n_64),
.B1(n_16),
.B2(n_20),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_60),
.B(n_28),
.Y(n_87)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_63),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_51),
.A2(n_39),
.B1(n_32),
.B2(n_26),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_15),
.B1(n_39),
.B2(n_32),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_66),
.A2(n_72),
.B1(n_35),
.B2(n_22),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_75),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

AO22x2_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_38),
.B1(n_35),
.B2(n_36),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_26),
.B1(n_28),
.B2(n_27),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_80),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_77),
.Y(n_102)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_79),
.A2(n_22),
.B1(n_17),
.B2(n_16),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_50),
.A2(n_26),
.B1(n_28),
.B2(n_27),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_81),
.Y(n_89)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_82),
.B(n_36),
.Y(n_98)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_47),
.B(n_1),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_86),
.A2(n_67),
.B(n_65),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_87),
.B(n_98),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_72),
.A2(n_16),
.B1(n_20),
.B2(n_27),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_88),
.A2(n_104),
.B1(n_77),
.B2(n_69),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_36),
.C(n_38),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_73),
.C(n_56),
.Y(n_112)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_95),
.Y(n_128)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_38),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_103),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_38),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_70),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_27),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_20),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_92),
.B1(n_63),
.B2(n_79),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_96),
.Y(n_151)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_89),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_17),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_120),
.B(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_124),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_27),
.C(n_62),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_137),
.C(n_105),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_74),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_57),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_129),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_126),
.A2(n_106),
.B1(n_91),
.B2(n_101),
.Y(n_139)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_87),
.B(n_99),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_104),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_138),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_0),
.B(n_2),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_134),
.A2(n_2),
.B(n_3),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_90),
.B1(n_93),
.B2(n_101),
.Y(n_147)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_2),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_12),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_0),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_139),
.A2(n_151),
.B(n_3),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_99),
.B1(n_85),
.B2(n_95),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_140),
.A2(n_166),
.B1(n_118),
.B2(n_123),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_112),
.A2(n_90),
.B1(n_85),
.B2(n_105),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_147),
.B1(n_150),
.B2(n_157),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_144),
.B(n_137),
.Y(n_173)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_146),
.Y(n_178)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_90),
.B1(n_96),
.B2(n_89),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_133),
.A2(n_101),
.B1(n_84),
.B2(n_107),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_84),
.Y(n_158)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_133),
.A2(n_135),
.B1(n_116),
.B2(n_111),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_121),
.B1(n_113),
.B2(n_114),
.Y(n_176)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_134),
.B(n_118),
.Y(n_171)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_126),
.A2(n_8),
.B1(n_12),
.B2(n_11),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_119),
.B(n_14),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_167),
.Y(n_186)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_120),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_169),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_R g202 ( 
.A(n_171),
.B(n_195),
.C(n_164),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_189),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_183),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_138),
.B1(n_131),
.B2(n_129),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_179),
.A2(n_191),
.B1(n_197),
.B2(n_166),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_180),
.A2(n_182),
.B1(n_160),
.B2(n_157),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_14),
.C(n_11),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_188),
.C(n_198),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_162),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_141),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_3),
.Y(n_185)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_8),
.C(n_11),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_14),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_168),
.A2(n_10),
.B(n_9),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_139),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_197),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_153),
.B(n_4),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_143),
.Y(n_206)
);

XOR2x1_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_5),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_152),
.A2(n_5),
.B(n_6),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_6),
.C(n_7),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_199),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_175),
.A2(n_149),
.B1(n_152),
.B2(n_141),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_203),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_202),
.A2(n_219),
.B(n_205),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_142),
.B1(n_154),
.B2(n_156),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_178),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_204),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_212),
.Y(n_225)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_211),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_184),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_209),
.B(n_216),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_195),
.B1(n_183),
.B2(n_172),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_213),
.A2(n_214),
.B1(n_187),
.B2(n_140),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_161),
.B1(n_163),
.B2(n_155),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_142),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_194),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_186),
.Y(n_216)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_170),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_196),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_208),
.B(n_154),
.Y(n_220)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_217),
.Y(n_223)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_212),
.B1(n_182),
.B2(n_174),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_205),
.A2(n_187),
.B1(n_185),
.B2(n_192),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_227),
.A2(n_202),
.B1(n_218),
.B2(n_171),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_217),
.A2(n_185),
.B(n_177),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_228),
.A2(n_237),
.B(n_155),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_232),
.C(n_234),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_177),
.C(n_181),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_214),
.B(n_219),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_233),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_189),
.C(n_198),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_231),
.B(n_210),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_248),
.Y(n_255)
);

O2A1O1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_233),
.A2(n_148),
.B(n_170),
.C(n_207),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_200),
.C(n_210),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_252),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_200),
.C(n_188),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_225),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_259),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_239),
.B(n_229),
.Y(n_259)
);

OAI221xp5_ASAP7_75t_L g260 ( 
.A1(n_250),
.A2(n_222),
.B1(n_231),
.B2(n_220),
.C(n_235),
.Y(n_260)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_230),
.Y(n_274)
);

XNOR2x1_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_228),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_264),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_255),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_269),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_263),
.A2(n_245),
.B(n_238),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_264),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_241),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_254),
.B(n_226),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_271),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_257),
.B(n_241),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_262),
.A2(n_230),
.B1(n_235),
.B2(n_236),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_272),
.A2(n_223),
.B1(n_243),
.B2(n_261),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_224),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_276),
.B(n_280),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_259),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_279),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_258),
.C(n_251),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_282),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_273),
.A2(n_245),
.B1(n_242),
.B2(n_227),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_266),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_285),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_275),
.A2(n_267),
.B(n_249),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_287),
.A2(n_280),
.B(n_249),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_L g289 ( 
.A1(n_286),
.A2(n_267),
.B(n_283),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_289),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_290),
.B(n_288),
.Y(n_292)
);

OAI321xp33_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_284),
.A3(n_277),
.B1(n_276),
.B2(n_268),
.C(n_253),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_293),
.A2(n_242),
.B(n_234),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_146),
.B(n_7),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_7),
.Y(n_296)
);


endmodule