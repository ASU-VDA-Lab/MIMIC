module fake_jpeg_3302_n_389 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_389);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_389;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_54),
.Y(n_134)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_56),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_24),
.B(n_9),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_57),
.B(n_67),
.Y(n_113)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_24),
.B(n_10),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_10),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_69),
.B(n_71),
.Y(n_126)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_70),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_19),
.B(n_44),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_73),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_33),
.B(n_8),
.C(n_15),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_78),
.Y(n_120)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_76),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_77),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_19),
.B(n_8),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_81),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_26),
.B(n_37),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_82),
.B(n_96),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_84),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_86),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_33),
.B(n_2),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g165 ( 
.A(n_87),
.B(n_98),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_88),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_95),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_26),
.B(n_8),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_97),
.B(n_107),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_20),
.B(n_7),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_20),
.B(n_12),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_102),
.Y(n_128)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_103),
.Y(n_168)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_105),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_108),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_39),
.B(n_12),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_109),
.B(n_57),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_96),
.A2(n_46),
.B1(n_43),
.B2(n_42),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_112),
.A2(n_129),
.B1(n_162),
.B2(n_163),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_57),
.A2(n_53),
.B1(n_48),
.B2(n_41),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_122),
.A2(n_133),
.B1(n_140),
.B2(n_20),
.Y(n_228)
);

OA22x2_ASAP7_75t_L g125 ( 
.A1(n_87),
.A2(n_50),
.B1(n_18),
.B2(n_48),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_125),
.B(n_117),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_65),
.A2(n_46),
.B1(n_53),
.B2(n_41),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_54),
.A2(n_50),
.B1(n_18),
.B2(n_52),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_131),
.A2(n_144),
.B1(n_145),
.B2(n_151),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_67),
.A2(n_39),
.B1(n_52),
.B2(n_32),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g140 ( 
.A1(n_66),
.A2(n_21),
.B1(n_36),
.B2(n_32),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_51),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_153),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_68),
.A2(n_51),
.B1(n_36),
.B2(n_31),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_72),
.A2(n_85),
.B1(n_73),
.B2(n_83),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_109),
.A2(n_21),
.B1(n_31),
.B2(n_14),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_71),
.B(n_14),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_86),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_154),
.A2(n_145),
.B1(n_144),
.B2(n_131),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_95),
.B(n_16),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_159),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_105),
.B(n_107),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_89),
.B(n_90),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_110),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_88),
.A2(n_3),
.B1(n_6),
.B2(n_102),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_84),
.A2(n_3),
.B1(n_35),
.B2(n_93),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_169),
.B(n_135),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_126),
.A2(n_172),
.B(n_128),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_175),
.A2(n_182),
.B(n_177),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_125),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_176),
.B(n_191),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_171),
.Y(n_178)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_178),
.Y(n_262)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_179),
.Y(n_232)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_181),
.A2(n_221),
.B1(n_200),
.B2(n_191),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_113),
.B(n_125),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_182),
.B(n_212),
.Y(n_230)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_183),
.Y(n_241)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_130),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_186),
.B(n_194),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_120),
.B(n_127),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

A2O1A1O1Ixp25_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_147),
.B(n_124),
.C(n_119),
.D(n_118),
.Y(n_190)
);

NOR3xp33_ASAP7_75t_L g231 ( 
.A(n_190),
.B(n_209),
.C(n_210),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_140),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_136),
.B(n_150),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_192),
.Y(n_247)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_171),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_L g249 ( 
.A1(n_195),
.A2(n_203),
.B(n_223),
.Y(n_249)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_197),
.B(n_202),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_115),
.A2(n_149),
.B1(n_134),
.B2(n_148),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_198),
.A2(n_224),
.B1(n_211),
.B2(n_183),
.Y(n_238)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_199),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_110),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_200),
.B(n_227),
.Y(n_258)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_201),
.B(n_215),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g203 ( 
.A1(n_162),
.A2(n_129),
.B(n_167),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_137),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_204),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_117),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_206),
.B(n_207),
.Y(n_263)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g208 ( 
.A(n_137),
.B(n_158),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_208),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_158),
.B(n_168),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_114),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_211),
.B(n_216),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_111),
.B(n_148),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_138),
.B(n_142),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_213),
.B(n_214),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_142),
.B(n_170),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_152),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_112),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_155),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_219),
.Y(n_245)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_114),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_218),
.Y(n_239)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_155),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_139),
.B(n_146),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_220),
.B(n_225),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_134),
.A2(n_164),
.B1(n_170),
.B2(n_156),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_139),
.B(n_146),
.C(n_156),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_208),
.C(n_178),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_164),
.B(n_87),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_141),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_120),
.B(n_153),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_226),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_141),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_228),
.A2(n_225),
.B1(n_195),
.B2(n_185),
.Y(n_260)
);

OR2x4_ASAP7_75t_L g233 ( 
.A(n_176),
.B(n_210),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_233),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_234),
.B(n_186),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_236),
.A2(n_217),
.B1(n_215),
.B2(n_189),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_238),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_190),
.A2(n_210),
.B(n_205),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_243),
.A2(n_250),
.B(n_252),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_202),
.A2(n_175),
.B(n_227),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_216),
.A2(n_209),
.B(n_212),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_228),
.A2(n_223),
.B1(n_224),
.B2(n_220),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_260),
.B1(n_222),
.B2(n_201),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_259),
.C(n_208),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_223),
.B(n_179),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_266),
.B(n_287),
.Y(n_308)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_232),
.Y(n_267)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_267),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_278),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_233),
.A2(n_218),
.B1(n_180),
.B2(n_219),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_269),
.A2(n_273),
.B1(n_274),
.B2(n_285),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_194),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_271),
.B(n_272),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_238),
.A2(n_240),
.B1(n_258),
.B2(n_260),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_178),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_275),
.B(n_277),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_193),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_184),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_240),
.B(n_204),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_279),
.B(n_282),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_229),
.B(n_196),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_281),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_246),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_234),
.B(n_199),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_283),
.Y(n_302)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_262),
.Y(n_284)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_284),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_258),
.A2(n_207),
.B1(n_253),
.B2(n_243),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_250),
.C(n_255),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_241),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_288),
.B(n_291),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_249),
.A2(n_231),
.B1(n_230),
.B2(n_265),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_289),
.A2(n_290),
.B1(n_293),
.B2(n_276),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_231),
.A2(n_230),
.B1(n_265),
.B2(n_251),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_251),
.B(n_242),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_261),
.A2(n_252),
.B1(n_241),
.B2(n_248),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_292),
.A2(n_261),
.B1(n_248),
.B2(n_242),
.Y(n_301)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_245),
.Y(n_294)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_294),
.Y(n_313)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_245),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_254),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_296),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_301),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_276),
.A2(n_263),
.B(n_245),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_306),
.A2(n_315),
.B(n_301),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_270),
.A2(n_246),
.B1(n_263),
.B2(n_239),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_295),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_271),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_297),
.Y(n_323)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_282),
.A2(n_239),
.A3(n_254),
.B1(n_264),
.B2(n_256),
.C1(n_237),
.C2(n_244),
.Y(n_315)
);

AOI221xp5_ASAP7_75t_L g335 ( 
.A1(n_317),
.A2(n_268),
.B1(n_296),
.B2(n_269),
.C(n_273),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_287),
.B(n_254),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_266),
.C(n_290),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_323),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_322),
.C(n_331),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_317),
.A2(n_292),
.B1(n_285),
.B2(n_291),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_321),
.A2(n_329),
.B1(n_333),
.B2(n_335),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_288),
.C(n_289),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_303),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_328),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_325),
.A2(n_336),
.B(n_298),
.Y(n_345)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_299),
.Y(n_326)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_326),
.Y(n_341)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_299),
.Y(n_327)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_327),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_314),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_278),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_306),
.A2(n_310),
.B(n_316),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_330),
.A2(n_332),
.B(n_313),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_308),
.B(n_279),
.C(n_272),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_316),
.A2(n_274),
.B(n_294),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_312),
.B(n_277),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_302),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_334),
.A2(n_300),
.B1(n_270),
.B2(n_305),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_338),
.A2(n_340),
.B1(n_345),
.B2(n_335),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_320),
.B(n_318),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_339),
.B(n_330),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_334),
.A2(n_300),
.B1(n_270),
.B2(n_305),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_322),
.C(n_325),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_346),
.B(n_348),
.C(n_350),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_322),
.B(n_314),
.C(n_309),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_349),
.B(n_329),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_332),
.B(n_309),
.C(n_313),
.Y(n_350)
);

OAI22x1_ASAP7_75t_L g351 ( 
.A1(n_347),
.A2(n_321),
.B1(n_323),
.B2(n_319),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_351),
.A2(n_340),
.B1(n_338),
.B2(n_342),
.Y(n_369)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_343),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_353),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_348),
.B(n_324),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_339),
.B(n_280),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_354),
.B(n_358),
.Y(n_368)
);

O2A1O1Ixp33_ASAP7_75t_L g363 ( 
.A1(n_355),
.A2(n_356),
.B(n_361),
.C(n_347),
.Y(n_363)
);

MAJx2_ASAP7_75t_L g366 ( 
.A(n_357),
.B(n_359),
.C(n_337),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_333),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_307),
.Y(n_359)
);

NOR3xp33_ASAP7_75t_SL g361 ( 
.A(n_344),
.B(n_336),
.C(n_327),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_351),
.A2(n_349),
.B(n_350),
.Y(n_362)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_362),
.Y(n_371)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_363),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_357),
.B(n_328),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_365),
.B(n_367),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_366),
.B(n_369),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_360),
.A2(n_359),
.B(n_346),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_365),
.B(n_360),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_372),
.B(n_375),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_364),
.B(n_368),
.Y(n_374)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_374),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_362),
.A2(n_361),
.B(n_341),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_376),
.B(n_326),
.C(n_304),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_378),
.B(n_379),
.C(n_286),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_372),
.B(n_304),
.C(n_311),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_373),
.B(n_302),
.Y(n_381)
);

NAND3xp33_ASAP7_75t_L g384 ( 
.A(n_381),
.B(n_371),
.C(n_275),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_377),
.B(n_375),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_382),
.A2(n_383),
.B(n_370),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_384),
.A2(n_381),
.B1(n_380),
.B2(n_286),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_385),
.B(n_386),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_387),
.A2(n_370),
.B(n_311),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_388),
.B(n_284),
.Y(n_389)
);


endmodule