module fake_ariane_3308_n_1754 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1754);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1754;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_2),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_159),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_103),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_49),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_46),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_99),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_62),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_116),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_45),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_81),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_64),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_101),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_142),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_23),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_53),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_33),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_40),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_3),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_2),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_160),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_33),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_127),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_80),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_26),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_86),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_8),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_57),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_49),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_22),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_131),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_37),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_5),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_9),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_108),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_41),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_74),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_51),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_115),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_68),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_143),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_73),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_132),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_27),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_93),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_14),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_5),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_162),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_117),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_84),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_56),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_24),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_133),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_3),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_138),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_85),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_112),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_13),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_125),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_60),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_48),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_48),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_146),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_82),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_157),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_70),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_12),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_92),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_149),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_129),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_91),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_7),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_124),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_114),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_19),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_88),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_139),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_55),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_76),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_145),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_130),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_98),
.Y(n_248)
);

BUFx8_ASAP7_75t_SL g249 ( 
.A(n_109),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_153),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_147),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_151),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_63),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_110),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_119),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_35),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_18),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_118),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_6),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_102),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_12),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_7),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_128),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_90),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_135),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_43),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_39),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_38),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_32),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_156),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_78),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_22),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_69),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_72),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_1),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_123),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_75),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_54),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_79),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_77),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_65),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_141),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_105),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_11),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_155),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_45),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_8),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_120),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_104),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_38),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_25),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_83),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_154),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_126),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_31),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_148),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_94),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_87),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_0),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_27),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_67),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_35),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_43),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_23),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_9),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_46),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_16),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_44),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_6),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_42),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_31),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_40),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_59),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_16),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_111),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_89),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_41),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_13),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_51),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_249),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_238),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_295),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_213),
.Y(n_323)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_295),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_165),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_174),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_290),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_295),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_187),
.B(n_0),
.Y(n_330)
);

INVxp33_ASAP7_75t_SL g331 ( 
.A(n_319),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_234),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_228),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_228),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_244),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_228),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_258),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_270),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_294),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_185),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_224),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_228),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_227),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_228),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_169),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_204),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_169),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_189),
.B(n_1),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_223),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_223),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_257),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_265),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_204),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_218),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_259),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_168),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_226),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_262),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_168),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_304),
.Y(n_360)
);

INVxp33_ASAP7_75t_SL g361 ( 
.A(n_163),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_306),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_307),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_226),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_273),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_266),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_273),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_232),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_277),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_267),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_292),
.B(n_4),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_170),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_272),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_277),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_286),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_163),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_212),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_178),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_191),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_166),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_166),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_309),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_L g383 ( 
.A(n_212),
.B(n_4),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_167),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_167),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_L g386 ( 
.A(n_284),
.B(n_10),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_199),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_L g388 ( 
.A(n_284),
.B(n_10),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_186),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_202),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_179),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_210),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_179),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_180),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_188),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_326),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_332),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_338),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_333),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_359),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_327),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_352),
.B(n_197),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_327),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_356),
.B(n_203),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_327),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_340),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_333),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_376),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_R g409 ( 
.A(n_320),
.B(n_201),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_339),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g411 ( 
.A(n_356),
.B(n_197),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_327),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_334),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_381),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_334),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_322),
.B(n_205),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_336),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_335),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_327),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_336),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_342),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_342),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_322),
.B(n_209),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_344),
.Y(n_424)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_372),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_337),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_341),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g428 ( 
.A1(n_345),
.A2(n_215),
.B(n_211),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_380),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_344),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_325),
.B(n_217),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_345),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_347),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_346),
.B(n_309),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_325),
.B(n_229),
.Y(n_435)
);

OA21x2_ASAP7_75t_L g436 ( 
.A1(n_347),
.A2(n_236),
.B(n_230),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_343),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_349),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_385),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_351),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_394),
.A2(n_269),
.B1(n_233),
.B2(n_173),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_355),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_372),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_349),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_384),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_354),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_360),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_350),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_350),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_368),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_357),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_357),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_358),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_382),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_366),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_364),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_370),
.B(n_164),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_359),
.B(n_263),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_329),
.B(n_243),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_364),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_365),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_373),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_365),
.Y(n_463)
);

OA21x2_ASAP7_75t_L g464 ( 
.A1(n_367),
.A2(n_251),
.B(n_247),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_367),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_369),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_369),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_434),
.B(n_443),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_432),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_399),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_400),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_432),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_402),
.B(n_382),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_438),
.Y(n_474)
);

AND2x6_ASAP7_75t_L g475 ( 
.A(n_458),
.B(n_174),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_457),
.B(n_331),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_400),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_400),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_451),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_427),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_399),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_437),
.B(n_375),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_404),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_439),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_420),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_420),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_353),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_420),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_454),
.B(n_440),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_421),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_442),
.Y(n_491)
);

AND2x6_ASAP7_75t_L g492 ( 
.A(n_458),
.B(n_174),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_407),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_407),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_434),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_458),
.B(n_329),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_425),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_413),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_451),
.Y(n_499)
);

BUFx10_ASAP7_75t_L g500 ( 
.A(n_453),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_451),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_443),
.B(n_389),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_413),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_454),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_436),
.A2(n_330),
.B1(n_348),
.B2(n_371),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_411),
.B(n_443),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_421),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_421),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_415),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_415),
.Y(n_510)
);

OAI21xp33_ASAP7_75t_L g511 ( 
.A1(n_416),
.A2(n_379),
.B(n_378),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_451),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_451),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_408),
.B(n_391),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_451),
.Y(n_515)
);

INVx6_ASAP7_75t_L g516 ( 
.A(n_425),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_L g517 ( 
.A(n_455),
.B(n_174),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_451),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_462),
.A2(n_383),
.B1(n_386),
.B2(n_388),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_411),
.B(n_389),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_408),
.B(n_323),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_417),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_443),
.B(n_395),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_401),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_429),
.B(n_324),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_460),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_417),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_409),
.B(n_393),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_436),
.A2(n_383),
.B1(n_395),
.B2(n_299),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_422),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_438),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_422),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_460),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_444),
.B(n_374),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_444),
.B(n_374),
.Y(n_535)
);

INVx1_ASAP7_75t_SL g536 ( 
.A(n_439),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_463),
.B(n_378),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_425),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_425),
.Y(n_539)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_404),
.Y(n_540)
);

AND2x6_ASAP7_75t_L g541 ( 
.A(n_463),
.B(n_174),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_445),
.B(n_321),
.Y(n_542)
);

NAND2xp33_ASAP7_75t_R g543 ( 
.A(n_396),
.B(n_328),
.Y(n_543)
);

BUFx10_ASAP7_75t_L g544 ( 
.A(n_397),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_425),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_424),
.Y(n_546)
);

NAND2xp33_ASAP7_75t_SL g547 ( 
.A(n_445),
.B(n_180),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_425),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_436),
.A2(n_220),
.B1(n_241),
.B2(n_318),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_460),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_L g551 ( 
.A(n_416),
.B(n_239),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_460),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_465),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_465),
.B(n_379),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_398),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_410),
.B(n_164),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_425),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_424),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_460),
.Y(n_559)
);

BUFx8_ASAP7_75t_SL g560 ( 
.A(n_414),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_430),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_423),
.B(n_387),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_430),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_460),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_460),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_423),
.B(n_171),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_450),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_431),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_433),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_433),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_433),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_448),
.B(n_387),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_448),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_448),
.B(n_390),
.Y(n_574)
);

NAND3xp33_ASAP7_75t_L g575 ( 
.A(n_431),
.B(n_377),
.C(n_182),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_449),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_449),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_435),
.B(n_390),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_435),
.B(n_392),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_436),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_449),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_436),
.A2(n_261),
.B1(n_302),
.B2(n_291),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_403),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_452),
.B(n_392),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_452),
.B(n_207),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_459),
.B(n_256),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_464),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_452),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_459),
.B(n_275),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_456),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_464),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_456),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_456),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_461),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_461),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_441),
.A2(n_308),
.B1(n_319),
.B2(n_317),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_464),
.A2(n_237),
.B1(n_214),
.B2(n_263),
.Y(n_597)
);

BUFx4f_ASAP7_75t_L g598 ( 
.A(n_464),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_441),
.B(n_450),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_464),
.A2(n_200),
.B1(n_317),
.B2(n_198),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_461),
.A2(n_200),
.B1(n_198),
.B2(n_196),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_466),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_403),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_466),
.Y(n_604)
);

OR2x6_ASAP7_75t_L g605 ( 
.A(n_414),
.B(n_253),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_466),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_467),
.B(n_280),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_467),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_467),
.B(n_171),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_428),
.B(n_172),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_401),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_428),
.A2(n_196),
.B1(n_181),
.B2(n_182),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_401),
.Y(n_613)
);

INVx1_ASAP7_75t_SL g614 ( 
.A(n_406),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_403),
.B(n_172),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_471),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_568),
.B(n_428),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_569),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_480),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_471),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_476),
.A2(n_194),
.B1(n_192),
.B2(n_190),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_483),
.B(n_540),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_600),
.A2(n_549),
.B1(n_582),
.B2(n_597),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_578),
.B(n_175),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_470),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_562),
.B(n_175),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_495),
.B(n_418),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_480),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_569),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_525),
.B(n_426),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_470),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_481),
.Y(n_632)
);

BUFx12f_ASAP7_75t_L g633 ( 
.A(n_500),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_484),
.B(n_446),
.Y(n_634)
);

AOI221xp5_ASAP7_75t_L g635 ( 
.A1(n_547),
.A2(n_181),
.B1(n_300),
.B2(n_287),
.C(n_183),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_612),
.A2(n_183),
.B1(n_193),
.B2(n_195),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_473),
.B(n_193),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_481),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_479),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_562),
.B(n_176),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_571),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_571),
.Y(n_642)
);

AOI22x1_ASAP7_75t_L g643 ( 
.A1(n_469),
.A2(n_472),
.B1(n_553),
.B2(n_474),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_514),
.B(n_176),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_579),
.B(n_177),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_493),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_581),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_579),
.B(n_177),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_493),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_468),
.B(n_495),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_598),
.B(n_184),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_593),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_468),
.B(n_184),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_598),
.B(n_190),
.Y(n_654)
);

BUFx12f_ASAP7_75t_L g655 ( 
.A(n_500),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_491),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_505),
.A2(n_310),
.B1(n_300),
.B2(n_303),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_586),
.B(n_192),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_586),
.B(n_194),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_590),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_589),
.B(n_531),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_589),
.B(n_289),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_494),
.Y(n_663)
);

NOR2x1p5_ASAP7_75t_L g664 ( 
.A(n_491),
.B(n_287),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_494),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_531),
.B(n_289),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_498),
.Y(n_667)
);

OR2x6_ASAP7_75t_L g668 ( 
.A(n_504),
.B(n_447),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_590),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_594),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_498),
.Y(n_671)
);

INVx8_ASAP7_75t_L g672 ( 
.A(n_475),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_537),
.B(n_296),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_536),
.Y(n_674)
);

A2O1A1Ixp33_ASAP7_75t_L g675 ( 
.A1(n_598),
.A2(n_281),
.B(n_288),
.C(n_293),
.Y(n_675)
);

A2O1A1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_511),
.A2(n_282),
.B(n_298),
.C(n_315),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_503),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_567),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_479),
.B(n_296),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_537),
.B(n_297),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_487),
.B(n_303),
.Y(n_681)
);

INVx8_ASAP7_75t_L g682 ( 
.A(n_475),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_566),
.B(n_305),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_556),
.B(n_305),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_502),
.B(n_297),
.Y(n_685)
);

INVx8_ASAP7_75t_L g686 ( 
.A(n_475),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_479),
.B(n_301),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_503),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_509),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_479),
.B(n_501),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_593),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_609),
.B(n_310),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_496),
.B(n_311),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_509),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_510),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_502),
.B(n_301),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_585),
.B(n_313),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_594),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_510),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_477),
.B(n_313),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_477),
.B(n_311),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_522),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_478),
.B(n_312),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_478),
.B(n_312),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_522),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_608),
.B(n_314),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_504),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_608),
.B(n_314),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_558),
.B(n_206),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_527),
.Y(n_710)
);

NOR3xp33_ASAP7_75t_L g711 ( 
.A(n_521),
.B(n_316),
.C(n_403),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_527),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_479),
.B(n_239),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_529),
.A2(n_363),
.B1(n_362),
.B2(n_285),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_501),
.B(n_239),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_561),
.B(n_208),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_530),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_575),
.B(n_11),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_530),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_532),
.Y(n_720)
);

OAI22xp33_ASAP7_75t_L g721 ( 
.A1(n_489),
.A2(n_596),
.B1(n_555),
.B2(n_519),
.Y(n_721)
);

O2A1O1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_554),
.A2(n_405),
.B(n_15),
.C(n_17),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_604),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_501),
.B(n_239),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_475),
.B(n_216),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_605),
.B(n_528),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_501),
.B(n_239),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_475),
.B(n_219),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_475),
.B(n_221),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_544),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_583),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_614),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_501),
.B(n_271),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_482),
.B(n_583),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_583),
.B(n_14),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_533),
.B(n_271),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_SL g737 ( 
.A(n_544),
.B(n_222),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_533),
.B(n_271),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_492),
.B(n_225),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_604),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_547),
.B(n_231),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_532),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_492),
.B(n_264),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_485),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_546),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_544),
.B(n_17),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_605),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_546),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_485),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_492),
.B(n_260),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_603),
.B(n_18),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_486),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_486),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_543),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_517),
.A2(n_235),
.B1(n_240),
.B2(n_248),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_492),
.B(n_276),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_605),
.B(n_405),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_563),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_517),
.A2(n_274),
.B1(n_245),
.B2(n_246),
.Y(n_759)
);

AO22x1_ASAP7_75t_L g760 ( 
.A1(n_542),
.A2(n_242),
.B1(n_250),
.B2(n_252),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_492),
.B(n_570),
.Y(n_761)
);

OR2x6_ASAP7_75t_L g762 ( 
.A(n_605),
.B(n_285),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_580),
.A2(n_271),
.B1(n_285),
.B2(n_405),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_533),
.B(n_271),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_SL g765 ( 
.A(n_599),
.B(n_283),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_563),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_492),
.A2(n_254),
.B1(n_255),
.B2(n_278),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_570),
.B(n_279),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_580),
.A2(n_591),
.B1(n_587),
.B2(n_573),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_573),
.B(n_405),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_488),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_576),
.B(n_419),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_572),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_576),
.B(n_419),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_577),
.B(n_419),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_587),
.A2(n_591),
.B1(n_577),
.B2(n_592),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_599),
.B(n_19),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_592),
.B(n_419),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_574),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_602),
.B(n_419),
.Y(n_780)
);

NOR2xp67_ASAP7_75t_L g781 ( 
.A(n_520),
.B(n_61),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_637),
.A2(n_607),
.B1(n_601),
.B2(n_615),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_622),
.A2(n_610),
.B(n_499),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_634),
.B(n_584),
.Y(n_784)
);

A2O1A1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_637),
.A2(n_606),
.B(n_602),
.C(n_588),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_661),
.B(n_606),
.Y(n_786)
);

O2A1O1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_657),
.A2(n_534),
.B(n_535),
.C(n_603),
.Y(n_787)
);

NOR3xp33_ASAP7_75t_L g788 ( 
.A(n_760),
.B(n_603),
.C(n_499),
.Y(n_788)
);

OR2x6_ASAP7_75t_L g789 ( 
.A(n_668),
.B(n_523),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_617),
.A2(n_499),
.B(n_526),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_650),
.B(n_595),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_624),
.B(n_488),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_625),
.Y(n_793)
);

OR2x6_ASAP7_75t_L g794 ( 
.A(n_668),
.B(n_506),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_690),
.A2(n_526),
.B(n_512),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_631),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_681),
.B(n_490),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_737),
.B(n_533),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_632),
.Y(n_799)
);

AOI21x1_ASAP7_75t_L g800 ( 
.A1(n_651),
.A2(n_512),
.B(n_515),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_638),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_618),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_681),
.B(n_490),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_646),
.A2(n_550),
.B1(n_513),
.B2(n_552),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_718),
.A2(n_552),
.B(n_518),
.C(n_550),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_651),
.A2(n_564),
.B(n_513),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_654),
.A2(n_564),
.B(n_613),
.Y(n_807)
);

O2A1O1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_626),
.A2(n_507),
.B(n_508),
.C(n_551),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_654),
.A2(n_613),
.B(n_533),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_721),
.B(n_565),
.Y(n_810)
);

OAI21xp5_ASAP7_75t_L g811 ( 
.A1(n_769),
.A2(n_507),
.B(n_508),
.Y(n_811)
);

OAI21xp33_ASAP7_75t_L g812 ( 
.A1(n_621),
.A2(n_551),
.B(n_559),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_639),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_640),
.B(n_565),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_645),
.B(n_565),
.Y(n_815)
);

OAI21xp33_ASAP7_75t_L g816 ( 
.A1(n_636),
.A2(n_559),
.B(n_565),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_770),
.A2(n_613),
.B(n_565),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_700),
.A2(n_559),
.B(n_611),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_623),
.A2(n_714),
.B1(n_777),
.B2(n_636),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_765),
.A2(n_559),
.B1(n_516),
.B2(n_541),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_630),
.A2(n_559),
.B1(n_516),
.B2(n_541),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_619),
.B(n_497),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_772),
.A2(n_611),
.B(n_524),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_774),
.A2(n_611),
.B(n_524),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_684),
.A2(n_516),
.B1(n_541),
.B2(n_557),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_775),
.A2(n_611),
.B(n_524),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_778),
.A2(n_611),
.B(n_524),
.Y(n_827)
);

AOI21x1_ASAP7_75t_L g828 ( 
.A1(n_761),
.A2(n_524),
.B(n_516),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_648),
.B(n_497),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_684),
.A2(n_541),
.B1(n_557),
.B2(n_548),
.Y(n_830)
);

NOR2xp67_ASAP7_75t_L g831 ( 
.A(n_674),
.B(n_560),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_627),
.B(n_560),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_780),
.A2(n_538),
.B(n_548),
.Y(n_833)
);

OR2x6_ASAP7_75t_L g834 ( 
.A(n_668),
.B(n_557),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_773),
.A2(n_548),
.B(n_545),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_779),
.A2(n_497),
.B(n_538),
.Y(n_836)
);

NOR3xp33_ASAP7_75t_L g837 ( 
.A(n_635),
.B(n_545),
.C(n_539),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_658),
.B(n_545),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_649),
.A2(n_538),
.B1(n_539),
.B2(n_285),
.Y(n_839)
);

O2A1O1Ixp33_ASAP7_75t_SL g840 ( 
.A1(n_644),
.A2(n_20),
.B(n_21),
.C(n_25),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_663),
.A2(n_539),
.B(n_419),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_659),
.B(n_541),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_619),
.B(n_401),
.Y(n_843)
);

INVxp67_ASAP7_75t_L g844 ( 
.A(n_678),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_639),
.Y(n_845)
);

INVx6_ASAP7_75t_L g846 ( 
.A(n_633),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_718),
.A2(n_285),
.B(n_401),
.C(n_412),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_732),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_639),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_665),
.A2(n_401),
.B1(n_412),
.B2(n_419),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_667),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_662),
.B(n_541),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_628),
.B(n_412),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_628),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_693),
.B(n_21),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_639),
.Y(n_856)
);

BUFx2_ASAP7_75t_L g857 ( 
.A(n_656),
.Y(n_857)
);

O2A1O1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_653),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_693),
.B(n_28),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_656),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_623),
.A2(n_412),
.B1(n_401),
.B2(n_32),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_726),
.B(n_29),
.Y(n_862)
);

BUFx8_ASAP7_75t_L g863 ( 
.A(n_655),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_747),
.B(n_412),
.Y(n_864)
);

NOR2xp67_ASAP7_75t_L g865 ( 
.A(n_754),
.B(n_95),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_673),
.B(n_30),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_680),
.B(n_30),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_671),
.A2(n_412),
.B(n_96),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_677),
.A2(n_412),
.B(n_71),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_688),
.A2(n_712),
.B(n_742),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_675),
.A2(n_66),
.B(n_152),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_689),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_694),
.A2(n_719),
.B(n_745),
.Y(n_873)
);

O2A1O1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_695),
.A2(n_36),
.B(n_39),
.C(n_42),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_699),
.A2(n_710),
.B(n_748),
.C(n_717),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_703),
.B(n_44),
.Y(n_876)
);

BUFx4f_ASAP7_75t_L g877 ( 
.A(n_762),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_730),
.B(n_47),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_702),
.A2(n_107),
.B(n_150),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_762),
.Y(n_880)
);

INVx3_ASAP7_75t_SL g881 ( 
.A(n_730),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_705),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_672),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_720),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_758),
.A2(n_766),
.B(n_731),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_731),
.A2(n_100),
.B(n_137),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_703),
.A2(n_47),
.B1(n_50),
.B2(n_52),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_726),
.B(n_52),
.Y(n_888)
);

O2A1O1Ixp33_ASAP7_75t_SL g889 ( 
.A1(n_679),
.A2(n_53),
.B(n_58),
.C(n_97),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_672),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_629),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_707),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_769),
.A2(n_113),
.B(n_121),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_734),
.B(n_122),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_757),
.Y(n_895)
);

NOR2xp67_ASAP7_75t_L g896 ( 
.A(n_701),
.B(n_134),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_768),
.A2(n_158),
.B(n_666),
.Y(n_897)
);

AO21x1_ASAP7_75t_L g898 ( 
.A1(n_679),
.A2(n_687),
.B(n_751),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_672),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_697),
.B(n_714),
.Y(n_900)
);

NOR2x1_ASAP7_75t_L g901 ( 
.A(n_762),
.B(n_664),
.Y(n_901)
);

O2A1O1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_685),
.A2(n_696),
.B(n_683),
.C(n_704),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_709),
.A2(n_716),
.B(n_734),
.Y(n_903)
);

AOI21xp33_ASAP7_75t_L g904 ( 
.A1(n_683),
.A2(n_692),
.B(n_706),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_687),
.A2(n_776),
.B(n_723),
.Y(n_905)
);

NAND3xp33_ASAP7_75t_L g906 ( 
.A(n_711),
.B(n_735),
.C(n_751),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_741),
.B(n_692),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_682),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_735),
.A2(n_708),
.B(n_691),
.C(n_652),
.Y(n_909)
);

OAI21xp33_ASAP7_75t_L g910 ( 
.A1(n_746),
.A2(n_643),
.B(n_755),
.Y(n_910)
);

AOI21xp33_ASAP7_75t_L g911 ( 
.A1(n_763),
.A2(n_691),
.B(n_652),
.Y(n_911)
);

OAI321xp33_ASAP7_75t_L g912 ( 
.A1(n_722),
.A2(n_676),
.A3(n_763),
.B1(n_776),
.B2(n_641),
.C(n_642),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_629),
.A2(n_723),
.B(n_749),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_641),
.A2(n_740),
.B(n_744),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_647),
.A2(n_752),
.B1(n_749),
.B2(n_771),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_647),
.A2(n_669),
.B(n_698),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_616),
.B(n_620),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_757),
.B(n_616),
.Y(n_918)
);

AOI21x1_ASAP7_75t_L g919 ( 
.A1(n_713),
.A2(n_733),
.B(n_764),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_682),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_682),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_660),
.Y(n_922)
);

OR2x2_ASAP7_75t_L g923 ( 
.A(n_669),
.B(n_670),
.Y(n_923)
);

AND2x4_ASAP7_75t_SL g924 ( 
.A(n_670),
.B(n_753),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_752),
.B(n_753),
.Y(n_925)
);

NOR3xp33_ASAP7_75t_L g926 ( 
.A(n_759),
.B(n_756),
.C(n_750),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_725),
.B(n_743),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_713),
.A2(n_733),
.B(n_715),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_715),
.A2(n_736),
.B(n_724),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_724),
.A2(n_738),
.B(n_727),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_686),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_686),
.B(n_767),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_781),
.A2(n_739),
.B(n_728),
.C(n_729),
.Y(n_933)
);

BUFx6f_ASAP7_75t_SL g934 ( 
.A(n_686),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_727),
.A2(n_764),
.B(n_736),
.C(n_738),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_765),
.B(n_326),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_622),
.A2(n_617),
.B(n_690),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_625),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_765),
.B(n_326),
.Y(n_939)
);

OAI21xp33_ASAP7_75t_L g940 ( 
.A1(n_637),
.A2(n_624),
.B(n_361),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_617),
.A2(n_598),
.B(n_610),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_637),
.A2(n_765),
.B1(n_476),
.B2(n_630),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_630),
.B(n_454),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_618),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_661),
.B(n_568),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_624),
.A2(n_625),
.B1(n_632),
.B2(n_631),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_661),
.B(n_568),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_622),
.A2(n_617),
.B(n_690),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_661),
.B(n_568),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_637),
.A2(n_718),
.B(n_661),
.C(n_476),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_625),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_661),
.B(n_568),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_625),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_637),
.A2(n_718),
.B(n_661),
.C(n_476),
.Y(n_954)
);

INVx4_ASAP7_75t_L g955 ( 
.A(n_672),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_765),
.B(n_326),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_737),
.B(n_480),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_622),
.A2(n_617),
.B(n_690),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_622),
.A2(n_617),
.B(n_690),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_661),
.B(n_568),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_661),
.B(n_568),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_622),
.A2(n_617),
.B(n_690),
.Y(n_962)
);

BUFx8_ASAP7_75t_SL g963 ( 
.A(n_633),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_661),
.B(n_568),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_903),
.A2(n_948),
.B(n_937),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_906),
.A2(n_959),
.B(n_958),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_793),
.Y(n_967)
);

AOI21x1_ASAP7_75t_L g968 ( 
.A1(n_800),
.A2(n_962),
.B(n_898),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_955),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_942),
.B(n_950),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_802),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_954),
.B(n_940),
.Y(n_972)
);

INVx6_ASAP7_75t_L g973 ( 
.A(n_863),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_946),
.A2(n_897),
.B(n_909),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_906),
.A2(n_941),
.B(n_885),
.Y(n_975)
);

AOI21xp33_ASAP7_75t_L g976 ( 
.A1(n_936),
.A2(n_956),
.B(n_939),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_783),
.A2(n_902),
.B(n_792),
.Y(n_977)
);

INVx6_ASAP7_75t_L g978 ( 
.A(n_863),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_945),
.A2(n_949),
.B(n_947),
.Y(n_979)
);

AOI22xp5_ASAP7_75t_L g980 ( 
.A1(n_943),
.A2(n_907),
.B1(n_832),
.B2(n_855),
.Y(n_980)
);

OAI21x1_ASAP7_75t_L g981 ( 
.A1(n_828),
.A2(n_916),
.B(n_914),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_895),
.B(n_860),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_819),
.B(n_860),
.Y(n_983)
);

AOI221x1_ASAP7_75t_L g984 ( 
.A1(n_816),
.A2(n_910),
.B1(n_871),
.B2(n_904),
.C(n_876),
.Y(n_984)
);

AOI21xp33_ASAP7_75t_L g985 ( 
.A1(n_900),
.A2(n_859),
.B(n_866),
.Y(n_985)
);

O2A1O1Ixp5_ASAP7_75t_L g986 ( 
.A1(n_785),
.A2(n_805),
.B(n_806),
.C(n_818),
.Y(n_986)
);

AOI21x1_ASAP7_75t_SL g987 ( 
.A1(n_867),
.A2(n_815),
.B(n_814),
.Y(n_987)
);

AO21x2_ASAP7_75t_L g988 ( 
.A1(n_905),
.A2(n_811),
.B(n_933),
.Y(n_988)
);

OAI21x1_ASAP7_75t_L g989 ( 
.A1(n_919),
.A2(n_807),
.B(n_913),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_881),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_952),
.A2(n_961),
.B(n_960),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_877),
.B(n_857),
.Y(n_992)
);

AO21x1_ASAP7_75t_L g993 ( 
.A1(n_894),
.A2(n_810),
.B(n_893),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_880),
.Y(n_994)
);

AOI21xp33_ASAP7_75t_L g995 ( 
.A1(n_784),
.A2(n_782),
.B(n_964),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_829),
.A2(n_838),
.B(n_803),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_796),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_799),
.B(n_801),
.Y(n_998)
);

O2A1O1Ixp5_ASAP7_75t_L g999 ( 
.A1(n_809),
.A2(n_798),
.B(n_804),
.C(n_847),
.Y(n_999)
);

OAI21x1_ASAP7_75t_L g1000 ( 
.A1(n_913),
.A2(n_811),
.B(n_929),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_846),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_870),
.A2(n_873),
.B(n_875),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_797),
.A2(n_817),
.B(n_841),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_851),
.B(n_882),
.Y(n_1004)
);

O2A1O1Ixp5_ASAP7_75t_L g1005 ( 
.A1(n_850),
.A2(n_843),
.B(n_853),
.C(n_852),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_884),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_787),
.A2(n_786),
.B(n_808),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_862),
.B(n_888),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_957),
.B(n_918),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_833),
.A2(n_791),
.B(n_917),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_836),
.A2(n_826),
.B(n_823),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_938),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_951),
.Y(n_1013)
);

INVx4_ASAP7_75t_L g1014 ( 
.A(n_890),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_824),
.A2(n_827),
.B(n_842),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_SL g1016 ( 
.A(n_963),
.B(n_877),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_953),
.B(n_844),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_912),
.A2(n_837),
.B(n_788),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_854),
.B(n_901),
.Y(n_1019)
);

INVx2_ASAP7_75t_SL g1020 ( 
.A(n_846),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_848),
.B(n_822),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_831),
.A2(n_789),
.B1(n_892),
.B2(n_834),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_890),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_835),
.A2(n_911),
.B(n_926),
.Y(n_1024)
);

CKINVDCx11_ASAP7_75t_R g1025 ( 
.A(n_834),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_789),
.B(n_834),
.Y(n_1026)
);

AO21x1_ASAP7_75t_L g1027 ( 
.A1(n_927),
.A2(n_928),
.B(n_930),
.Y(n_1027)
);

OAI22x1_ASAP7_75t_L g1028 ( 
.A1(n_887),
.A2(n_878),
.B1(n_864),
.B2(n_821),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_SL g1029 ( 
.A1(n_955),
.A2(n_934),
.B(n_932),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_922),
.B(n_861),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_812),
.A2(n_830),
.B(n_825),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_858),
.A2(n_874),
.B(n_896),
.C(n_865),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_890),
.B(n_921),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_891),
.B(n_944),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_794),
.B(n_923),
.Y(n_1035)
);

NAND2xp33_ASAP7_75t_L g1036 ( 
.A(n_813),
.B(n_849),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_839),
.A2(n_915),
.B(n_925),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_868),
.A2(n_869),
.B(n_935),
.Y(n_1038)
);

AOI21xp33_ASAP7_75t_L g1039 ( 
.A1(n_794),
.A2(n_924),
.B(n_820),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_794),
.B(n_872),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_886),
.A2(n_879),
.B(n_889),
.Y(n_1041)
);

AO31x2_ASAP7_75t_L g1042 ( 
.A1(n_840),
.A2(n_813),
.A3(n_845),
.B(n_849),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_813),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_920),
.Y(n_1044)
);

AOI21x1_ASAP7_75t_SL g1045 ( 
.A1(n_845),
.A2(n_849),
.B(n_856),
.Y(n_1045)
);

NAND2x1p5_ASAP7_75t_L g1046 ( 
.A(n_920),
.B(n_921),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_883),
.A2(n_899),
.B(n_908),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_883),
.A2(n_899),
.B(n_908),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_931),
.A2(n_790),
.B(n_800),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_921),
.B(n_942),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_950),
.A2(n_954),
.B(n_904),
.C(n_942),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_903),
.A2(n_948),
.B(n_937),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_906),
.A2(n_948),
.B(n_937),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_903),
.A2(n_948),
.B(n_937),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_790),
.A2(n_800),
.B(n_795),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_942),
.A2(n_950),
.B1(n_954),
.B2(n_906),
.Y(n_1056)
);

AND3x2_ASAP7_75t_L g1057 ( 
.A(n_936),
.B(n_956),
.C(n_939),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_942),
.B(n_495),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_943),
.B(n_630),
.Y(n_1059)
);

NAND2xp33_ASAP7_75t_L g1060 ( 
.A(n_855),
.B(n_859),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_793),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_943),
.Y(n_1062)
);

INVx4_ASAP7_75t_L g1063 ( 
.A(n_881),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_942),
.B(n_495),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_943),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_950),
.A2(n_954),
.B(n_904),
.C(n_942),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_790),
.A2(n_800),
.B(n_795),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_790),
.A2(n_800),
.B(n_795),
.Y(n_1068)
);

AOI21x1_ASAP7_75t_L g1069 ( 
.A1(n_800),
.A2(n_959),
.B(n_958),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_790),
.A2(n_800),
.B(n_795),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_903),
.A2(n_948),
.B(n_937),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_942),
.B(n_495),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_943),
.B(n_630),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_906),
.A2(n_948),
.B(n_937),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_793),
.Y(n_1075)
);

AO31x2_ASAP7_75t_L g1076 ( 
.A1(n_898),
.A2(n_805),
.A3(n_905),
.B(n_937),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_942),
.A2(n_630),
.B1(n_939),
.B2(n_936),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_903),
.A2(n_948),
.B(n_937),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_942),
.B(n_495),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_942),
.B(n_495),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_942),
.B(n_495),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_942),
.A2(n_950),
.B1(n_954),
.B2(n_906),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_942),
.B(n_495),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_903),
.A2(n_948),
.B(n_937),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_950),
.A2(n_954),
.B(n_904),
.C(n_942),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_890),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_802),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_906),
.A2(n_948),
.B(n_937),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_955),
.Y(n_1089)
);

AOI21x1_ASAP7_75t_L g1090 ( 
.A1(n_800),
.A2(n_959),
.B(n_958),
.Y(n_1090)
);

NAND2x1p5_ASAP7_75t_L g1091 ( 
.A(n_955),
.B(n_890),
.Y(n_1091)
);

INVxp67_ASAP7_75t_SL g1092 ( 
.A(n_877),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_942),
.B(n_495),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_890),
.Y(n_1094)
);

NAND2x1p5_ASAP7_75t_L g1095 ( 
.A(n_955),
.B(n_890),
.Y(n_1095)
);

INVx5_ASAP7_75t_L g1096 ( 
.A(n_890),
.Y(n_1096)
);

AOI21xp33_ASAP7_75t_L g1097 ( 
.A1(n_936),
.A2(n_956),
.B(n_939),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_802),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_SL g1099 ( 
.A1(n_894),
.A2(n_762),
.B(n_955),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_881),
.Y(n_1100)
);

AOI21x1_ASAP7_75t_L g1101 ( 
.A1(n_800),
.A2(n_959),
.B(n_958),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_790),
.A2(n_800),
.B(n_795),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_942),
.B(n_495),
.Y(n_1103)
);

AO31x2_ASAP7_75t_L g1104 ( 
.A1(n_898),
.A2(n_805),
.A3(n_905),
.B(n_937),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_903),
.A2(n_948),
.B(n_937),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_1062),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1077),
.A2(n_980),
.B1(n_970),
.B2(n_1056),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_967),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1059),
.A2(n_1073),
.B1(n_976),
.B2(n_1097),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_973),
.Y(n_1110)
);

OR2x6_ASAP7_75t_L g1111 ( 
.A(n_1099),
.B(n_982),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_990),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_971),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_1065),
.B(n_1008),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_1082),
.A2(n_1051),
.B1(n_1066),
.B2(n_1085),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_1100),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_1057),
.B(n_1009),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_1092),
.B(n_982),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_996),
.A2(n_1052),
.B(n_965),
.Y(n_1119)
);

AOI21xp33_ASAP7_75t_SL g1120 ( 
.A1(n_1001),
.A2(n_1020),
.B(n_1017),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_997),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_1050),
.B(n_995),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_994),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_1063),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1057),
.B(n_1017),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_SL g1126 ( 
.A(n_1063),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1058),
.B(n_1064),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1072),
.B(n_1079),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1080),
.B(n_1081),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1083),
.B(n_1093),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_973),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1006),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_973),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_1091),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1012),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_978),
.Y(n_1136)
);

OA21x2_ASAP7_75t_L g1137 ( 
.A1(n_1054),
.A2(n_1105),
.B(n_1084),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_1021),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1013),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_SL g1140 ( 
.A(n_1016),
.B(n_1092),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_994),
.Y(n_1141)
);

INVx3_ASAP7_75t_SL g1142 ( 
.A(n_978),
.Y(n_1142)
);

INVx3_ASAP7_75t_SL g1143 ( 
.A(n_978),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1087),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_998),
.B(n_1004),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_983),
.A2(n_1060),
.B1(n_1098),
.B2(n_972),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1103),
.A2(n_985),
.B(n_1018),
.C(n_1032),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1061),
.B(n_1075),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1034),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1025),
.B(n_1040),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_974),
.A2(n_1002),
.B(n_975),
.C(n_1074),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1035),
.Y(n_1152)
);

O2A1O1Ixp5_ASAP7_75t_L g1153 ( 
.A1(n_993),
.A2(n_974),
.B(n_1053),
.C(n_966),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1022),
.A2(n_991),
.B1(n_979),
.B2(n_1030),
.Y(n_1154)
);

AOI21xp33_ASAP7_75t_L g1155 ( 
.A1(n_1028),
.A2(n_1024),
.B(n_1009),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1019),
.Y(n_1156)
);

INVxp67_ASAP7_75t_L g1157 ( 
.A(n_992),
.Y(n_1157)
);

BUFx12f_ASAP7_75t_L g1158 ( 
.A(n_1023),
.Y(n_1158)
);

NAND2x1p5_ASAP7_75t_L g1159 ( 
.A(n_1096),
.B(n_1033),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1043),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_1026),
.B(n_1044),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_1086),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_1086),
.Y(n_1163)
);

INVx4_ASAP7_75t_SL g1164 ( 
.A(n_1033),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_1086),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1096),
.B(n_1014),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1042),
.Y(n_1167)
);

O2A1O1Ixp5_ASAP7_75t_SL g1168 ( 
.A1(n_1088),
.A2(n_1007),
.B(n_1041),
.C(n_1039),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1031),
.A2(n_977),
.B1(n_1037),
.B2(n_1089),
.Y(n_1169)
);

INVxp67_ASAP7_75t_L g1170 ( 
.A(n_1094),
.Y(n_1170)
);

BUFx4_ASAP7_75t_SL g1171 ( 
.A(n_1045),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1044),
.B(n_1014),
.Y(n_1172)
);

AND2x6_ASAP7_75t_L g1173 ( 
.A(n_969),
.B(n_1089),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_1036),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_977),
.A2(n_969),
.B1(n_1078),
.B2(n_1071),
.Y(n_1175)
);

INVx2_ASAP7_75t_SL g1176 ( 
.A(n_1094),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_1095),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1094),
.B(n_1046),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1042),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1029),
.B(n_1095),
.Y(n_1180)
);

INVxp67_ASAP7_75t_L g1181 ( 
.A(n_988),
.Y(n_1181)
);

OR2x2_ASAP7_75t_L g1182 ( 
.A(n_1076),
.B(n_1104),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_984),
.B(n_1027),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1010),
.B(n_988),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1010),
.A2(n_1038),
.B1(n_1048),
.B2(n_1003),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1047),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_SL g1187 ( 
.A(n_1038),
.B(n_1015),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1076),
.B(n_1104),
.Y(n_1188)
);

NAND3xp33_ASAP7_75t_L g1189 ( 
.A(n_986),
.B(n_1003),
.C(n_1005),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_1011),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_1045),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_968),
.B(n_1090),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1104),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_987),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1000),
.B(n_1104),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_986),
.A2(n_1005),
.B(n_1102),
.Y(n_1196)
);

HB1xp67_ASAP7_75t_L g1197 ( 
.A(n_989),
.Y(n_1197)
);

INVx4_ASAP7_75t_L g1198 ( 
.A(n_987),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1049),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1069),
.B(n_1101),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_999),
.A2(n_981),
.B(n_1055),
.C(n_1067),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1068),
.B(n_1070),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_996),
.A2(n_1052),
.B(n_965),
.Y(n_1203)
);

BUFx16f_ASAP7_75t_R g1204 ( 
.A(n_1057),
.Y(n_1204)
);

NAND2x1p5_ASAP7_75t_L g1205 ( 
.A(n_1096),
.B(n_877),
.Y(n_1205)
);

NAND2xp33_ASAP7_75t_L g1206 ( 
.A(n_1056),
.B(n_940),
.Y(n_1206)
);

O2A1O1Ixp5_ASAP7_75t_SL g1207 ( 
.A1(n_985),
.A2(n_1082),
.B(n_1056),
.C(n_966),
.Y(n_1207)
);

NAND2x1p5_ASAP7_75t_L g1208 ( 
.A(n_1096),
.B(n_877),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_996),
.A2(n_1052),
.B(n_965),
.Y(n_1209)
);

INVxp67_ASAP7_75t_L g1210 ( 
.A(n_1062),
.Y(n_1210)
);

OR2x6_ASAP7_75t_L g1211 ( 
.A(n_1099),
.B(n_762),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_967),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1077),
.A2(n_942),
.B1(n_954),
.B2(n_950),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_990),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1062),
.B(n_1065),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1059),
.B(n_1073),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_967),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1059),
.B(n_1073),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_967),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1077),
.B(n_439),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1077),
.A2(n_942),
.B(n_954),
.C(n_950),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_990),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1077),
.A2(n_942),
.B1(n_630),
.B2(n_939),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_967),
.Y(n_1224)
);

AOI222xp33_ASAP7_75t_L g1225 ( 
.A1(n_1059),
.A2(n_819),
.B1(n_636),
.B2(n_304),
.C1(n_185),
.C2(n_307),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1051),
.A2(n_1085),
.B(n_1066),
.Y(n_1226)
);

AO22x1_ASAP7_75t_L g1227 ( 
.A1(n_1092),
.A2(n_936),
.B1(n_956),
.B2(n_939),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_973),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_967),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1077),
.A2(n_942),
.B1(n_630),
.B2(n_939),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1062),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1059),
.B(n_936),
.Y(n_1232)
);

OR2x2_ASAP7_75t_SL g1233 ( 
.A(n_973),
.B(n_978),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_976),
.A2(n_936),
.B1(n_956),
.B2(n_939),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1092),
.B(n_895),
.Y(n_1235)
);

OR2x2_ASAP7_75t_L g1236 ( 
.A(n_1062),
.B(n_1065),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1077),
.A2(n_942),
.B1(n_954),
.B2(n_950),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1077),
.A2(n_942),
.B1(n_954),
.B2(n_950),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_996),
.A2(n_1052),
.B(n_965),
.Y(n_1239)
);

AO21x2_ASAP7_75t_L g1240 ( 
.A1(n_1183),
.A2(n_1201),
.B(n_1196),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_SL g1241 ( 
.A1(n_1226),
.A2(n_1115),
.B(n_1213),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_SL g1242 ( 
.A1(n_1226),
.A2(n_1115),
.B(n_1213),
.Y(n_1242)
);

OR2x6_ASAP7_75t_L g1243 ( 
.A(n_1111),
.B(n_1211),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1145),
.B(n_1220),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1225),
.A2(n_1107),
.B1(n_1206),
.B2(n_1234),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1148),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1108),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1121),
.Y(n_1248)
);

OAI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1223),
.A2(n_1230),
.B1(n_1232),
.B2(n_1107),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1132),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1207),
.A2(n_1221),
.B(n_1147),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1188),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1225),
.A2(n_1237),
.B1(n_1238),
.B2(n_1218),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1182),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1237),
.A2(n_1238),
.B1(n_1216),
.B2(n_1155),
.Y(n_1255)
);

AO21x2_ASAP7_75t_L g1256 ( 
.A1(n_1184),
.A2(n_1154),
.B(n_1167),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1135),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1112),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1139),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1212),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1193),
.B(n_1217),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1117),
.A2(n_1122),
.B1(n_1113),
.B2(n_1144),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1219),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1224),
.B(n_1229),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1116),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1195),
.B(n_1190),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1127),
.B(n_1128),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1129),
.B(n_1130),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1123),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1227),
.B(n_1106),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1110),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1198),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_1106),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1171),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1181),
.Y(n_1275)
);

BUFx4f_ASAP7_75t_SL g1276 ( 
.A(n_1142),
.Y(n_1276)
);

CKINVDCx11_ASAP7_75t_R g1277 ( 
.A(n_1143),
.Y(n_1277)
);

AO21x2_ASAP7_75t_L g1278 ( 
.A1(n_1154),
.A2(n_1179),
.B(n_1209),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1197),
.Y(n_1279)
);

AO21x2_ASAP7_75t_L g1280 ( 
.A1(n_1119),
.A2(n_1239),
.B(n_1203),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1111),
.A2(n_1125),
.B1(n_1152),
.B2(n_1109),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1111),
.A2(n_1156),
.B1(n_1211),
.B2(n_1149),
.Y(n_1282)
);

AOI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1140),
.A2(n_1150),
.B1(n_1118),
.B2(n_1157),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1202),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1141),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1160),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_1215),
.Y(n_1287)
);

INVx6_ASAP7_75t_L g1288 ( 
.A(n_1164),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_SL g1289 ( 
.A1(n_1140),
.A2(n_1204),
.B1(n_1211),
.B2(n_1118),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1137),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1231),
.A2(n_1146),
.B1(n_1138),
.B2(n_1236),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1137),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1114),
.B(n_1210),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1161),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1165),
.Y(n_1295)
);

CKINVDCx16_ASAP7_75t_R g1296 ( 
.A(n_1126),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1158),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1169),
.B(n_1153),
.Y(n_1298)
);

INVxp33_ASAP7_75t_L g1299 ( 
.A(n_1235),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1191),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1169),
.B(n_1194),
.Y(n_1301)
);

NAND2x1p5_ASAP7_75t_L g1302 ( 
.A(n_1174),
.B(n_1180),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1162),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_1186),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1228),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1168),
.B(n_1151),
.Y(n_1306)
);

OAI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1131),
.A2(n_1133),
.B1(n_1136),
.B2(n_1120),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1163),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1172),
.Y(n_1309)
);

AND2x4_ASAP7_75t_SL g1310 ( 
.A(n_1214),
.B(n_1222),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1189),
.A2(n_1124),
.B1(n_1233),
.B2(n_1222),
.Y(n_1311)
);

AO21x2_ASAP7_75t_L g1312 ( 
.A1(n_1189),
.A2(n_1192),
.B(n_1200),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1170),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1175),
.B(n_1134),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1202),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1173),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1176),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1178),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1164),
.B(n_1166),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1185),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1173),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1199),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1185),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1187),
.Y(n_1324)
);

BUFx8_ASAP7_75t_L g1325 ( 
.A(n_1214),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1214),
.A2(n_1222),
.B1(n_1208),
.B2(n_1205),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1187),
.A2(n_1177),
.B(n_1159),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1173),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1226),
.B(n_1107),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1148),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1225),
.A2(n_1220),
.B1(n_939),
.B2(n_956),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1223),
.A2(n_942),
.B1(n_1230),
.B2(n_1077),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1145),
.B(n_1220),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1148),
.Y(n_1334)
);

INVxp67_ASAP7_75t_L g1335 ( 
.A(n_1216),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1171),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1148),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1148),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1148),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1225),
.A2(n_1220),
.B1(n_939),
.B2(n_956),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1225),
.A2(n_1220),
.B1(n_939),
.B2(n_956),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_1233),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1225),
.A2(n_1220),
.B1(n_939),
.B2(n_956),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1148),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_SL g1345 ( 
.A1(n_1220),
.A2(n_936),
.B1(n_956),
.B2(n_939),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1223),
.A2(n_942),
.B1(n_1230),
.B2(n_1077),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1225),
.A2(n_1220),
.B1(n_939),
.B2(n_956),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1226),
.B(n_1107),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_SL g1349 ( 
.A1(n_1220),
.A2(n_936),
.B1(n_956),
.B2(n_939),
.Y(n_1349)
);

AO21x2_ASAP7_75t_L g1350 ( 
.A1(n_1251),
.A2(n_1306),
.B(n_1292),
.Y(n_1350)
);

AO21x2_ASAP7_75t_L g1351 ( 
.A1(n_1306),
.A2(n_1292),
.B(n_1290),
.Y(n_1351)
);

INVx3_ASAP7_75t_SL g1352 ( 
.A(n_1274),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1269),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1266),
.B(n_1254),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1267),
.B(n_1268),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1244),
.B(n_1333),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1332),
.A2(n_1346),
.B(n_1345),
.Y(n_1357)
);

INVx3_ASAP7_75t_L g1358 ( 
.A(n_1272),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1266),
.B(n_1254),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1325),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1329),
.B(n_1348),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1329),
.B(n_1348),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1325),
.Y(n_1363)
);

INVxp67_ASAP7_75t_L g1364 ( 
.A(n_1293),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1252),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1252),
.Y(n_1366)
);

INVxp67_ASAP7_75t_L g1367 ( 
.A(n_1285),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1261),
.B(n_1298),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1261),
.B(n_1298),
.Y(n_1369)
);

OAI21xp33_ASAP7_75t_SL g1370 ( 
.A1(n_1245),
.A2(n_1253),
.B(n_1255),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1296),
.B(n_1258),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1314),
.B(n_1284),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1314),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1295),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1284),
.B(n_1315),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1320),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1320),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1323),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1310),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1323),
.Y(n_1380)
);

INVx6_ASAP7_75t_L g1381 ( 
.A(n_1325),
.Y(n_1381)
);

AO21x1_ASAP7_75t_SL g1382 ( 
.A1(n_1324),
.A2(n_1300),
.B(n_1283),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1265),
.B(n_1335),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1272),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1247),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1264),
.B(n_1301),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1248),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1250),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1257),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1279),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1275),
.B(n_1279),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1312),
.B(n_1324),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1312),
.B(n_1259),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1260),
.Y(n_1394)
);

BUFx2_ASAP7_75t_SL g1395 ( 
.A(n_1274),
.Y(n_1395)
);

CKINVDCx6p67_ASAP7_75t_R g1396 ( 
.A(n_1277),
.Y(n_1396)
);

OR2x6_ASAP7_75t_L g1397 ( 
.A(n_1243),
.B(n_1288),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1309),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1327),
.B(n_1243),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1263),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1286),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1256),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1294),
.B(n_1256),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1278),
.B(n_1275),
.Y(n_1404)
);

INVx4_ASAP7_75t_L g1405 ( 
.A(n_1316),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1278),
.B(n_1240),
.Y(n_1406)
);

AO22x1_ASAP7_75t_L g1407 ( 
.A1(n_1328),
.A2(n_1336),
.B1(n_1299),
.B2(n_1270),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1287),
.B(n_1302),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1243),
.B(n_1327),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1304),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1278),
.B(n_1246),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1304),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1273),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1303),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1330),
.B(n_1334),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_1310),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1308),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1337),
.B(n_1338),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1339),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1316),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_1390),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1368),
.B(n_1280),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1351),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1351),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1368),
.B(n_1280),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1361),
.B(n_1280),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1369),
.B(n_1322),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1361),
.B(n_1328),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1357),
.A2(n_1249),
.B(n_1349),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1362),
.B(n_1321),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1403),
.B(n_1241),
.Y(n_1431)
);

CKINVDCx14_ASAP7_75t_R g1432 ( 
.A(n_1396),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1372),
.Y(n_1433)
);

NOR3xp33_ASAP7_75t_L g1434 ( 
.A(n_1370),
.B(n_1311),
.C(n_1336),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1373),
.B(n_1344),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1351),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1390),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1386),
.B(n_1406),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1350),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1396),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1350),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1372),
.B(n_1319),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1350),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1391),
.B(n_1354),
.Y(n_1444)
);

AO21x2_ASAP7_75t_L g1445 ( 
.A1(n_1402),
.A2(n_1241),
.B(n_1242),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1391),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1403),
.B(n_1242),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1372),
.B(n_1319),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1353),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1354),
.B(n_1291),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1393),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1376),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1411),
.B(n_1281),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_SL g1454 ( 
.A1(n_1392),
.A2(n_1347),
.B1(n_1343),
.B2(n_1341),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1392),
.B(n_1318),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1449),
.B(n_1398),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1449),
.B(n_1367),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1446),
.B(n_1374),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1446),
.B(n_1419),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1438),
.B(n_1375),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1438),
.B(n_1375),
.Y(n_1461)
);

AOI211xp5_ASAP7_75t_SL g1462 ( 
.A1(n_1434),
.A2(n_1371),
.B(n_1364),
.C(n_1420),
.Y(n_1462)
);

OAI221xp5_ASAP7_75t_L g1463 ( 
.A1(n_1429),
.A2(n_1340),
.B1(n_1331),
.B2(n_1355),
.C(n_1282),
.Y(n_1463)
);

OAI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1429),
.A2(n_1359),
.B1(n_1397),
.B2(n_1299),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1454),
.A2(n_1359),
.B1(n_1395),
.B2(n_1352),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1438),
.B(n_1404),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1435),
.B(n_1413),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1434),
.B(n_1352),
.Y(n_1468)
);

NOR2x1_ASAP7_75t_L g1469 ( 
.A(n_1445),
.B(n_1405),
.Y(n_1469)
);

AOI221xp5_ASAP7_75t_SL g1470 ( 
.A1(n_1431),
.A2(n_1383),
.B1(n_1395),
.B2(n_1404),
.C(n_1400),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1435),
.B(n_1414),
.Y(n_1471)
);

NAND3xp33_ASAP7_75t_L g1472 ( 
.A(n_1454),
.B(n_1417),
.C(n_1387),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_SL g1473 ( 
.A1(n_1432),
.A2(n_1289),
.B(n_1307),
.Y(n_1473)
);

NAND4xp25_ASAP7_75t_L g1474 ( 
.A(n_1421),
.B(n_1410),
.C(n_1356),
.D(n_1376),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1452),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1435),
.B(n_1418),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1433),
.B(n_1428),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1453),
.A2(n_1382),
.B1(n_1262),
.B2(n_1399),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1447),
.B(n_1352),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1435),
.B(n_1455),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1433),
.B(n_1377),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1433),
.B(n_1377),
.Y(n_1482)
);

NOR3xp33_ASAP7_75t_SL g1483 ( 
.A(n_1440),
.B(n_1305),
.C(n_1271),
.Y(n_1483)
);

OAI21xp5_ASAP7_75t_SL g1484 ( 
.A1(n_1432),
.A2(n_1326),
.B(n_1420),
.Y(n_1484)
);

NOR3xp33_ASAP7_75t_L g1485 ( 
.A(n_1431),
.B(n_1407),
.C(n_1358),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_SL g1486 ( 
.A(n_1447),
.B(n_1408),
.Y(n_1486)
);

NAND4xp25_ASAP7_75t_L g1487 ( 
.A(n_1421),
.B(n_1380),
.C(n_1378),
.D(n_1384),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1455),
.B(n_1418),
.Y(n_1488)
);

AND2x2_ASAP7_75t_SL g1489 ( 
.A(n_1442),
.B(n_1399),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1455),
.B(n_1385),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1428),
.B(n_1380),
.Y(n_1491)
);

OAI21xp33_ASAP7_75t_L g1492 ( 
.A1(n_1422),
.A2(n_1388),
.B(n_1401),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1455),
.B(n_1385),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1422),
.B(n_1412),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1444),
.B(n_1387),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1450),
.A2(n_1381),
.B1(n_1389),
.B2(n_1401),
.Y(n_1496)
);

NAND3xp33_ASAP7_75t_L g1497 ( 
.A(n_1439),
.B(n_1400),
.C(n_1388),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1453),
.A2(n_1382),
.B1(n_1409),
.B2(n_1397),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1422),
.B(n_1425),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1444),
.B(n_1389),
.Y(n_1500)
);

AOI221xp5_ASAP7_75t_L g1501 ( 
.A1(n_1439),
.A2(n_1394),
.B1(n_1415),
.B2(n_1366),
.C(n_1365),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1422),
.B(n_1412),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1425),
.B(n_1412),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1499),
.B(n_1426),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1499),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1466),
.B(n_1425),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1466),
.B(n_1460),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1480),
.B(n_1426),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1475),
.B(n_1425),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1475),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1489),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1495),
.B(n_1426),
.Y(n_1512)
);

NAND2x1p5_ASAP7_75t_L g1513 ( 
.A(n_1469),
.B(n_1489),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1489),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1461),
.B(n_1477),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1481),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1469),
.B(n_1442),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1481),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1497),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1500),
.B(n_1426),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1494),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_1456),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1492),
.B(n_1501),
.Y(n_1523)
);

NAND2x1_ASAP7_75t_L g1524 ( 
.A(n_1485),
.B(n_1421),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1502),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1503),
.B(n_1442),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1459),
.B(n_1444),
.Y(n_1527)
);

INVxp67_ASAP7_75t_SL g1528 ( 
.A(n_1497),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1482),
.B(n_1442),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1457),
.B(n_1440),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1458),
.B(n_1444),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1492),
.B(n_1491),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1490),
.Y(n_1533)
);

AND2x2_ASAP7_75t_SL g1534 ( 
.A(n_1498),
.B(n_1442),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1483),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1493),
.B(n_1452),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1523),
.B(n_1471),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1507),
.B(n_1470),
.Y(n_1538)
);

OR2x6_ASAP7_75t_L g1539 ( 
.A(n_1513),
.B(n_1407),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1523),
.B(n_1467),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1507),
.B(n_1470),
.Y(n_1541)
);

NAND4xp75_ASAP7_75t_L g1542 ( 
.A(n_1534),
.B(n_1468),
.C(n_1453),
.D(n_1486),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1531),
.B(n_1488),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1531),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1512),
.B(n_1520),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1522),
.B(n_1476),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1512),
.B(n_1474),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1535),
.B(n_1277),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1511),
.B(n_1442),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1507),
.B(n_1437),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1531),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1515),
.B(n_1437),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1522),
.B(n_1437),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1515),
.B(n_1430),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1527),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1527),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1527),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1530),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1519),
.B(n_1474),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1515),
.B(n_1506),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1512),
.B(n_1487),
.Y(n_1561)
);

OAI211xp5_ASAP7_75t_L g1562 ( 
.A1(n_1528),
.A2(n_1462),
.B(n_1472),
.C(n_1487),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1506),
.B(n_1427),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1508),
.B(n_1520),
.Y(n_1564)
);

INVxp67_ASAP7_75t_SL g1565 ( 
.A(n_1528),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1506),
.B(n_1427),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1526),
.B(n_1427),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1526),
.B(n_1427),
.Y(n_1568)
);

INVxp67_ASAP7_75t_L g1569 ( 
.A(n_1519),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1510),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1520),
.B(n_1451),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1533),
.B(n_1462),
.Y(n_1572)
);

AOI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1524),
.A2(n_1472),
.B(n_1465),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1508),
.B(n_1451),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1538),
.B(n_1524),
.Y(n_1575)
);

INVxp67_ASAP7_75t_SL g1576 ( 
.A(n_1565),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1563),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1538),
.B(n_1541),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1569),
.B(n_1533),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1570),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1541),
.B(n_1526),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1544),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1551),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1560),
.B(n_1526),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1558),
.B(n_1271),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1555),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1556),
.Y(n_1587)
);

AOI33xp33_ASAP7_75t_L g1588 ( 
.A1(n_1557),
.A2(n_1560),
.A3(n_1562),
.B1(n_1550),
.B2(n_1552),
.B3(n_1510),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1571),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1573),
.A2(n_1465),
.B(n_1484),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1572),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1571),
.Y(n_1592)
);

AND2x4_ASAP7_75t_SL g1593 ( 
.A(n_1549),
.B(n_1448),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1554),
.B(n_1526),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1540),
.B(n_1504),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1540),
.B(n_1504),
.Y(n_1596)
);

O2A1O1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1559),
.A2(n_1473),
.B(n_1463),
.C(n_1532),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1545),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1554),
.B(n_1529),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1546),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1567),
.B(n_1529),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1563),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1567),
.B(n_1529),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1566),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1549),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1545),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1568),
.B(n_1566),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1537),
.B(n_1504),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1548),
.B(n_1305),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1537),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1543),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1564),
.B(n_1509),
.Y(n_1612)
);

NAND2x1_ASAP7_75t_SL g1613 ( 
.A(n_1549),
.B(n_1517),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1574),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1542),
.A2(n_1534),
.B1(n_1496),
.B2(n_1464),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1547),
.B(n_1509),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1574),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1605),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1584),
.B(n_1576),
.Y(n_1619)
);

NOR2x1_ASAP7_75t_L g1620 ( 
.A(n_1590),
.B(n_1547),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1591),
.B(n_1561),
.Y(n_1621)
);

BUFx3_ASAP7_75t_L g1622 ( 
.A(n_1585),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1584),
.B(n_1511),
.Y(n_1623)
);

INVx1_ASAP7_75t_SL g1624 ( 
.A(n_1579),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_1615),
.B(n_1511),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1580),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1578),
.B(n_1568),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1610),
.B(n_1561),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1580),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1597),
.B(n_1550),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1609),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1595),
.B(n_1553),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1578),
.A2(n_1539),
.B1(n_1453),
.B2(n_1514),
.Y(n_1633)
);

NAND3xp33_ASAP7_75t_L g1634 ( 
.A(n_1588),
.B(n_1539),
.C(n_1473),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1595),
.B(n_1508),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_1598),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1605),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1605),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1575),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1598),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1575),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1582),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1600),
.A2(n_1539),
.B1(n_1514),
.B2(n_1534),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1596),
.B(n_1536),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1606),
.B(n_1276),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1606),
.B(n_1552),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1582),
.Y(n_1647)
);

INVxp67_ASAP7_75t_SL g1648 ( 
.A(n_1613),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1583),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1581),
.B(n_1601),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1581),
.B(n_1529),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1596),
.B(n_1536),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1583),
.Y(n_1653)
);

O2A1O1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1620),
.A2(n_1616),
.B(n_1608),
.C(n_1587),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1620),
.A2(n_1634),
.B1(n_1625),
.B2(n_1630),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1621),
.B(n_1608),
.Y(n_1656)
);

AOI21xp33_ASAP7_75t_L g1657 ( 
.A1(n_1634),
.A2(n_1587),
.B(n_1586),
.Y(n_1657)
);

NAND3xp33_ASAP7_75t_L g1658 ( 
.A(n_1642),
.B(n_1616),
.C(n_1592),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1622),
.Y(n_1659)
);

NAND4xp25_ASAP7_75t_L g1660 ( 
.A(n_1639),
.B(n_1617),
.C(n_1589),
.D(n_1614),
.Y(n_1660)
);

O2A1O1Ixp33_ASAP7_75t_L g1661 ( 
.A1(n_1624),
.A2(n_1539),
.B(n_1592),
.C(n_1614),
.Y(n_1661)
);

AOI211xp5_ASAP7_75t_L g1662 ( 
.A1(n_1624),
.A2(n_1484),
.B(n_1589),
.C(n_1617),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1643),
.A2(n_1611),
.B1(n_1514),
.B2(n_1496),
.Y(n_1663)
);

AO21x1_ASAP7_75t_L g1664 ( 
.A1(n_1648),
.A2(n_1593),
.B(n_1513),
.Y(n_1664)
);

NOR2x1_ASAP7_75t_L g1665 ( 
.A(n_1622),
.B(n_1360),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1650),
.Y(n_1666)
);

NOR3xp33_ASAP7_75t_L g1667 ( 
.A(n_1628),
.B(n_1612),
.C(n_1602),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1647),
.Y(n_1668)
);

OAI222xp33_ASAP7_75t_L g1669 ( 
.A1(n_1633),
.A2(n_1513),
.B1(n_1478),
.B2(n_1602),
.C1(n_1604),
.C2(n_1577),
.Y(n_1669)
);

NAND2x1p5_ASAP7_75t_L g1670 ( 
.A(n_1622),
.B(n_1360),
.Y(n_1670)
);

OAI211xp5_ASAP7_75t_SL g1671 ( 
.A1(n_1639),
.A2(n_1612),
.B(n_1577),
.C(n_1604),
.Y(n_1671)
);

OAI32xp33_ASAP7_75t_L g1672 ( 
.A1(n_1641),
.A2(n_1513),
.A3(n_1607),
.B1(n_1603),
.B2(n_1601),
.Y(n_1672)
);

AOI222xp33_ASAP7_75t_L g1673 ( 
.A1(n_1636),
.A2(n_1443),
.B1(n_1441),
.B2(n_1423),
.C1(n_1424),
.C2(n_1436),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1641),
.A2(n_1593),
.B(n_1594),
.Y(n_1674)
);

A2O1A1Ixp33_ASAP7_75t_L g1675 ( 
.A1(n_1636),
.A2(n_1613),
.B(n_1517),
.C(n_1607),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1626),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1636),
.B(n_1599),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1619),
.A2(n_1517),
.B1(n_1342),
.B2(n_1443),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1650),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1676),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1668),
.Y(n_1681)
);

NOR2x1_ASAP7_75t_L g1682 ( 
.A(n_1659),
.B(n_1631),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1667),
.B(n_1627),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1666),
.B(n_1627),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1656),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1679),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1654),
.B(n_1653),
.Y(n_1687)
);

INVx1_ASAP7_75t_SL g1688 ( 
.A(n_1665),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1658),
.Y(n_1689)
);

INVx1_ASAP7_75t_SL g1690 ( 
.A(n_1670),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1655),
.B(n_1653),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1662),
.B(n_1631),
.Y(n_1692)
);

INVxp67_ASAP7_75t_SL g1693 ( 
.A(n_1661),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1658),
.Y(n_1694)
);

OAI21xp33_ASAP7_75t_L g1695 ( 
.A1(n_1657),
.A2(n_1619),
.B(n_1646),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1677),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1660),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1663),
.Y(n_1698)
);

BUFx2_ASAP7_75t_L g1699 ( 
.A(n_1664),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1698),
.A2(n_1678),
.B1(n_1619),
.B2(n_1640),
.Y(n_1700)
);

NAND3xp33_ASAP7_75t_SL g1701 ( 
.A(n_1699),
.B(n_1662),
.C(n_1675),
.Y(n_1701)
);

NAND3xp33_ASAP7_75t_L g1702 ( 
.A(n_1689),
.B(n_1671),
.C(n_1640),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1682),
.B(n_1631),
.Y(n_1703)
);

AOI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1692),
.A2(n_1669),
.B(n_1672),
.Y(n_1704)
);

OAI21xp33_ASAP7_75t_L g1705 ( 
.A1(n_1694),
.A2(n_1619),
.B(n_1674),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1692),
.A2(n_1640),
.B(n_1649),
.Y(n_1706)
);

AOI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1693),
.A2(n_1645),
.B1(n_1618),
.B2(n_1638),
.Y(n_1707)
);

AOI211xp5_ASAP7_75t_L g1708 ( 
.A1(n_1687),
.A2(n_1638),
.B(n_1618),
.C(n_1637),
.Y(n_1708)
);

O2A1O1Ixp33_ASAP7_75t_L g1709 ( 
.A1(n_1691),
.A2(n_1649),
.B(n_1629),
.C(n_1626),
.Y(n_1709)
);

O2A1O1Ixp33_ASAP7_75t_SL g1710 ( 
.A1(n_1697),
.A2(n_1618),
.B(n_1638),
.C(n_1637),
.Y(n_1710)
);

NAND3xp33_ASAP7_75t_L g1711 ( 
.A(n_1699),
.B(n_1637),
.C(n_1629),
.Y(n_1711)
);

NOR2x1_ASAP7_75t_L g1712 ( 
.A(n_1701),
.B(n_1680),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1711),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1706),
.B(n_1685),
.Y(n_1714)
);

NOR2x1_ASAP7_75t_L g1715 ( 
.A(n_1703),
.B(n_1680),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1708),
.B(n_1697),
.Y(n_1716)
);

NOR2x1_ASAP7_75t_L g1717 ( 
.A(n_1702),
.B(n_1681),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1710),
.Y(n_1718)
);

AOI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1704),
.A2(n_1698),
.B1(n_1700),
.B2(n_1707),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1709),
.Y(n_1720)
);

NOR3x1_ASAP7_75t_L g1721 ( 
.A(n_1705),
.B(n_1686),
.C(n_1696),
.Y(n_1721)
);

NOR4xp25_ASAP7_75t_L g1722 ( 
.A(n_1713),
.B(n_1695),
.C(n_1688),
.D(n_1683),
.Y(n_1722)
);

O2A1O1Ixp5_ASAP7_75t_SL g1723 ( 
.A1(n_1718),
.A2(n_1684),
.B(n_1690),
.C(n_1632),
.Y(n_1723)
);

NOR3x1_ASAP7_75t_L g1724 ( 
.A(n_1716),
.B(n_1632),
.C(n_1644),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1715),
.Y(n_1725)
);

NAND3xp33_ASAP7_75t_SL g1726 ( 
.A(n_1719),
.B(n_1635),
.C(n_1651),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1712),
.A2(n_1635),
.B(n_1623),
.Y(n_1727)
);

AO22x1_ASAP7_75t_L g1728 ( 
.A1(n_1725),
.A2(n_1717),
.B1(n_1721),
.B2(n_1720),
.Y(n_1728)
);

AND3x4_ASAP7_75t_L g1729 ( 
.A(n_1722),
.B(n_1714),
.C(n_1623),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1727),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1724),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1726),
.Y(n_1732)
);

INVxp67_ASAP7_75t_SL g1733 ( 
.A(n_1723),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1724),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1730),
.B(n_1651),
.Y(n_1735)
);

NOR2x1p5_ASAP7_75t_L g1736 ( 
.A(n_1731),
.B(n_1297),
.Y(n_1736)
);

NOR3xp33_ASAP7_75t_L g1737 ( 
.A(n_1728),
.B(n_1297),
.C(n_1644),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1733),
.A2(n_1623),
.B(n_1652),
.Y(n_1738)
);

OAI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1730),
.A2(n_1652),
.B1(n_1673),
.B2(n_1363),
.C(n_1603),
.Y(n_1739)
);

OR3x2_ASAP7_75t_L g1740 ( 
.A(n_1736),
.B(n_1734),
.C(n_1732),
.Y(n_1740)
);

INVx2_ASAP7_75t_SL g1741 ( 
.A(n_1735),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1739),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1741),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1743),
.B(n_1738),
.Y(n_1744)
);

INVx3_ASAP7_75t_L g1745 ( 
.A(n_1744),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1744),
.A2(n_1729),
.B1(n_1740),
.B2(n_1742),
.Y(n_1746)
);

OR2x6_ASAP7_75t_L g1747 ( 
.A(n_1745),
.B(n_1737),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1746),
.A2(n_1623),
.B1(n_1441),
.B2(n_1313),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1747),
.B(n_1599),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1748),
.A2(n_1594),
.B1(n_1363),
.B2(n_1381),
.Y(n_1750)
);

AOI222xp33_ASAP7_75t_SL g1751 ( 
.A1(n_1749),
.A2(n_1750),
.B1(n_1521),
.B2(n_1525),
.C1(n_1516),
.C2(n_1518),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1751),
.A2(n_1381),
.B1(n_1317),
.B2(n_1394),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1752),
.A2(n_1342),
.B1(n_1381),
.B2(n_1505),
.Y(n_1753)
);

AOI211xp5_ASAP7_75t_L g1754 ( 
.A1(n_1753),
.A2(n_1379),
.B(n_1416),
.C(n_1479),
.Y(n_1754)
);


endmodule