module fake_jpeg_17136_n_291 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_291);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_291;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_24),
.B(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_30),
.B1(n_33),
.B2(n_17),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_23),
.B1(n_34),
.B2(n_31),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_23),
.B1(n_34),
.B2(n_31),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_23),
.B1(n_34),
.B2(n_35),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_35),
.B1(n_26),
.B2(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_62),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_35),
.B1(n_26),
.B2(n_32),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_63),
.B1(n_30),
.B2(n_28),
.Y(n_77)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_20),
.B1(n_32),
.B2(n_21),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_24),
.B(n_40),
.C(n_37),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_85),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_49),
.A2(n_33),
.B1(n_19),
.B2(n_17),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_65),
.A2(n_61),
.B1(n_54),
.B2(n_29),
.Y(n_112)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_66),
.B(n_67),
.Y(n_124)
);

CKINVDCx12_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_59),
.A2(n_43),
.B1(n_39),
.B2(n_38),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_68),
.A2(n_74),
.B1(n_90),
.B2(n_83),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_42),
.B1(n_44),
.B2(n_39),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_70),
.A2(n_77),
.B1(n_79),
.B2(n_93),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_42),
.B1(n_50),
.B2(n_44),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_71),
.A2(n_88),
.B1(n_94),
.B2(n_55),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_57),
.A2(n_44),
.B1(n_43),
.B2(n_38),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_72),
.A2(n_81),
.B1(n_41),
.B2(n_29),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_48),
.B(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_76),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_19),
.C(n_22),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_96),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_39),
.B1(n_38),
.B2(n_43),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_18),
.B1(n_29),
.B2(n_39),
.Y(n_81)
);

XOR2x2_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_43),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_0),
.C(n_1),
.Y(n_130)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_22),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_22),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_92),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_43),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_21),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_91),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_61),
.B(n_28),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_22),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_54),
.B1(n_58),
.B2(n_53),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_39),
.B1(n_38),
.B2(n_43),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

CKINVDCx12_ASAP7_75t_R g97 ( 
.A(n_61),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_97),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_60),
.B(n_25),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_98),
.B(n_99),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_22),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_25),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_100),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_54),
.B(n_25),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_61),
.B(n_10),
.Y(n_102)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_112),
.A2(n_113),
.B1(n_122),
.B2(n_95),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_66),
.A2(n_38),
.B1(n_41),
.B2(n_29),
.Y(n_113)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_88),
.B1(n_69),
.B2(n_94),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_119),
.A2(n_95),
.B1(n_87),
.B2(n_3),
.Y(n_159)
);

NAND2xp33_ASAP7_75t_SL g120 ( 
.A(n_71),
.B(n_41),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_130),
.B(n_98),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_70),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

NOR2x1_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_76),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_132),
.A2(n_137),
.B(n_141),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_85),
.C(n_86),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_138),
.C(n_145),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_106),
.B(n_82),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_136),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_82),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_64),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_111),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_110),
.B(n_73),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_140),
.B(n_149),
.Y(n_163)
);

NOR2xp67_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_75),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_SL g173 ( 
.A1(n_144),
.A2(n_158),
.B(n_103),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_92),
.C(n_72),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_88),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_150),
.B(n_153),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_68),
.B(n_1),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_0),
.B(n_1),
.Y(n_165)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_68),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_68),
.B1(n_90),
.B2(n_96),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_160),
.B1(n_105),
.B2(n_109),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_79),
.Y(n_155)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_125),
.B(n_108),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_93),
.Y(n_157)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_9),
.B(n_15),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_126),
.B1(n_121),
.B2(n_108),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_164),
.A2(n_174),
.B1(n_175),
.B2(n_179),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_165),
.A2(n_177),
.B1(n_189),
.B2(n_147),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_119),
.C(n_130),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_167),
.B(n_176),
.C(n_182),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_120),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_168),
.B(n_185),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_173),
.A2(n_187),
.B1(n_152),
.B2(n_139),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_117),
.B1(n_122),
.B2(n_103),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_154),
.A2(n_117),
.B1(n_115),
.B2(n_109),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_117),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_178),
.B(n_181),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_141),
.A2(n_117),
.B1(n_107),
.B2(n_123),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_123),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_104),
.C(n_87),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_183),
.B(n_184),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_137),
.B(n_114),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_134),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_186),
.B(n_148),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_144),
.A2(n_105),
.B1(n_114),
.B2(n_104),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_132),
.A2(n_0),
.B(n_1),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_166),
.Y(n_191)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_132),
.Y(n_192)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_136),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_202),
.C(n_167),
.Y(n_214)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_198),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_135),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_206),
.Y(n_228)
);

AOI322xp5_ASAP7_75t_SL g200 ( 
.A1(n_180),
.A2(n_156),
.A3(n_143),
.B1(n_140),
.B2(n_159),
.C1(n_151),
.C2(n_157),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_200),
.B(n_203),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_155),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_143),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_222)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_184),
.Y(n_226)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_216),
.C(n_223),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_162),
.C(n_168),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_192),
.A2(n_180),
.B(n_189),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_207),
.B1(n_199),
.B2(n_197),
.Y(n_236)
);

NAND2x1_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_179),
.Y(n_221)
);

BUFx12f_ASAP7_75t_SL g238 ( 
.A(n_221),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_185),
.C(n_172),
.Y(n_223)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

XNOR2x1_ASAP7_75t_SL g227 ( 
.A(n_190),
.B(n_165),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_227),
.A2(n_231),
.B1(n_3),
.B2(n_4),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_196),
.C(n_195),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_190),
.C(n_204),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_212),
.A2(n_210),
.B1(n_209),
.B2(n_204),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_245),
.C(n_223),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_211),
.Y(n_235)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_248),
.B1(n_226),
.B2(n_228),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_228),
.B(n_193),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_237),
.B(n_242),
.Y(n_250)
);

AOI322xp5_ASAP7_75t_L g239 ( 
.A1(n_230),
.A2(n_191),
.A3(n_201),
.B1(n_194),
.B2(n_148),
.C1(n_104),
.C2(n_8),
.Y(n_239)
);

BUFx24_ASAP7_75t_SL g258 ( 
.A(n_239),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_243),
.B1(n_220),
.B2(n_14),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_9),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_222),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_7),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_244),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_11),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_217),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_249),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_225),
.B1(n_218),
.B2(n_224),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_221),
.B1(n_225),
.B2(n_224),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_260),
.B1(n_261),
.B2(n_246),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_238),
.A2(n_227),
.B1(n_222),
.B2(n_231),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_259),
.Y(n_271)
);

XNOR2x1_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_216),
.Y(n_254)
);

AO22x1_ASAP7_75t_L g270 ( 
.A1(n_254),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_270)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_240),
.A2(n_229),
.B1(n_4),
.B2(n_5),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_3),
.C(n_4),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_245),
.C(n_234),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_257),
.B(n_247),
.Y(n_263)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_266),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_265),
.B(n_267),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_233),
.C(n_254),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_247),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_248),
.C(n_236),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_268),
.B(n_256),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_270),
.A2(n_253),
.B(n_250),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_274),
.B(n_268),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_271),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g277 ( 
.A1(n_269),
.A2(n_258),
.B(n_261),
.Y(n_277)
);

OAI211xp5_ASAP7_75t_L g281 ( 
.A1(n_277),
.A2(n_278),
.B(n_265),
.C(n_266),
.Y(n_281)
);

NOR2x1_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_251),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_11),
.C(n_12),
.Y(n_285)
);

AOI322xp5_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_281),
.A3(n_282),
.B1(n_283),
.B2(n_274),
.C1(n_272),
.C2(n_273),
.Y(n_284)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_278),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_275),
.B(n_11),
.Y(n_283)
);

A2O1A1Ixp33_ASAP7_75t_SL g287 ( 
.A1(n_284),
.A2(n_6),
.B(n_263),
.C(n_283),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_286),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_281),
.A2(n_12),
.B(n_15),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_287),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_288),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_6),
.Y(n_291)
);


endmodule