module real_aes_8691_n_382 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_382);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_382;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_618;
wire n_1170;
wire n_778;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_1110;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_1014;
wire n_421;
wire n_742;
wire n_852;
wire n_555;
wire n_766;
wire n_974;
wire n_1113;
wire n_919;
wire n_1089;
wire n_857;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_1034;
wire n_571;
wire n_491;
wire n_894;
wire n_694;
wire n_1123;
wire n_923;
wire n_952;
wire n_429;
wire n_1166;
wire n_1137;
wire n_752;
wire n_556;
wire n_448;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_666;
wire n_537;
wire n_884;
wire n_551;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_1146;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_958;
wire n_677;
wire n_1021;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_961;
wire n_870;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_1160;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_892;
wire n_495;
wire n_1078;
wire n_994;
wire n_1072;
wire n_384;
wire n_744;
wire n_938;
wire n_1128;
wire n_935;
wire n_1098;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_559;
wire n_1049;
wire n_636;
wire n_466;
wire n_976;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_1070;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_1168;
wire n_755;
wire n_1025;
wire n_1148;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_996;
wire n_860;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_1152;
wire n_801;
wire n_1126;
wire n_383;
wire n_529;
wire n_1115;
wire n_455;
wire n_725;
wire n_504;
wire n_973;
wire n_1081;
wire n_671;
wire n_960;
wire n_1084;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_1017;
wire n_1013;
wire n_737;
wire n_936;
wire n_581;
wire n_610;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_1135;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_398;
wire n_1167;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1103;
wire n_1131;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_1145;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_1077;
wire n_501;
wire n_488;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_1163;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_756;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_1171;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1157;
wire n_1158;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_1136;
wire n_579;
wire n_1033;
wire n_533;
wire n_699;
wire n_1028;
wire n_1003;
wire n_1000;
wire n_727;
wire n_1083;
wire n_397;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_1155;
wire n_1165;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1169;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_1043;
wire n_850;
wire n_720;
wire n_1127;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_1068;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_691;
wire n_765;
wire n_481;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_679;
wire n_520;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_1071;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_1133;
wire n_1164;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_1162;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_639;
wire n_587;
wire n_1010;
wire n_811;
wire n_823;
wire n_459;
wire n_558;
wire n_1015;
wire n_1172;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1150;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_929;
wire n_1143;
wire n_686;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_949;
wire n_507;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_1045;
wire n_1114;
wire n_465;
wire n_473;
wire n_566;
wire n_837;
wire n_967;
wire n_719;
wire n_871;
wire n_474;
wire n_1159;
wire n_1156;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1151;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_968;
wire n_710;
wire n_650;
wire n_743;
wire n_646;
wire n_1040;
wire n_652;
wire n_1097;
wire n_393;
wire n_601;
wire n_500;
wire n_1102;
wire n_661;
wire n_463;
wire n_703;
wire n_396;
wire n_804;
wire n_1076;
wire n_447;
wire n_1101;
wire n_1173;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_1119;
wire n_1039;
wire n_868;
wire n_802;
wire n_877;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_0), .A2(n_288), .B1(n_596), .B2(n_705), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g952 ( .A(n_1), .Y(n_952) );
CKINVDCx20_ASAP7_75t_R g1077 ( .A(n_2), .Y(n_1077) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_3), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_4), .A2(n_54), .B1(n_521), .B2(n_524), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g1024 ( .A(n_5), .Y(n_1024) );
AOI221xp5_ASAP7_75t_L g564 ( .A1(n_6), .A2(n_14), .B1(n_565), .B2(n_567), .C(n_568), .Y(n_564) );
AOI221xp5_ASAP7_75t_L g545 ( .A1(n_7), .A2(n_272), .B1(n_546), .B2(n_548), .C(n_549), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g1131 ( .A1(n_8), .A2(n_141), .B1(n_587), .B2(n_919), .Y(n_1131) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_9), .Y(n_814) );
AO22x2_ASAP7_75t_L g402 ( .A1(n_10), .A2(n_224), .B1(n_403), .B2(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g1110 ( .A(n_10), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_11), .A2(n_158), .B1(n_455), .B2(n_774), .Y(n_939) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_12), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g902 ( .A(n_13), .Y(n_902) );
CKINVDCx20_ASAP7_75t_R g955 ( .A(n_15), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_16), .A2(n_291), .B1(n_638), .B2(n_652), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g887 ( .A(n_17), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_18), .A2(n_108), .B1(n_455), .B2(n_772), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_19), .A2(n_57), .B1(n_427), .B2(n_528), .Y(n_871) );
CKINVDCx20_ASAP7_75t_R g1034 ( .A(n_20), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_21), .A2(n_249), .B1(n_943), .B2(n_944), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1125 ( .A(n_22), .B(n_608), .Y(n_1125) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_23), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_24), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g931 ( .A(n_25), .Y(n_931) );
AOI222xp33_ASAP7_75t_L g669 ( .A1(n_26), .A2(n_59), .B1(n_341), .B2(n_575), .C1(n_577), .C2(n_670), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g1042 ( .A(n_27), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_28), .A2(n_128), .B1(n_479), .B2(n_763), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_29), .A2(n_58), .B1(n_485), .B2(n_776), .Y(n_1009) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_30), .Y(n_751) );
AO22x2_ASAP7_75t_L g406 ( .A1(n_31), .A2(n_115), .B1(n_403), .B2(n_407), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_32), .A2(n_544), .B1(n_579), .B2(n_580), .Y(n_543) );
INVx1_ASAP7_75t_L g579 ( .A(n_32), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_33), .A2(n_373), .B1(n_636), .B2(n_834), .Y(n_833) );
AOI22xp5_ASAP7_75t_L g1016 ( .A1(n_34), .A2(n_1017), .B1(n_1045), .B2(n_1046), .Y(n_1016) );
CKINVDCx20_ASAP7_75t_R g1045 ( .A(n_34), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_35), .A2(n_250), .B1(n_479), .B2(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_SL g1151 ( .A1(n_36), .A2(n_96), .B1(n_427), .B2(n_436), .Y(n_1151) );
INVx1_ASAP7_75t_L g440 ( .A(n_37), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_38), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_39), .A2(n_120), .B1(n_456), .B2(n_487), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_40), .A2(n_160), .B1(n_498), .B2(n_499), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g918 ( .A1(n_41), .A2(n_276), .B1(n_831), .B2(n_919), .Y(n_918) );
CKINVDCx20_ASAP7_75t_R g1124 ( .A(n_42), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_43), .B(n_567), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_44), .B(n_525), .Y(n_1002) );
CKINVDCx20_ASAP7_75t_R g1005 ( .A(n_45), .Y(n_1005) );
AOI22xp5_ASAP7_75t_SL g708 ( .A1(n_46), .A2(n_709), .B1(n_710), .B2(n_733), .Y(n_708) );
INVx1_ASAP7_75t_L g733 ( .A(n_46), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g1004 ( .A(n_47), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_48), .A2(n_189), .B1(n_455), .B2(n_664), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_49), .A2(n_332), .B1(n_474), .B2(n_477), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g932 ( .A1(n_50), .A2(n_217), .B1(n_428), .B2(n_578), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_51), .A2(n_248), .B1(n_499), .B2(n_728), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g951 ( .A(n_52), .Y(n_951) );
CKINVDCx20_ASAP7_75t_R g893 ( .A(n_53), .Y(n_893) );
CKINVDCx20_ASAP7_75t_R g1001 ( .A(n_55), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_56), .A2(n_129), .B1(n_779), .B2(n_780), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_60), .A2(n_148), .B1(n_467), .B2(n_501), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_61), .A2(n_247), .B1(n_943), .B2(n_944), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_62), .A2(n_289), .B1(n_482), .B2(n_1136), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_63), .A2(n_112), .B1(n_591), .B2(n_593), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_64), .A2(n_315), .B1(n_501), .B2(n_503), .Y(n_500) );
AOI22xp33_ASAP7_75t_SL g1064 ( .A1(n_65), .A2(n_275), .B1(n_502), .B2(n_868), .Y(n_1064) );
CKINVDCx20_ASAP7_75t_R g1080 ( .A(n_66), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_67), .A2(n_343), .B1(n_943), .B2(n_944), .Y(n_1011) );
CKINVDCx20_ASAP7_75t_R g910 ( .A(n_68), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_69), .A2(n_298), .B1(n_482), .B2(n_486), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_70), .Y(n_413) );
INVx1_ASAP7_75t_L g972 ( .A(n_71), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_72), .A2(n_355), .B1(n_501), .B2(n_650), .Y(n_866) );
CKINVDCx20_ASAP7_75t_R g1028 ( .A(n_73), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_74), .A2(n_106), .B1(n_479), .B2(n_813), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_75), .A2(n_340), .B1(n_501), .B2(n_785), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_76), .A2(n_100), .B1(n_758), .B2(n_760), .Y(n_757) );
AOI222xp33_ASAP7_75t_L g911 ( .A1(n_77), .A2(n_282), .B1(n_339), .B2(n_521), .C1(n_575), .C2(n_608), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_78), .B(n_524), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_79), .A2(n_292), .B1(n_666), .B2(n_668), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_80), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g847 ( .A1(n_81), .A2(n_214), .B1(n_436), .B2(n_670), .Y(n_847) );
INVx1_ASAP7_75t_L g915 ( .A(n_82), .Y(n_915) );
CKINVDCx20_ASAP7_75t_R g1036 ( .A(n_83), .Y(n_1036) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_84), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_85), .A2(n_210), .B1(n_587), .B2(n_588), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_86), .A2(n_136), .B1(n_537), .B2(n_540), .Y(n_536) );
AO22x2_ASAP7_75t_L g410 ( .A1(n_87), .A2(n_254), .B1(n_403), .B2(n_404), .Y(n_410) );
INVx1_ASAP7_75t_L g1107 ( .A(n_87), .Y(n_1107) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_88), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_89), .A2(n_90), .B1(n_638), .B2(n_668), .Y(n_1088) );
AOI22xp33_ASAP7_75t_SL g1160 ( .A1(n_91), .A2(n_312), .B1(n_1161), .B2(n_1162), .Y(n_1160) );
AOI22xp5_ASAP7_75t_L g922 ( .A1(n_92), .A2(n_113), .B1(n_642), .B2(n_765), .Y(n_922) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_93), .A2(n_231), .B1(n_437), .B2(n_625), .Y(n_694) );
AOI22x1_ASAP7_75t_L g991 ( .A1(n_94), .A2(n_992), .B1(n_1013), .B2(n_1014), .Y(n_991) );
INVx1_ASAP7_75t_L g1013 ( .A(n_94), .Y(n_1013) );
AOI222xp33_ASAP7_75t_L g574 ( .A1(n_95), .A2(n_109), .B1(n_139), .B2(n_427), .C1(n_575), .C2(n_577), .Y(n_574) );
CKINVDCx20_ASAP7_75t_R g822 ( .A(n_97), .Y(n_822) );
AOI211xp5_ASAP7_75t_L g1164 ( .A1(n_98), .A2(n_728), .B(n_1165), .C(n_1169), .Y(n_1164) );
AOI22xp33_ASAP7_75t_SL g1153 ( .A1(n_99), .A2(n_284), .B1(n_1154), .B2(n_1155), .Y(n_1153) );
INVx1_ASAP7_75t_L g957 ( .A(n_101), .Y(n_957) );
AOI221xp5_ASAP7_75t_L g907 ( .A1(n_102), .A2(n_327), .B1(n_628), .B2(n_630), .C(n_908), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_103), .A2(n_146), .B1(n_532), .B2(n_716), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g1081 ( .A(n_104), .Y(n_1081) );
CKINVDCx20_ASAP7_75t_R g1075 ( .A(n_105), .Y(n_1075) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_107), .A2(n_183), .B1(n_660), .B2(n_661), .Y(n_659) );
AOI22xp33_ASAP7_75t_SL g723 ( .A1(n_110), .A2(n_358), .B1(n_724), .B2(n_725), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_111), .A2(n_364), .B1(n_728), .B2(n_756), .Y(n_874) );
CKINVDCx20_ASAP7_75t_R g995 ( .A(n_114), .Y(n_995) );
INVx1_ASAP7_75t_L g1111 ( .A(n_115), .Y(n_1111) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_116), .Y(n_519) );
AOI22xp33_ASAP7_75t_SL g719 ( .A1(n_117), .A2(n_166), .B1(n_633), .B2(n_660), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g926 ( .A(n_118), .Y(n_926) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_119), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g889 ( .A(n_121), .Y(n_889) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_122), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g1033 ( .A(n_123), .Y(n_1033) );
CKINVDCx20_ASAP7_75t_R g1053 ( .A(n_124), .Y(n_1053) );
AOI22xp5_ASAP7_75t_L g1113 ( .A1(n_125), .A2(n_1114), .B1(n_1115), .B2(n_1137), .Y(n_1113) );
CKINVDCx20_ASAP7_75t_R g1137 ( .A(n_125), .Y(n_1137) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_126), .B(n_608), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_127), .A2(n_293), .B1(n_455), .B2(n_763), .Y(n_1008) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_130), .A2(n_303), .B1(n_459), .B2(n_479), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_131), .A2(n_212), .B1(n_784), .B2(n_785), .Y(n_783) );
AOI22xp33_ASAP7_75t_SL g632 ( .A1(n_132), .A2(n_178), .B1(n_523), .B2(n_633), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_133), .Y(n_816) );
AOI22xp33_ASAP7_75t_SL g637 ( .A1(n_134), .A2(n_299), .B1(n_638), .B2(n_639), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_135), .A2(n_331), .B1(n_437), .B2(n_633), .Y(n_1078) );
CKINVDCx20_ASAP7_75t_R g1128 ( .A(n_137), .Y(n_1128) );
AOI22xp33_ASAP7_75t_SL g1060 ( .A1(n_138), .A2(n_322), .B1(n_625), .B2(n_661), .Y(n_1060) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_140), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_142), .A2(n_328), .B1(n_462), .B2(n_650), .Y(n_649) );
AOI222xp33_ASAP7_75t_L g875 ( .A1(n_143), .A2(n_225), .B1(n_307), .B2(n_421), .C1(n_534), .C2(n_876), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_144), .A2(n_204), .B1(n_774), .B2(n_861), .Y(n_860) );
CKINVDCx20_ASAP7_75t_R g925 ( .A(n_145), .Y(n_925) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_147), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_149), .B(n_1057), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_150), .A2(n_203), .B1(n_756), .B2(n_831), .Y(n_830) );
AND2x6_ASAP7_75t_L g385 ( .A(n_151), .B(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g1104 ( .A(n_151), .Y(n_1104) );
AOI22xp33_ASAP7_75t_SL g527 ( .A1(n_152), .A2(n_277), .B1(n_528), .B2(n_532), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_153), .A2(n_176), .B1(n_666), .B2(n_835), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_154), .A2(n_265), .B1(n_605), .B2(n_765), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_155), .A2(n_279), .B1(n_467), .B2(n_834), .Y(n_1012) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_156), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_157), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_159), .A2(n_185), .B1(n_782), .B2(n_856), .Y(n_855) );
AOI22xp5_ASAP7_75t_SL g963 ( .A1(n_161), .A2(n_964), .B1(n_985), .B2(n_986), .Y(n_963) );
INVx1_ASAP7_75t_L g986 ( .A(n_161), .Y(n_986) );
AOI22xp33_ASAP7_75t_SL g1054 ( .A1(n_162), .A2(n_281), .B1(n_578), .B2(n_852), .Y(n_1054) );
AOI22xp5_ASAP7_75t_L g920 ( .A1(n_163), .A2(n_302), .B1(n_835), .B2(n_861), .Y(n_920) );
NAND2xp5_ASAP7_75t_SL g629 ( .A(n_164), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g967 ( .A(n_165), .Y(n_967) );
AOI22xp33_ASAP7_75t_SL g1156 ( .A1(n_167), .A2(n_236), .B1(n_628), .B2(n_631), .Y(n_1156) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_168), .Y(n_610) );
AO22x2_ASAP7_75t_L g412 ( .A1(n_169), .A2(n_245), .B1(n_403), .B2(n_407), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g1108 ( .A(n_169), .B(n_1109), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_170), .A2(n_180), .B1(n_462), .B2(n_467), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g1170 ( .A(n_171), .Y(n_1170) );
AOI22xp33_ASAP7_75t_SL g643 ( .A1(n_172), .A2(n_261), .B1(n_499), .B2(n_644), .Y(n_643) );
AOI22xp33_ASAP7_75t_SL g1158 ( .A1(n_173), .A2(n_262), .B1(n_765), .B2(n_1159), .Y(n_1158) );
XNOR2x2_ASAP7_75t_L g863 ( .A(n_174), .B(n_864), .Y(n_863) );
CKINVDCx20_ASAP7_75t_R g897 ( .A(n_175), .Y(n_897) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_177), .A2(n_269), .B1(n_436), .B2(n_625), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g999 ( .A(n_179), .Y(n_999) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_181), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_182), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_184), .A2(n_316), .B1(n_774), .B2(n_868), .Y(n_867) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_186), .Y(n_689) );
AOI22xp33_ASAP7_75t_SL g641 ( .A1(n_187), .A2(n_202), .B1(n_588), .B2(n_642), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g923 ( .A1(n_188), .A2(n_234), .B1(n_638), .B2(n_702), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_190), .A2(n_228), .B1(n_537), .B2(n_540), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_191), .A2(n_394), .B1(n_490), .B2(n_491), .Y(n_393) );
INVx1_ASAP7_75t_L g490 ( .A(n_191), .Y(n_490) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_192), .A2(n_360), .B1(n_650), .B2(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g714 ( .A(n_193), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_194), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_195), .A2(n_311), .B1(n_467), .B2(n_834), .Y(n_945) );
CKINVDCx20_ASAP7_75t_R g1120 ( .A(n_196), .Y(n_1120) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_197), .B(n_1040), .Y(n_1039) );
CKINVDCx20_ASAP7_75t_R g1150 ( .A(n_198), .Y(n_1150) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_199), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g671 ( .A(n_200), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_201), .A2(n_367), .B1(n_638), .B2(n_652), .Y(n_651) );
AOI22xp33_ASAP7_75t_SL g635 ( .A1(n_205), .A2(n_354), .B1(n_462), .B2(n_636), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_206), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_207), .B(n_608), .Y(n_953) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_208), .Y(n_819) );
AOI22xp33_ASAP7_75t_SL g1063 ( .A1(n_209), .A2(n_258), .B1(n_479), .B2(n_666), .Y(n_1063) );
CKINVDCx20_ASAP7_75t_R g949 ( .A(n_211), .Y(n_949) );
INVxp67_ASAP7_75t_L g1145 ( .A(n_213), .Y(n_1145) );
XNOR2xp5_ASAP7_75t_L g1146 ( .A(n_213), .B(n_1147), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_215), .A2(n_223), .B1(n_436), .B2(n_748), .Y(n_747) );
AOI211xp5_ASAP7_75t_L g382 ( .A1(n_216), .A2(n_383), .B(n_391), .C(n_1112), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g899 ( .A(n_218), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_219), .A2(n_257), .B1(n_588), .B2(n_668), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_220), .A2(n_226), .B1(n_477), .B2(n_596), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g909 ( .A(n_221), .Y(n_909) );
CKINVDCx20_ASAP7_75t_R g1122 ( .A(n_222), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_227), .A2(n_346), .B1(n_592), .B2(n_983), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_229), .B(n_1168), .Y(n_1167) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_230), .A2(n_320), .B1(n_638), .B2(n_652), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g600 ( .A(n_232), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_233), .A2(n_274), .B1(n_779), .B2(n_780), .Y(n_984) );
OA22x2_ASAP7_75t_L g1069 ( .A1(n_235), .A2(n_1070), .B1(n_1071), .B2(n_1089), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_235), .Y(n_1070) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_237), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g996 ( .A(n_238), .Y(n_996) );
CKINVDCx20_ASAP7_75t_R g1043 ( .A(n_239), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_240), .B(n_628), .Y(n_627) );
XNOR2x2_ASAP7_75t_L g493 ( .A(n_241), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g390 ( .A(n_242), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g935 ( .A1(n_243), .A2(n_936), .B1(n_958), .B2(n_959), .Y(n_935) );
INVx1_ASAP7_75t_L g958 ( .A(n_243), .Y(n_958) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_244), .Y(n_799) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_246), .A2(n_256), .B1(n_482), .B2(n_763), .Y(n_762) );
AOI22xp33_ASAP7_75t_SL g1067 ( .A1(n_251), .A2(n_375), .B1(n_485), .B2(n_702), .Y(n_1067) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_252), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g1066 ( .A1(n_253), .A2(n_370), .B1(n_474), .B2(n_919), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_255), .A2(n_347), .B1(n_530), .B2(n_852), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g1026 ( .A(n_259), .Y(n_1026) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_260), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g1038 ( .A(n_263), .Y(n_1038) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_264), .A2(n_583), .B1(n_615), .B2(n_616), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g615 ( .A(n_264), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_266), .A2(n_365), .B1(n_462), .B2(n_785), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_267), .A2(n_372), .B1(n_644), .B2(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_268), .B(n_658), .Y(n_849) );
AOI22xp5_ASAP7_75t_L g883 ( .A1(n_270), .A2(n_884), .B1(n_912), .B2(n_913), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g912 ( .A(n_270), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_271), .A2(n_351), .B1(n_503), .B2(n_1022), .Y(n_1021) );
CKINVDCx20_ASAP7_75t_R g1074 ( .A(n_273), .Y(n_1074) );
INVx1_ASAP7_75t_L g971 ( .A(n_278), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_280), .A2(n_300), .B1(n_639), .B2(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g975 ( .A(n_283), .Y(n_975) );
INVx1_ASAP7_75t_L g403 ( .A(n_285), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_285), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_286), .A2(n_369), .B1(n_479), .B2(n_765), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_287), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_290), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g555 ( .A1(n_294), .A2(n_306), .B1(n_482), .B2(n_556), .C(n_559), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g905 ( .A(n_295), .Y(n_905) );
CKINVDCx20_ASAP7_75t_R g838 ( .A(n_296), .Y(n_838) );
INVx1_ASAP7_75t_L g948 ( .A(n_297), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_301), .B(n_658), .Y(n_657) );
AOI22xp33_ASAP7_75t_SL g859 ( .A1(n_304), .A2(n_363), .B1(n_596), .B2(n_705), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_305), .A2(n_326), .B1(n_455), .B2(n_459), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_308), .A2(n_353), .B1(n_666), .B2(n_702), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_309), .A2(n_338), .B1(n_530), .B2(n_534), .Y(n_927) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_310), .Y(n_434) );
AND2x2_ASAP7_75t_L g389 ( .A(n_313), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g445 ( .A(n_314), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_317), .Y(n_645) );
INVx1_ASAP7_75t_L g386 ( .A(n_318), .Y(n_386) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_319), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_321), .Y(n_560) );
OA22x2_ASAP7_75t_L g1048 ( .A1(n_323), .A2(n_1049), .B1(n_1050), .B2(n_1068), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_323), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_324), .A2(n_359), .B1(n_587), .B2(n_668), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_325), .B(n_631), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_329), .A2(n_333), .B1(n_537), .B2(n_540), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_330), .A2(n_342), .B1(n_588), .B2(n_782), .Y(n_873) );
CKINVDCx20_ASAP7_75t_R g613 ( .A(n_334), .Y(n_613) );
CKINVDCx20_ASAP7_75t_R g1029 ( .A(n_335), .Y(n_1029) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_336), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_337), .B(n_524), .Y(n_973) );
CKINVDCx20_ASAP7_75t_R g846 ( .A(n_344), .Y(n_846) );
INVx1_ASAP7_75t_L g766 ( .A(n_345), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g1119 ( .A(n_348), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_349), .B(n_532), .Y(n_817) );
INVx1_ASAP7_75t_L g969 ( .A(n_350), .Y(n_969) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_352), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g1166 ( .A(n_356), .Y(n_1166) );
CKINVDCx20_ASAP7_75t_R g603 ( .A(n_357), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g892 ( .A(n_361), .Y(n_892) );
INVx1_ASAP7_75t_L g707 ( .A(n_362), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_366), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_368), .B(n_436), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_371), .Y(n_788) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_374), .A2(n_768), .B1(n_800), .B2(n_801), .Y(n_767) );
INVx1_ASAP7_75t_L g800 ( .A(n_374), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_376), .Y(n_397) );
CKINVDCx20_ASAP7_75t_R g1127 ( .A(n_377), .Y(n_1127) );
INVx1_ASAP7_75t_L g976 ( .A(n_378), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_379), .A2(n_381), .B1(n_774), .B2(n_776), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_380), .Y(n_425) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
HB1xp67_ASAP7_75t_L g1103 ( .A(n_386), .Y(n_1103) );
OAI21xp5_ASAP7_75t_L g1143 ( .A1(n_387), .A2(n_1102), .B(n_1144), .Y(n_1143) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_388), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_679), .B1(n_1097), .B2(n_1098), .C(n_1099), .Y(n_391) );
INVxp67_ASAP7_75t_L g1097 ( .A(n_392), .Y(n_1097) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_492), .B1(n_677), .B2(n_678), .Y(n_392) );
INVx1_ASAP7_75t_L g677 ( .A(n_393), .Y(n_677) );
INVx2_ASAP7_75t_L g491 ( .A(n_394), .Y(n_491) );
AND2x2_ASAP7_75t_SL g394 ( .A(n_395), .B(n_452), .Y(n_394) );
NOR3xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_419), .C(n_439), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B1(n_413), .B2(n_414), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_398), .A2(n_689), .B1(n_690), .B2(n_691), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_398), .A2(n_655), .B1(n_1074), .B2(n_1075), .Y(n_1073) );
BUFx3_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g612 ( .A(n_399), .Y(n_612) );
BUFx6f_ASAP7_75t_L g789 ( .A(n_399), .Y(n_789) );
OAI221xp5_ASAP7_75t_L g924 ( .A1(n_399), .A2(n_416), .B1(n_925), .B2(n_926), .C(n_927), .Y(n_924) );
OR2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_408), .Y(n_399) );
INVx2_ASAP7_75t_L g460 ( .A(n_400), .Y(n_460) );
OR2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_406), .Y(n_400) );
AND2x2_ASAP7_75t_L g418 ( .A(n_401), .B(n_406), .Y(n_418) );
AND2x2_ASAP7_75t_L g458 ( .A(n_401), .B(n_432), .Y(n_458) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g422 ( .A(n_402), .B(n_406), .Y(n_422) );
AND2x2_ASAP7_75t_L g433 ( .A(n_402), .B(n_412), .Y(n_433) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_405), .Y(n_407) );
INVx2_ASAP7_75t_L g432 ( .A(n_406), .Y(n_432) );
INVx1_ASAP7_75t_L g470 ( .A(n_406), .Y(n_470) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND2x1p5_ASAP7_75t_L g417 ( .A(n_409), .B(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g485 ( .A(n_409), .B(n_458), .Y(n_485) );
AND2x4_ASAP7_75t_L g539 ( .A(n_409), .B(n_460), .Y(n_539) );
AND2x6_ASAP7_75t_L g541 ( .A(n_409), .B(n_418), .Y(n_541) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g424 ( .A(n_410), .Y(n_424) );
INVx1_ASAP7_75t_L g431 ( .A(n_410), .Y(n_431) );
INVx1_ASAP7_75t_L g451 ( .A(n_410), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_410), .B(n_412), .Y(n_471) );
AND2x2_ASAP7_75t_L g423 ( .A(n_411), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g466 ( .A(n_412), .B(n_451), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_414), .A2(n_611), .B1(n_742), .B2(n_743), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_414), .A2(n_819), .B1(n_820), .B2(n_822), .Y(n_818) );
OAI22xp5_ASAP7_75t_L g1118 ( .A1(n_414), .A2(n_968), .B1(n_1119), .B2(n_1120), .Y(n_1118) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx3_ASAP7_75t_L g614 ( .A(n_416), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g947 ( .A1(n_416), .A2(n_789), .B1(n_948), .B2(n_949), .Y(n_947) );
BUFx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g656 ( .A(n_417), .Y(n_656) );
AND2x2_ASAP7_75t_L g465 ( .A(n_418), .B(n_466), .Y(n_465) );
AND2x4_ASAP7_75t_L g476 ( .A(n_418), .B(n_423), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_418), .B(n_466), .Y(n_552) );
OAI221xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_425), .B1(n_426), .B2(n_434), .C(n_435), .Y(n_419) );
OAI221xp5_ASAP7_75t_SL g602 ( .A1(n_420), .A2(n_603), .B1(n_604), .B2(n_606), .C(n_607), .Y(n_602) );
OAI21xp5_ASAP7_75t_SL g622 ( .A1(n_420), .A2(n_623), .B(n_624), .Y(n_622) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g518 ( .A(n_421), .Y(n_518) );
INVx4_ASAP7_75t_L g576 ( .A(n_421), .Y(n_576) );
BUFx6f_ASAP7_75t_L g813 ( .A(n_421), .Y(n_813) );
BUFx3_ASAP7_75t_L g930 ( .A(n_421), .Y(n_930) );
AND2x6_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g448 ( .A(n_422), .Y(n_448) );
AND2x4_ASAP7_75t_L g535 ( .A(n_422), .B(n_450), .Y(n_535) );
AND2x2_ASAP7_75t_L g457 ( .A(n_423), .B(n_458), .Y(n_457) );
AND2x6_ASAP7_75t_L g459 ( .A(n_423), .B(n_460), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_426), .A2(n_443), .B1(n_696), .B2(n_697), .Y(n_695) );
INVx2_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_SL g1037 ( .A(n_427), .Y(n_1037) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g825 ( .A(n_428), .Y(n_825) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_429), .Y(n_523) );
BUFx2_ASAP7_75t_L g605 ( .A(n_429), .Y(n_605) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_429), .Y(n_660) );
BUFx4f_ASAP7_75t_SL g852 ( .A(n_429), .Y(n_852) );
AND2x4_ASAP7_75t_L g429 ( .A(n_430), .B(n_433), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_L g438 ( .A(n_431), .Y(n_438) );
INVx1_ASAP7_75t_L g444 ( .A(n_432), .Y(n_444) );
AND2x4_ASAP7_75t_L g437 ( .A(n_433), .B(n_438), .Y(n_437) );
NAND2x1p5_ASAP7_75t_L g443 ( .A(n_433), .B(n_444), .Y(n_443) );
AND2x4_ASAP7_75t_L g530 ( .A(n_433), .B(n_531), .Y(n_530) );
BUFx3_ASAP7_75t_L g608 ( .A(n_436), .Y(n_608) );
INVx2_ASAP7_75t_L g877 ( .A(n_436), .Y(n_877) );
BUFx2_ASAP7_75t_L g1040 ( .A(n_436), .Y(n_1040) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_437), .Y(n_525) );
BUFx12f_ASAP7_75t_L g578 ( .A(n_437), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B1(n_445), .B2(n_446), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_441), .A2(n_572), .B1(n_600), .B2(n_601), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_441), .A2(n_750), .B1(n_751), .B2(n_752), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g1126 ( .A1(n_441), .A2(n_572), .B1(n_1127), .B2(n_1128), .Y(n_1126) );
INVx3_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g570 ( .A(n_442), .Y(n_570) );
INVx4_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx3_ASAP7_75t_L g798 ( .A(n_443), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_443), .A2(n_447), .B1(n_909), .B2(n_910), .Y(n_908) );
HB1xp67_ASAP7_75t_L g956 ( .A(n_443), .Y(n_956) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_443), .A2(n_752), .B1(n_975), .B2(n_976), .Y(n_974) );
OAI22xp5_ASAP7_75t_L g1032 ( .A1(n_443), .A2(n_752), .B1(n_1033), .B2(n_1034), .Y(n_1032) );
AND2x2_ASAP7_75t_L g861 ( .A(n_444), .B(n_489), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_446), .A2(n_797), .B1(n_798), .B2(n_799), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_446), .A2(n_798), .B1(n_1004), .B2(n_1005), .Y(n_1003) );
BUFx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
CKINVDCx16_ASAP7_75t_R g573 ( .A(n_447), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g1079 ( .A1(n_447), .A2(n_469), .B1(n_1080), .B2(n_1081), .Y(n_1079) );
OR2x6_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_472), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_461), .Y(n_453) );
BUFx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_456), .Y(n_498) );
INVx3_ASAP7_75t_L g547 ( .A(n_456), .Y(n_547) );
BUFx3_ASAP7_75t_L g587 ( .A(n_456), .Y(n_587) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_SL g644 ( .A(n_457), .Y(n_644) );
INVx2_ASAP7_75t_L g667 ( .A(n_457), .Y(n_667) );
BUFx2_ASAP7_75t_SL g728 ( .A(n_457), .Y(n_728) );
AND2x2_ASAP7_75t_L g480 ( .A(n_458), .B(n_466), .Y(n_480) );
AND2x4_ASAP7_75t_L g488 ( .A(n_458), .B(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_458), .B(n_466), .Y(n_515) );
INVx11_ASAP7_75t_L g508 ( .A(n_459), .Y(n_508) );
INVx11_ASAP7_75t_L g589 ( .A(n_459), .Y(n_589) );
INVx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx4_ASAP7_75t_L g502 ( .A(n_464), .Y(n_502) );
INVx3_ASAP7_75t_L g705 ( .A(n_464), .Y(n_705) );
INVx1_ASAP7_75t_L g731 ( .A(n_464), .Y(n_731) );
INVx2_ASAP7_75t_L g784 ( .A(n_464), .Y(n_784) );
INVx5_ASAP7_75t_L g835 ( .A(n_464), .Y(n_835) );
INVx8_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx4f_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
BUFx2_ASAP7_75t_L g503 ( .A(n_468), .Y(n_503) );
BUFx2_ASAP7_75t_L g639 ( .A(n_468), .Y(n_639) );
BUFx2_ASAP7_75t_L g652 ( .A(n_468), .Y(n_652) );
BUFx2_ASAP7_75t_L g785 ( .A(n_468), .Y(n_785) );
INVx6_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g760 ( .A(n_469), .Y(n_760) );
INVx1_ASAP7_75t_SL g868 ( .A(n_469), .Y(n_868) );
INVx1_ASAP7_75t_SL g1168 ( .A(n_469), .Y(n_1168) );
OR2x6_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx1_ASAP7_75t_L g531 ( .A(n_470), .Y(n_531) );
INVx1_ASAP7_75t_L g489 ( .A(n_471), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_481), .Y(n_472) );
INVx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_475), .A2(n_511), .B1(n_512), .B2(n_513), .Y(n_510) );
INVx2_ASAP7_75t_L g596 ( .A(n_475), .Y(n_596) );
INVx2_ASAP7_75t_L g636 ( .A(n_475), .Y(n_636) );
INVx2_ASAP7_75t_L g650 ( .A(n_475), .Y(n_650) );
INVx6_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx3_ASAP7_75t_L g562 ( .A(n_476), .Y(n_562) );
BUFx3_ASAP7_75t_L g765 ( .A(n_476), .Y(n_765) );
BUFx3_ASAP7_75t_L g943 ( .A(n_476), .Y(n_943) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g1159 ( .A(n_479), .Y(n_1159) );
BUFx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx3_ASAP7_75t_L g642 ( .A(n_480), .Y(n_642) );
BUFx3_ASAP7_75t_L g726 ( .A(n_480), .Y(n_726) );
BUFx3_ASAP7_75t_L g782 ( .A(n_480), .Y(n_782) );
INVx4_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_483), .A2(n_505), .B1(n_506), .B2(n_509), .Y(n_504) );
INVx4_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx3_ASAP7_75t_L g592 ( .A(n_485), .Y(n_592) );
BUFx3_ASAP7_75t_L g638 ( .A(n_485), .Y(n_638) );
INVx2_ASAP7_75t_L g775 ( .A(n_485), .Y(n_775) );
BUFx3_ASAP7_75t_L g837 ( .A(n_485), .Y(n_837) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g890 ( .A(n_487), .Y(n_890) );
BUFx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_SL g499 ( .A(n_488), .Y(n_499) );
BUFx3_ASAP7_75t_L g548 ( .A(n_488), .Y(n_548) );
BUFx3_ASAP7_75t_L g593 ( .A(n_488), .Y(n_593) );
BUFx3_ASAP7_75t_L g668 ( .A(n_488), .Y(n_668) );
BUFx2_ASAP7_75t_L g702 ( .A(n_488), .Y(n_702) );
BUFx2_ASAP7_75t_SL g756 ( .A(n_488), .Y(n_756) );
INVx1_ASAP7_75t_L g1163 ( .A(n_488), .Y(n_1163) );
INVx1_ASAP7_75t_L g678 ( .A(n_492), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_542), .B1(n_675), .B2(n_676), .Y(n_492) );
INVx2_ASAP7_75t_L g676 ( .A(n_493), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_495), .B(n_516), .Y(n_494) );
NOR3xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_504), .C(n_510), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_500), .Y(n_496) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g759 ( .A(n_502), .Y(n_759) );
INVx1_ASAP7_75t_L g554 ( .A(n_503), .Y(n_554) );
INVx2_ASAP7_75t_L g772 ( .A(n_506), .Y(n_772) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
HB1xp67_ASAP7_75t_L g904 ( .A(n_507), .Y(n_904) );
INVx5_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_SL g558 ( .A(n_508), .Y(n_558) );
INVx1_ASAP7_75t_L g664 ( .A(n_508), .Y(n_664) );
INVx4_ASAP7_75t_L g856 ( .A(n_508), .Y(n_856) );
INVx2_ASAP7_75t_L g983 ( .A(n_508), .Y(n_983) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_513), .A2(n_560), .B1(n_561), .B2(n_563), .Y(n_559) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g900 ( .A(n_514), .Y(n_900) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_517), .B(n_526), .Y(n_516) );
OAI21xp5_ASAP7_75t_SL g517 ( .A1(n_518), .A2(n_519), .B(n_520), .Y(n_517) );
INVx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx4_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx2_ASAP7_75t_L g748 ( .A(n_523), .Y(n_748) );
INVx2_ASAP7_75t_L g793 ( .A(n_523), .Y(n_793) );
BUFx4f_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g815 ( .A(n_525), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_536), .Y(n_526) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx2_ASAP7_75t_L g633 ( .A(n_530), .Y(n_633) );
BUFx3_ASAP7_75t_L g661 ( .A(n_530), .Y(n_661) );
BUFx2_ASAP7_75t_L g1154 ( .A(n_530), .Y(n_1154) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx2_ASAP7_75t_SL g625 ( .A(n_535), .Y(n_625) );
BUFx2_ASAP7_75t_SL g670 ( .A(n_535), .Y(n_670) );
BUFx3_ASAP7_75t_L g1155 ( .A(n_535), .Y(n_1155) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g566 ( .A(n_538), .Y(n_566) );
INVx5_ASAP7_75t_L g631 ( .A(n_538), .Y(n_631) );
INVx2_ASAP7_75t_L g658 ( .A(n_538), .Y(n_658) );
INVx4_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
BUFx4f_ASAP7_75t_L g567 ( .A(n_541), .Y(n_567) );
BUFx2_ASAP7_75t_L g628 ( .A(n_541), .Y(n_628) );
INVx1_ASAP7_75t_SL g1058 ( .A(n_541), .Y(n_1058) );
INVx1_ASAP7_75t_L g675 ( .A(n_542), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_581), .B1(n_673), .B2(n_674), .Y(n_542) );
INVx1_ASAP7_75t_L g673 ( .A(n_543), .Y(n_673) );
INVx1_ASAP7_75t_L g580 ( .A(n_544), .Y(n_580) );
AND4x1_ASAP7_75t_L g544 ( .A(n_545), .B(n_555), .C(n_564), .D(n_574), .Y(n_544) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_551), .B1(n_553), .B2(n_554), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_551), .A2(n_892), .B1(n_893), .B2(n_894), .Y(n_891) );
OAI21xp33_ASAP7_75t_L g1165 ( .A1(n_551), .A2(n_1166), .B(n_1167), .Y(n_1165) );
BUFx2_ASAP7_75t_R g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g779 ( .A(n_561), .Y(n_779) );
INVx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B1(n_571), .B2(n_572), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g954 ( .A1(n_572), .A2(n_955), .B1(n_956), .B2(n_957), .Y(n_954) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g752 ( .A(n_573), .Y(n_752) );
INVx2_ASAP7_75t_L g713 ( .A(n_575), .Y(n_713) );
INVx4_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OAI21xp5_ASAP7_75t_SL g692 ( .A1(n_576), .A2(n_693), .B(n_694), .Y(n_692) );
BUFx2_ASAP7_75t_L g746 ( .A(n_576), .Y(n_746) );
BUFx4f_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g717 ( .A(n_578), .Y(n_717) );
INVx2_ASAP7_75t_L g674 ( .A(n_581), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_617), .B1(n_618), .B2(n_672), .Y(n_581) );
INVx1_ASAP7_75t_L g672 ( .A(n_582), .Y(n_672) );
INVx1_ASAP7_75t_SL g616 ( .A(n_583), .Y(n_616) );
AND2x2_ASAP7_75t_SL g583 ( .A(n_584), .B(n_598), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_585), .B(n_594), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_590), .Y(n_585) );
INVx4_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx3_ASAP7_75t_L g724 ( .A(n_589), .Y(n_724) );
INVx2_ASAP7_75t_SL g763 ( .A(n_589), .Y(n_763) );
INVx4_ASAP7_75t_L g919 ( .A(n_589), .Y(n_919) );
OAI21xp33_ASAP7_75t_SL g1076 ( .A1(n_589), .A2(n_1077), .B(n_1078), .Y(n_1076) );
NOR2xp33_ASAP7_75t_L g1169 ( .A(n_589), .B(n_1170), .Y(n_1169) );
BUFx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g906 ( .A(n_592), .Y(n_906) );
BUFx2_ASAP7_75t_L g776 ( .A(n_593), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
INVxp67_ASAP7_75t_L g898 ( .A(n_596), .Y(n_898) );
NOR3xp33_ASAP7_75t_SL g598 ( .A(n_599), .B(n_602), .C(n_609), .Y(n_598) );
OAI221xp5_ASAP7_75t_SL g950 ( .A1(n_604), .A2(n_713), .B1(n_951), .B2(n_952), .C(n_953), .Y(n_950) );
OAI221xp5_ASAP7_75t_SL g970 ( .A1(n_604), .A2(n_713), .B1(n_971), .B2(n_972), .C(n_973), .Y(n_970) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B1(n_613), .B2(n_614), .Y(n_609) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g968 ( .A(n_612), .Y(n_968) );
INVx2_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
XNOR2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_646), .Y(n_618) );
XOR2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_645), .Y(n_619) );
NAND3x1_ASAP7_75t_L g620 ( .A(n_621), .B(n_634), .C(n_640), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_626), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .C(n_632), .Y(n_626) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .Y(n_634) );
INVx2_ASAP7_75t_L g1025 ( .A(n_636), .Y(n_1025) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
BUFx3_ASAP7_75t_L g944 ( .A(n_642), .Y(n_944) );
XOR2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_671), .Y(n_646) );
NAND4xp75_ASAP7_75t_L g647 ( .A(n_648), .B(n_653), .C(n_662), .D(n_669), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
OA211x2_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .B(n_657), .C(n_659), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_655), .A2(n_788), .B1(n_789), .B2(n_790), .Y(n_787) );
INVx1_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g691 ( .A(n_656), .Y(n_691) );
INVx2_ASAP7_75t_L g1044 ( .A(n_656), .Y(n_1044) );
CKINVDCx20_ASAP7_75t_R g1123 ( .A(n_660), .Y(n_1123) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
INVx3_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx3_ASAP7_75t_L g831 ( .A(n_667), .Y(n_831) );
INVxp67_ASAP7_75t_L g1030 ( .A(n_668), .Y(n_1030) );
INVx1_ASAP7_75t_L g1098 ( .A(n_679), .Y(n_1098) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_961), .B1(n_1095), .B2(n_1096), .Y(n_679) );
INVx1_ASAP7_75t_L g1095 ( .A(n_680), .Y(n_1095) );
XOR2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_804), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_683), .B1(n_735), .B2(n_803), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OA22x2_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_685), .B1(n_708), .B2(n_734), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
XNOR2xp5_ASAP7_75t_L g737 ( .A(n_685), .B(n_738), .Y(n_737) );
XOR2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_707), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_698), .Y(n_686) );
NOR3xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_692), .C(n_695), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g966 ( .A1(n_691), .A2(n_967), .B1(n_968), .B2(n_969), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g994 ( .A1(n_691), .A2(n_968), .B1(n_995), .B2(n_996), .Y(n_994) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_703), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_706), .Y(n_703) );
INVx1_ASAP7_75t_L g734 ( .A(n_708), .Y(n_734) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_711), .B(n_721), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_712), .B(n_718), .Y(n_711) );
OAI21xp5_ASAP7_75t_SL g712 ( .A1(n_713), .A2(n_714), .B(n_715), .Y(n_712) );
OAI221xp5_ASAP7_75t_L g791 ( .A1(n_713), .A2(n_792), .B1(n_793), .B2(n_794), .C(n_795), .Y(n_791) );
OAI221xp5_ASAP7_75t_L g1035 ( .A1(n_713), .A2(n_1036), .B1(n_1037), .B2(n_1038), .C(n_1039), .Y(n_1035) );
OAI221xp5_ASAP7_75t_SL g1121 ( .A1(n_713), .A2(n_1122), .B1(n_1123), .B2(n_1124), .C(n_1125), .Y(n_1121) );
INVx3_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_729), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_727), .Y(n_722) );
BUFx4f_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .Y(n_729) );
HB1xp67_ASAP7_75t_L g1022 ( .A(n_731), .Y(n_1022) );
INVx1_ASAP7_75t_L g803 ( .A(n_735), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .B1(n_767), .B2(n_802), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
XOR2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_766), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_753), .Y(n_739) );
NOR3xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_744), .C(n_749), .Y(n_740) );
OAI21xp33_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B(n_747), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_761), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_757), .Y(n_754) );
INVx3_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_764), .Y(n_761) );
INVx1_ASAP7_75t_L g802 ( .A(n_767), .Y(n_802) );
INVx2_ASAP7_75t_L g801 ( .A(n_768), .Y(n_801) );
AND2x2_ASAP7_75t_SL g768 ( .A(n_769), .B(n_786), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g769 ( .A(n_770), .B(n_777), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_773), .Y(n_770) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_778), .B(n_783), .Y(n_777) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVxp67_ASAP7_75t_L g894 ( .A(n_785), .Y(n_894) );
NOR3xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_791), .C(n_796), .Y(n_786) );
INVx1_ASAP7_75t_L g821 ( .A(n_789), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_789), .A2(n_1042), .B1(n_1043), .B2(n_1044), .Y(n_1041) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_798), .A2(n_824), .B1(n_825), .B2(n_826), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_806), .B1(n_879), .B2(n_880), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_808), .B1(n_839), .B2(n_840), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
XOR2x2_ASAP7_75t_L g808 ( .A(n_809), .B(n_838), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_827), .Y(n_809) );
NOR3xp33_ASAP7_75t_L g810 ( .A(n_811), .B(n_818), .C(n_823), .Y(n_810) );
OAI221xp5_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_814), .B1(n_815), .B2(n_816), .C(n_817), .Y(n_811) );
OAI21xp5_ASAP7_75t_L g845 ( .A1(n_812), .A2(n_846), .B(n_847), .Y(n_845) );
OAI21xp5_ASAP7_75t_SL g1149 ( .A1(n_812), .A2(n_1150), .B(n_1151), .Y(n_1149) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx2_ASAP7_75t_SL g998 ( .A(n_813), .Y(n_998) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_828), .B(n_832), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
INVxp67_ASAP7_75t_L g888 ( .A(n_831), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_836), .Y(n_832) );
BUFx6f_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
BUFx2_ASAP7_75t_L g1161 ( .A(n_837), .Y(n_1161) );
INVx1_ASAP7_75t_SL g839 ( .A(n_840), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_842), .B1(n_863), .B2(n_878), .Y(n_840) );
INVx3_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
XOR2x2_ASAP7_75t_L g842 ( .A(n_843), .B(n_862), .Y(n_842) );
NAND2xp5_ASAP7_75t_SL g843 ( .A(n_844), .B(n_853), .Y(n_843) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_845), .B(n_848), .Y(n_844) );
NAND3xp33_ASAP7_75t_L g848 ( .A(n_849), .B(n_850), .C(n_851), .Y(n_848) );
INVx1_ASAP7_75t_L g1000 ( .A(n_852), .Y(n_1000) );
NOR2x1_ASAP7_75t_L g853 ( .A(n_854), .B(n_858), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_855), .B(n_857), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_860), .Y(n_858) );
INVx1_ASAP7_75t_L g878 ( .A(n_863), .Y(n_878) );
NAND4xp75_ASAP7_75t_L g864 ( .A(n_865), .B(n_869), .C(n_872), .D(n_875), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
AND2x2_ASAP7_75t_SL g869 ( .A(n_870), .B(n_871), .Y(n_869) );
AND2x2_ASAP7_75t_L g872 ( .A(n_873), .B(n_874), .Y(n_872) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
OAI22xp5_ASAP7_75t_SL g880 ( .A1(n_881), .A2(n_882), .B1(n_935), .B2(n_960), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g882 ( .A1(n_883), .A2(n_914), .B1(n_933), .B2(n_934), .Y(n_882) );
INVx1_ASAP7_75t_L g933 ( .A(n_883), .Y(n_933) );
INVx1_ASAP7_75t_L g913 ( .A(n_884), .Y(n_913) );
AND4x1_ASAP7_75t_L g884 ( .A(n_885), .B(n_895), .C(n_907), .D(n_911), .Y(n_884) );
NOR2xp33_ASAP7_75t_SL g885 ( .A(n_886), .B(n_891), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_887), .A2(n_888), .B1(n_889), .B2(n_890), .Y(n_886) );
INVx2_ASAP7_75t_L g1136 ( .A(n_890), .Y(n_1136) );
NOR2xp33_ASAP7_75t_L g895 ( .A(n_896), .B(n_901), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_897), .A2(n_898), .B1(n_899), .B2(n_900), .Y(n_896) );
OAI22xp5_ASAP7_75t_L g1023 ( .A1(n_900), .A2(n_1024), .B1(n_1025), .B2(n_1026), .Y(n_1023) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_902), .A2(n_903), .B1(n_905), .B2(n_906), .Y(n_901) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g1027 ( .A1(n_906), .A2(n_1028), .B1(n_1029), .B2(n_1030), .Y(n_1027) );
INVx2_ASAP7_75t_SL g934 ( .A(n_914), .Y(n_934) );
OAI22xp5_ASAP7_75t_L g989 ( .A1(n_914), .A2(n_934), .B1(n_990), .B2(n_991), .Y(n_989) );
XNOR2x2_ASAP7_75t_L g914 ( .A(n_915), .B(n_916), .Y(n_914) );
NOR4xp75_ASAP7_75t_L g916 ( .A(n_917), .B(n_921), .C(n_924), .D(n_928), .Y(n_916) );
NAND2xp5_ASAP7_75t_SL g917 ( .A(n_918), .B(n_920), .Y(n_917) );
NAND2xp5_ASAP7_75t_SL g921 ( .A(n_922), .B(n_923), .Y(n_921) );
OAI21xp5_ASAP7_75t_SL g928 ( .A1(n_929), .A2(n_931), .B(n_932), .Y(n_928) );
OAI21xp5_ASAP7_75t_SL g1052 ( .A1(n_929), .A2(n_1053), .B(n_1054), .Y(n_1052) );
INVx3_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g960 ( .A(n_935), .Y(n_960) );
INVx1_ASAP7_75t_L g959 ( .A(n_936), .Y(n_959) );
AND2x2_ASAP7_75t_SL g936 ( .A(n_937), .B(n_946), .Y(n_936) );
NOR2xp33_ASAP7_75t_L g937 ( .A(n_938), .B(n_941), .Y(n_937) );
NAND2xp33_ASAP7_75t_SL g938 ( .A(n_939), .B(n_940), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_942), .B(n_945), .Y(n_941) );
NOR3xp33_ASAP7_75t_L g946 ( .A(n_947), .B(n_950), .C(n_954), .Y(n_946) );
INVx2_ASAP7_75t_L g1096 ( .A(n_961), .Y(n_1096) );
AOI22xp5_ASAP7_75t_L g961 ( .A1(n_962), .A2(n_987), .B1(n_1093), .B2(n_1094), .Y(n_961) );
INVxp67_ASAP7_75t_L g1093 ( .A(n_962), .Y(n_1093) );
HB1xp67_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx1_ASAP7_75t_SL g985 ( .A(n_964), .Y(n_985) );
AND2x2_ASAP7_75t_SL g964 ( .A(n_965), .B(n_977), .Y(n_964) );
NOR3xp33_ASAP7_75t_L g965 ( .A(n_966), .B(n_970), .C(n_974), .Y(n_965) );
NOR2xp33_ASAP7_75t_L g977 ( .A(n_978), .B(n_981), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_979), .B(n_980), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_982), .B(n_984), .Y(n_981) );
INVx1_ASAP7_75t_L g1094 ( .A(n_987), .Y(n_1094) );
AOI22xp5_ASAP7_75t_L g987 ( .A1(n_988), .A2(n_989), .B1(n_1015), .B2(n_1092), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx2_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx2_ASAP7_75t_SL g1014 ( .A(n_992), .Y(n_1014) );
AND2x2_ASAP7_75t_L g992 ( .A(n_993), .B(n_1006), .Y(n_992) );
NOR3xp33_ASAP7_75t_L g993 ( .A(n_994), .B(n_997), .C(n_1003), .Y(n_993) );
OAI221xp5_ASAP7_75t_SL g997 ( .A1(n_998), .A2(n_999), .B1(n_1000), .B2(n_1001), .C(n_1002), .Y(n_997) );
NOR2xp33_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1010), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1009), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1012), .Y(n_1010) );
INVx2_ASAP7_75t_SL g1092 ( .A(n_1015), .Y(n_1092) );
OA22x2_ASAP7_75t_L g1015 ( .A1(n_1016), .A2(n_1047), .B1(n_1090), .B2(n_1091), .Y(n_1015) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1016), .Y(n_1090) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1017), .Y(n_1046) );
AND2x2_ASAP7_75t_SL g1017 ( .A(n_1018), .B(n_1031), .Y(n_1017) );
NOR3xp33_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1023), .C(n_1027), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1021), .Y(n_1019) );
NOR3xp33_ASAP7_75t_SL g1031 ( .A(n_1032), .B(n_1035), .C(n_1041), .Y(n_1031) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1047), .Y(n_1091) );
XOR2x2_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1069), .Y(n_1047) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1050), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1061), .Y(n_1050) );
NOR2xp67_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1055), .Y(n_1051) );
NAND3xp33_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1059), .C(n_1060), .Y(n_1055) );
INVx1_ASAP7_75t_SL g1057 ( .A(n_1058), .Y(n_1057) );
NOR2x1_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1065), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1064), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1067), .Y(n_1065) );
INVx2_ASAP7_75t_L g1089 ( .A(n_1071), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1082), .Y(n_1071) );
NOR3xp33_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1076), .C(n_1079), .Y(n_1072) );
NOR2xp33_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1086), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1085), .Y(n_1083) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_1087), .B(n_1088), .Y(n_1086) );
INVx1_ASAP7_75t_SL g1099 ( .A(n_1100), .Y(n_1099) );
NOR2x1_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1105), .Y(n_1100) );
OR2x2_ASAP7_75t_SL g1173 ( .A(n_1101), .B(n_1106), .Y(n_1173) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1104), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g1138 ( .A(n_1103), .Y(n_1138) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_1103), .B(n_1141), .Y(n_1144) );
CKINVDCx16_ASAP7_75t_R g1141 ( .A(n_1104), .Y(n_1141) );
CKINVDCx20_ASAP7_75t_R g1105 ( .A(n_1106), .Y(n_1105) );
NAND2xp5_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1108), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1111), .Y(n_1109) );
OAI322xp33_ASAP7_75t_L g1112 ( .A1(n_1113), .A2(n_1138), .A3(n_1139), .B1(n_1142), .B2(n_1145), .C1(n_1146), .C2(n_1171), .Y(n_1112) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx2_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1117), .B(n_1129), .Y(n_1116) );
NOR3xp33_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1121), .C(n_1126), .Y(n_1117) );
NOR2xp33_ASAP7_75t_L g1129 ( .A(n_1130), .B(n_1133), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1132), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1135), .Y(n_1133) );
HB1xp67_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
CKINVDCx20_ASAP7_75t_R g1142 ( .A(n_1143), .Y(n_1142) );
NAND3x1_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1157), .C(n_1164), .Y(n_1147) );
NOR2xp33_ASAP7_75t_L g1148 ( .A(n_1149), .B(n_1152), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_1153), .B(n_1156), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1160), .Y(n_1157) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
CKINVDCx20_ASAP7_75t_R g1171 ( .A(n_1172), .Y(n_1171) );
CKINVDCx20_ASAP7_75t_R g1172 ( .A(n_1173), .Y(n_1172) );
endmodule