module fake_netlist_1_1212_n_18 (n_1, n_2, n_0, n_18);
input n_1;
input n_2;
input n_0;
output n_18;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_17;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
NAND2xp5_ASAP7_75t_SL g3 ( .A(n_1), .B(n_2), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_1), .Y(n_5) );
NOR2xp33_ASAP7_75t_SL g6 ( .A(n_4), .B(n_0), .Y(n_6) );
INVx2_ASAP7_75t_SL g7 ( .A(n_5), .Y(n_7) );
NAND2xp33_ASAP7_75t_R g8 ( .A(n_3), .B(n_2), .Y(n_8) );
AND2x2_ASAP7_75t_L g9 ( .A(n_7), .B(n_6), .Y(n_9) );
AND2x2_ASAP7_75t_L g10 ( .A(n_7), .B(n_3), .Y(n_10) );
INVxp67_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
NAND2xp5_ASAP7_75t_SL g12 ( .A(n_9), .B(n_6), .Y(n_12) );
OAI21xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_10), .B(n_7), .Y(n_13) );
OAI31xp33_ASAP7_75t_SL g14 ( .A1(n_11), .A2(n_8), .A3(n_1), .B(n_2), .Y(n_14) );
NAND4xp75_ASAP7_75t_L g15 ( .A(n_13), .B(n_0), .C(n_1), .D(n_2), .Y(n_15) );
OR2x2_ASAP7_75t_L g16 ( .A(n_14), .B(n_0), .Y(n_16) );
NAND2x1_ASAP7_75t_SL g17 ( .A(n_15), .B(n_14), .Y(n_17) );
OAI21xp5_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_16), .B(n_12), .Y(n_18) );
endmodule