module fake_jpeg_27763_n_291 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_291);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_291;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVxp33_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_23),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_54),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_51),
.B(n_57),
.Y(n_97)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_20),
.B1(n_33),
.B2(n_30),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_64),
.B1(n_70),
.B2(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_59),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_26),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_62),
.B(n_67),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_30),
.B1(n_27),
.B2(n_26),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_48),
.A2(n_38),
.B1(n_29),
.B2(n_21),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_65),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_66),
.A2(n_28),
.B(n_32),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_22),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_35),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_47),
.A2(n_22),
.B1(n_27),
.B2(n_21),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_38),
.B1(n_29),
.B2(n_28),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_43),
.A2(n_28),
.B1(n_35),
.B2(n_34),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_28),
.B1(n_18),
.B2(n_34),
.Y(n_110)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_36),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_23),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_81),
.A2(n_36),
.B1(n_25),
.B2(n_18),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_83),
.A2(n_110),
.B1(n_113),
.B2(n_1),
.Y(n_138)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_99),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_80),
.A2(n_79),
.B1(n_60),
.B2(n_58),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_89),
.B(n_32),
.Y(n_133)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_23),
.C(n_25),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_91),
.B(n_2),
.C(n_4),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_23),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_93),
.A2(n_106),
.B(n_0),
.Y(n_137)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_105),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_60),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_31),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_104),
.B(n_109),
.Y(n_126)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_31),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_34),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_61),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_16),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_116),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_78),
.A2(n_18),
.B1(n_32),
.B2(n_2),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

BUFx8_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_68),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_118),
.A2(n_73),
.B1(n_71),
.B2(n_63),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_131),
.B1(n_83),
.B2(n_93),
.Y(n_150)
);

NOR2x1_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_66),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_135),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_54),
.B(n_50),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_123),
.A2(n_134),
.B(n_141),
.Y(n_172)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_129),
.B(n_132),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_130),
.B(n_133),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_73),
.B1(n_71),
.B2(n_63),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_61),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_132),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_146),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_117),
.B1(n_97),
.B2(n_91),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_82),
.A2(n_93),
.B(n_111),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_106),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

BUFx16f_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_167),
.B1(n_174),
.B2(n_140),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_150),
.A2(n_168),
.B1(n_157),
.B2(n_152),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_114),
.C(n_87),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_151),
.B(n_166),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_153),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_105),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_122),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_157),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_94),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_159),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_123),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_126),
.B(n_4),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_169),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_87),
.C(n_94),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_138),
.A2(n_90),
.B1(n_88),
.B2(n_108),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_120),
.A2(n_88),
.B1(n_98),
.B2(n_107),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_134),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_170),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_107),
.Y(n_171)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_173),
.A2(n_176),
.B(n_147),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_140),
.A2(n_92),
.B1(n_84),
.B2(n_115),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_122),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_92),
.Y(n_177)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_84),
.Y(n_178)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

XNOR2x1_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_137),
.Y(n_180)
);

FAx1_ASAP7_75t_SL g208 ( 
.A(n_180),
.B(n_175),
.CI(n_150),
.CON(n_208),
.SN(n_208)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_181),
.A2(n_183),
.B(n_198),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_193),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_166),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_130),
.B1(n_125),
.B2(n_144),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_187),
.A2(n_190),
.B1(n_196),
.B2(n_197),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_125),
.B1(n_128),
.B2(n_121),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_172),
.A2(n_147),
.B(n_146),
.Y(n_193)
);

AO22x1_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_124),
.B1(n_128),
.B2(n_121),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_190),
.Y(n_216)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_201),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_124),
.B1(n_5),
.B2(n_6),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_149),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_7),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_158),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_199)
);

OAI22x1_ASAP7_75t_L g206 ( 
.A1(n_199),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_170),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_200)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_206),
.Y(n_243)
);

AOI221xp5_ASAP7_75t_L g207 ( 
.A1(n_203),
.A2(n_156),
.B1(n_161),
.B2(n_164),
.C(n_175),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_193),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_208),
.A2(n_216),
.B(n_219),
.Y(n_227)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_202),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_210),
.Y(n_229)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

OAI22x1_ASAP7_75t_L g212 ( 
.A1(n_180),
.A2(n_174),
.B1(n_161),
.B2(n_155),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_212),
.A2(n_225),
.B(n_226),
.Y(n_242)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_217),
.Y(n_233)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_185),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_222),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_163),
.Y(n_224)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_176),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_204),
.C(n_183),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_236),
.C(n_238),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_232),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_183),
.B1(n_184),
.B2(n_198),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_234),
.A2(n_239),
.B1(n_220),
.B2(n_154),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_204),
.C(n_189),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_224),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_182),
.C(n_179),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_225),
.A2(n_196),
.B1(n_197),
.B2(n_200),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_226),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_240),
.Y(n_252)
);

A2O1A1O1Ixp25_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_212),
.B(n_208),
.C(n_218),
.D(n_214),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_238),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_226),
.B(n_223),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_250),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_248),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_247),
.B(n_228),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_230),
.A2(n_214),
.B(n_198),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_229),
.A2(n_213),
.B(n_206),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_254),
.Y(n_262)
);

NOR3xp33_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_213),
.C(n_208),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_215),
.B(n_220),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_242),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_229),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_233),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_227),
.A2(n_165),
.B(n_173),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_237),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_258),
.A2(n_263),
.B(n_266),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_260),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_243),
.B1(n_241),
.B2(n_231),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_267),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_265),
.B(n_233),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_241),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_261),
.B(n_247),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_271),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_253),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_234),
.B(n_236),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_251),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_274),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_274),
.A2(n_239),
.B1(n_259),
.B2(n_244),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_275),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_253),
.C(n_260),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_278),
.C(n_269),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_245),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_279),
.A2(n_14),
.B(n_15),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_280),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_246),
.C(n_160),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_279),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_284),
.Y(n_285)
);

AOI322xp5_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_14),
.A3(n_15),
.B1(n_148),
.B2(n_160),
.C1(n_281),
.C2(n_285),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_288),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_286),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_290),
.Y(n_291)
);


endmodule