module fake_netlist_5_2079_n_162 (n_29, n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_162);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_162;

wire n_137;
wire n_91;
wire n_82;
wire n_122;
wire n_142;
wire n_140;
wire n_136;
wire n_86;
wire n_146;
wire n_124;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_111;
wire n_108;
wire n_129;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_69;
wire n_58;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_125;
wire n_35;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_30;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_79;
wire n_131;
wire n_151;
wire n_47;
wire n_53;
wire n_160;
wire n_158;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_154;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_95;
wire n_119;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_150;
wire n_64;
wire n_77;
wire n_106;
wire n_102;
wire n_161;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_134;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_141;
wire n_63;
wire n_51;
wire n_97;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

INVxp67_ASAP7_75t_SL g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

AND2x6_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_15),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_0),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

AND3x1_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_0),
.C(n_2),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_35),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_52),
.B1(n_50),
.B2(n_37),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_72),
.Y(n_76)
);

AND2x4_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_69),
.Y(n_77)
);

NAND2x1p5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_41),
.Y(n_78)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_52),
.B1(n_50),
.B2(n_30),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_41),
.Y(n_81)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_31),
.C(n_38),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

AND2x4_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_31),
.B1(n_38),
.B2(n_44),
.Y(n_88)
);

AO22x2_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_45),
.B1(n_42),
.B2(n_8),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_32),
.B1(n_40),
.B2(n_58),
.Y(n_92)
);

AOI22x1_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_56),
.B1(n_57),
.B2(n_73),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_81),
.B(n_76),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_67),
.B(n_66),
.C(n_64),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_64),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_56),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_88),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_74),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_92),
.Y(n_109)
);

OR2x6_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

NOR2x1_ASAP7_75t_SL g112 ( 
.A(n_108),
.B(n_95),
.Y(n_112)
);

AOI221xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_79),
.B1(n_82),
.B2(n_89),
.C(n_78),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_96),
.B(n_82),
.C(n_86),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_105),
.B(n_107),
.Y(n_116)
);

OAI21x1_ASAP7_75t_L g117 ( 
.A1(n_113),
.A2(n_93),
.B(n_106),
.Y(n_117)
);

AO21x2_ASAP7_75t_L g118 ( 
.A1(n_114),
.A2(n_106),
.B(n_102),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_115),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_103),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_102),
.B(n_93),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_110),
.Y(n_125)
);

AO21x2_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_112),
.B(n_90),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_117),
.Y(n_128)
);

INVxp67_ASAP7_75t_SL g129 ( 
.A(n_119),
.Y(n_129)
);

NAND2x1_ASAP7_75t_SL g130 ( 
.A(n_127),
.B(n_123),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g136 ( 
.A(n_131),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_134),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_130),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_120),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_130),
.Y(n_143)
);

AND2x4_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_126),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

AOI221xp5_ASAP7_75t_L g149 ( 
.A1(n_147),
.A2(n_51),
.B1(n_62),
.B2(n_137),
.C(n_3),
.Y(n_149)
);

OR3x2_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_5),
.C(n_9),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_121),
.B(n_119),
.Y(n_152)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_146),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

NAND5xp2_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_121),
.C(n_9),
.D(n_144),
.E(n_16),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_152),
.Y(n_156)
);

NAND4xp25_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_150),
.C(n_51),
.D(n_22),
.Y(n_157)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_153),
.A2(n_11),
.A3(n_12),
.B1(n_24),
.B2(n_25),
.C1(n_27),
.C2(n_28),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_156),
.A2(n_58),
.B1(n_97),
.B2(n_124),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_154),
.Y(n_160)
);

OAI322xp33_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_158),
.A3(n_159),
.B1(n_58),
.B2(n_97),
.C1(n_95),
.C2(n_124),
.Y(n_161)
);

AOI221xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_95),
.B1(n_97),
.B2(n_160),
.C(n_150),
.Y(n_162)
);


endmodule