module fake_jpeg_19058_n_345 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_29),
.Y(n_58)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_20),
.B1(n_44),
.B2(n_42),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_50),
.A2(n_31),
.B1(n_30),
.B2(n_23),
.Y(n_88)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_37),
.B(n_34),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_64),
.B(n_26),
.Y(n_78)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_38),
.A2(n_20),
.B1(n_25),
.B2(n_22),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_23),
.B1(n_31),
.B2(n_30),
.Y(n_83)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_41),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_79),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_20),
.B1(n_25),
.B2(n_22),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_72),
.A2(n_55),
.B1(n_23),
.B2(n_47),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_50),
.B(n_58),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_93),
.B(n_48),
.Y(n_103)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_25),
.B1(n_28),
.B2(n_22),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_75),
.A2(n_83),
.B1(n_89),
.B2(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_78),
.B(n_27),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_46),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_85),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_18),
.C(n_46),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_94),
.Y(n_110)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_61),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_86),
.Y(n_116)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_97),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_43),
.B1(n_41),
.B2(n_38),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_25),
.B1(n_28),
.B2(n_26),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

BUFx24_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_28),
.B(n_21),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_14),
.B(n_16),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_51),
.A2(n_53),
.B(n_56),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_62),
.B(n_48),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_21),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_98),
.B(n_43),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_32),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_101),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_117),
.B(n_110),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_106),
.B(n_129),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_109),
.B(n_119),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_47),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_79),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_120),
.A2(n_14),
.B(n_16),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_131),
.B1(n_132),
.B2(n_85),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_84),
.B(n_13),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_122),
.B(n_129),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_36),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_128),
.Y(n_151)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_91),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_18),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_98),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_84),
.A2(n_24),
.B1(n_33),
.B2(n_19),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_93),
.B(n_33),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_82),
.C(n_94),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_113),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_156),
.B1(n_115),
.B2(n_130),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_128),
.B(n_94),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_137),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_18),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_139),
.A2(n_144),
.B1(n_113),
.B2(n_102),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_132),
.A2(n_90),
.B(n_74),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_142),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_91),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_113),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_70),
.B1(n_69),
.B2(n_68),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_146),
.A2(n_149),
.B1(n_154),
.B2(n_126),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_101),
.B(n_87),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_103),
.A2(n_119),
.B1(n_105),
.B2(n_117),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_161),
.B1(n_133),
.B2(n_116),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_80),
.B1(n_76),
.B2(n_24),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_150),
.B(n_152),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_160),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_105),
.A2(n_123),
.B1(n_107),
.B2(n_106),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_155),
.A2(n_122),
.B(n_109),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_102),
.A2(n_76),
.B1(n_100),
.B2(n_77),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_18),
.C(n_35),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_133),
.C(n_35),
.Y(n_162)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_127),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_107),
.B(n_18),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_108),
.A2(n_24),
.B1(n_33),
.B2(n_19),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_163),
.A2(n_183),
.B1(n_140),
.B2(n_161),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_L g217 ( 
.A1(n_164),
.A2(n_182),
.B(n_166),
.Y(n_217)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_188),
.Y(n_193)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_172),
.Y(n_196)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_174),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_180),
.B1(n_152),
.B2(n_178),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_35),
.C(n_24),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_116),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_190),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_115),
.B1(n_118),
.B2(n_126),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

AND2x6_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_113),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_143),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_191),
.Y(n_197)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_126),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_150),
.B(n_125),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_124),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_112),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_151),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_220),
.C(n_223),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_136),
.B1(n_140),
.B2(n_137),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_198),
.A2(n_200),
.B1(n_206),
.B2(n_217),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_199),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_137),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_213),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_137),
.B1(n_139),
.B2(n_134),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_203),
.A2(n_216),
.B1(n_175),
.B2(n_173),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_176),
.A2(n_139),
.B1(n_157),
.B2(n_159),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_168),
.A2(n_124),
.B(n_158),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_209),
.A2(n_0),
.B(n_1),
.Y(n_249)
);

INVxp67_ASAP7_75t_SL g211 ( 
.A(n_182),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_211),
.B(n_222),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_171),
.Y(n_212)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_19),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_19),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_218),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_168),
.A2(n_158),
.B1(n_112),
.B2(n_124),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_175),
.B(n_33),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_180),
.Y(n_221)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g222 ( 
.A(n_188),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_173),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_238),
.B(n_239),
.Y(n_253)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_207),
.Y(n_260)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_192),
.C(n_162),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_230),
.B(n_242),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_240),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_200),
.A2(n_172),
.B1(n_167),
.B2(n_112),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_219),
.A2(n_29),
.B1(n_32),
.B2(n_35),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_235),
.A2(n_250),
.B1(n_249),
.B2(n_214),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_35),
.B(n_9),
.Y(n_238)
);

AND2x4_ASAP7_75t_SL g239 ( 
.A(n_209),
.B(n_210),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_221),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_208),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_241),
.B(n_204),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_193),
.B(n_15),
.C(n_13),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_208),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_244),
.B(n_245),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_193),
.B(n_15),
.C(n_12),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_201),
.Y(n_246)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_246),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_215),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_250)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_228),
.Y(n_256)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_201),
.Y(n_258)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_258),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_266),
.Y(n_278)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_260),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_205),
.Y(n_262)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_224),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_264),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_267),
.Y(n_272)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_246),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_248),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_269),
.A2(n_218),
.B(n_194),
.Y(n_287)
);

AOI21xp33_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_202),
.B(n_234),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_259),
.A2(n_236),
.B1(n_247),
.B2(n_232),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_273),
.A2(n_269),
.B1(n_266),
.B2(n_258),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_225),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_283),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_271),
.A2(n_203),
.B1(n_239),
.B2(n_207),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_276),
.A2(n_285),
.B1(n_257),
.B2(n_240),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_225),
.C(n_230),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_220),
.C(n_255),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_226),
.B(n_231),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_252),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_223),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_284),
.A2(n_289),
.B(n_268),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_271),
.A2(n_235),
.B1(n_210),
.B2(n_226),
.Y(n_285)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_287),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_261),
.A2(n_194),
.B(n_245),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_292),
.B(n_296),
.Y(n_310)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_294),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_256),
.C(n_251),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_292),
.C(n_301),
.Y(n_318)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_251),
.C(n_255),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_287),
.C(n_277),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_298),
.A2(n_302),
.B1(n_305),
.B2(n_278),
.Y(n_311)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_303),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_301),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_283),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_252),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_273),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_276),
.A2(n_278),
.B1(n_285),
.B2(n_275),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_250),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_306),
.A2(n_282),
.B1(n_233),
.B2(n_9),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_314),
.Y(n_323)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_311),
.Y(n_319)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_297),
.A2(n_279),
.B1(n_242),
.B2(n_286),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_229),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_315),
.B(n_318),
.Y(n_321)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_316),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_291),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_317),
.A2(n_10),
.B(n_3),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_309),
.A2(n_305),
.B1(n_295),
.B2(n_303),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_320),
.A2(n_327),
.B1(n_308),
.B2(n_312),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_325),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_307),
.A2(n_293),
.B(n_3),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_310),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_326),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_328),
.B(n_329),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_318),
.C(n_315),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_332),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_312),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_313),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_333),
.A2(n_334),
.B(n_314),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_323),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_336),
.B(n_328),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_335),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_337),
.B(n_330),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_340),
.A2(n_4),
.B(n_5),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_4),
.B(n_5),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_7),
.C(n_5),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_6),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_6),
.B(n_270),
.Y(n_345)
);


endmodule