module fake_jpeg_19637_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_33),
.Y(n_63)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_43),
.Y(n_74)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_57),
.Y(n_95)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_20),
.Y(n_57)
);

NAND2x1_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_32),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_63),
.Y(n_78)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_40),
.B(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_68),
.Y(n_106)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_23),
.B1(n_44),
.B2(n_17),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_72),
.A2(n_43),
.B1(n_34),
.B2(n_19),
.Y(n_105)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

BUFx4f_ASAP7_75t_SL g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_85),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_51),
.B(n_64),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_48),
.Y(n_116)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_83),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_17),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_86),
.B(n_93),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_45),
.B1(n_44),
.B2(n_23),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_87),
.A2(n_96),
.B1(n_101),
.B2(n_47),
.Y(n_129)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_92),
.Y(n_127)
);

AO22x1_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_43),
.B1(n_44),
.B2(n_50),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_89),
.A2(n_96),
.B1(n_111),
.B2(n_101),
.Y(n_121)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_30),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_61),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_94),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_58),
.A2(n_19),
.B1(n_42),
.B2(n_41),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_98),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_31),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_68),
.A2(n_19),
.B1(n_42),
.B2(n_41),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

FAx1_ASAP7_75t_SL g104 ( 
.A(n_73),
.B(n_42),
.CI(n_32),
.CON(n_104),
.SN(n_104)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_104),
.A2(n_76),
.A3(n_89),
.B1(n_114),
.B2(n_95),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_107),
.B1(n_109),
.B2(n_111),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_56),
.A2(n_43),
.B1(n_48),
.B2(n_46),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_62),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_108),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_65),
.A2(n_43),
.B1(n_34),
.B2(n_25),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_67),
.A2(n_70),
.B(n_74),
.C(n_25),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_115),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_116),
.A2(n_134),
.B(n_144),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_121),
.A2(n_129),
.B1(n_150),
.B2(n_1),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_46),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_136),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_78),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_133),
.A2(n_115),
.B1(n_113),
.B2(n_100),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_82),
.A2(n_106),
.B(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_28),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_146),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_112),
.A2(n_37),
.B1(n_26),
.B2(n_31),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_102),
.A2(n_28),
.B(n_27),
.C(n_37),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_91),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_84),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_92),
.B(n_36),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_97),
.A2(n_26),
.B1(n_36),
.B2(n_29),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_153),
.B(n_172),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_155),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_80),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_165),
.C(n_166),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_137),
.A2(n_79),
.B1(n_77),
.B2(n_94),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_18),
.B1(n_29),
.B2(n_36),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_118),
.A2(n_29),
.B1(n_36),
.B2(n_18),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_118),
.A2(n_29),
.B1(n_33),
.B2(n_32),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_161),
.A2(n_171),
.B1(n_177),
.B2(n_185),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_168),
.B1(n_173),
.B2(n_176),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_33),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_84),
.C(n_33),
.Y(n_166)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_121),
.A2(n_136),
.B1(n_142),
.B2(n_116),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_167),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_116),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_33),
.B1(n_32),
.B2(n_24),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_32),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_146),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_24),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_174),
.B(n_178),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_124),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_120),
.A2(n_7),
.B1(n_11),
.B2(n_8),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_130),
.B(n_24),
.Y(n_178)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_184),
.Y(n_190)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

FAx1_ASAP7_75t_SL g183 ( 
.A(n_133),
.B(n_21),
.CI(n_16),
.CON(n_183),
.SN(n_183)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_131),
.Y(n_187)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_144),
.A2(n_21),
.B1(n_16),
.B2(n_3),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_131),
.B(n_138),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_186),
.A2(n_187),
.B(n_201),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_169),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_189),
.B(n_193),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_179),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_170),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_194),
.B(n_208),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_122),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_196),
.Y(n_227)
);

AO221x1_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_147),
.B1(n_125),
.B2(n_117),
.C(n_122),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_126),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_206),
.Y(n_233)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

AND2x4_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_163),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_160),
.A2(n_149),
.B(n_119),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_203),
.A2(n_205),
.B(n_1),
.Y(n_234)
);

NAND2x1_ASAP7_75t_L g205 ( 
.A(n_152),
.B(n_125),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_139),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_167),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_117),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_209),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_156),
.B(n_119),
.C(n_128),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_165),
.C(n_183),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_132),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_217),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_176),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_213),
.Y(n_231)
);

MAJx2_ASAP7_75t_L g215 ( 
.A(n_167),
.B(n_21),
.C(n_16),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_183),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_166),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_192),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_219),
.B(n_223),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_216),
.A2(n_164),
.B1(n_162),
.B2(n_159),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_221),
.A2(n_229),
.B1(n_230),
.B2(n_232),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_238),
.C(n_204),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_192),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_222),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_216),
.A2(n_162),
.B1(n_161),
.B2(n_173),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_214),
.A2(n_185),
.B1(n_168),
.B2(n_132),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_214),
.A2(n_128),
.B1(n_147),
.B2(n_177),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_234),
.A2(n_187),
.B(n_206),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_190),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_237),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_202),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_6),
.C(n_8),
.Y(n_238)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_2),
.Y(n_241)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_241),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_186),
.B(n_204),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_211),
.Y(n_262)
);

OAI22x1_ASAP7_75t_SL g244 ( 
.A1(n_239),
.A2(n_201),
.B1(n_205),
.B2(n_212),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_244),
.A2(n_231),
.B1(n_232),
.B2(n_218),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_205),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_245),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_243),
.A2(n_203),
.B(n_201),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_246),
.A2(n_248),
.B(n_252),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_250),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_215),
.B(n_201),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_201),
.B(n_200),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_259),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_195),
.C(n_217),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_260),
.C(n_261),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_191),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_262),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_227),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_188),
.C(n_208),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_188),
.C(n_207),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_228),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_264),
.Y(n_283)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_267),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_263),
.A2(n_244),
.B1(n_220),
.B2(n_245),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_273),
.B1(n_274),
.B2(n_246),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_233),
.C(n_235),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_270),
.C(n_271),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_233),
.C(n_238),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_236),
.C(n_220),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_245),
.A2(n_199),
.B1(n_240),
.B2(n_223),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_260),
.A2(n_230),
.B1(n_198),
.B2(n_219),
.Y(n_274)
);

AOI21xp33_ASAP7_75t_L g276 ( 
.A1(n_251),
.A2(n_226),
.B(n_199),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_276),
.A2(n_4),
.B(n_2),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_256),
.A2(n_198),
.B1(n_237),
.B2(n_241),
.Y(n_277)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_277),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_258),
.B(n_253),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_279),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_228),
.C(n_189),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_11),
.C(n_3),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_261),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_284),
.Y(n_302)
);

BUFx4f_ASAP7_75t_SL g285 ( 
.A(n_283),
.Y(n_285)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_269),
.Y(n_287)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_291),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_275),
.A2(n_252),
.B1(n_249),
.B2(n_255),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_248),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_292),
.A2(n_282),
.B1(n_265),
.B2(n_270),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_193),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_295),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_4),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_297),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_290),
.B(n_271),
.Y(n_298)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_298),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_294),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_295),
.C(n_293),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_278),
.B1(n_272),
.B2(n_281),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_303),
.B(n_292),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_306),
.A2(n_284),
.B(n_282),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_309),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_286),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_313),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_293),
.C(n_266),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_300),
.A2(n_285),
.B(n_274),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_304),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_307),
.A2(n_285),
.B1(n_296),
.B2(n_280),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_301),
.B1(n_305),
.B2(n_280),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_311),
.B(n_306),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_316),
.B(n_310),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_320),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_321),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_323),
.A2(n_319),
.B(n_312),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_324),
.B(n_317),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_325),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_322),
.C(n_326),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_318),
.B1(n_3),
.B2(n_4),
.Y(n_329)
);

BUFx24_ASAP7_75t_SL g330 ( 
.A(n_329),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_2),
.Y(n_331)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_331),
.Y(n_332)
);


endmodule