module fake_jpeg_10525_n_178 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx8_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_6),
.B(n_1),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_35),
.Y(n_58)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_17),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_16),
.Y(n_46)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_15),
.B1(n_16),
.B2(n_29),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_15),
.Y(n_44)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_20),
.B1(n_31),
.B2(n_22),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_50),
.B1(n_63),
.B2(n_19),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_46),
.B(n_25),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_48),
.A2(n_57),
.B1(n_15),
.B2(n_28),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_22),
.B1(n_31),
.B2(n_20),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_30),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_60),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_30),
.B(n_25),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_15),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_34),
.A2(n_29),
.B1(n_18),
.B2(n_30),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

AND2x6_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_2),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_SL g91 ( 
.A(n_66),
.B(n_85),
.C(n_86),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_68),
.Y(n_98)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_17),
.B1(n_40),
.B2(n_19),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_69),
.A2(n_32),
.B(n_27),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_89),
.B1(n_27),
.B2(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_14),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_73),
.B(n_75),
.Y(n_100)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_26),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_76),
.B(n_79),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_35),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_78),
.B(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_12),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_43),
.B1(n_47),
.B2(n_51),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_87),
.B1(n_32),
.B2(n_3),
.Y(n_105)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_2),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_49),
.A2(n_41),
.B1(n_44),
.B2(n_28),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_55),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_32),
.C(n_3),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_32),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_32),
.C(n_3),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_66),
.A2(n_51),
.B1(n_61),
.B2(n_55),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_94),
.B1(n_95),
.B2(n_105),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_99),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_68),
.A2(n_61),
.B1(n_53),
.B2(n_64),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_71),
.B(n_83),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_97),
.B(n_69),
.Y(n_113)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_109),
.Y(n_114)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_104),
.B(n_72),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_11),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_83),
.B(n_2),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_122),
.B(n_124),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_117),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_90),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_119),
.Y(n_137)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_120),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_121),
.A2(n_108),
.B(n_102),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_86),
.C(n_87),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_126),
.C(n_127),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_82),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_70),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_70),
.B(n_99),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_77),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_77),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_126),
.A2(n_104),
.B1(n_105),
.B2(n_96),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_128),
.A2(n_129),
.B1(n_131),
.B2(n_134),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_120),
.A2(n_92),
.B1(n_109),
.B2(n_103),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_123),
.A2(n_112),
.B1(n_122),
.B2(n_116),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_118),
.C(n_114),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_8),
.C(n_130),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_110),
.B1(n_101),
.B2(n_100),
.Y(n_134)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_101),
.C(n_100),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_116),
.C(n_113),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_132),
.C(n_138),
.Y(n_156)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_148),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_140),
.A2(n_127),
.B1(n_115),
.B2(n_107),
.Y(n_147)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_107),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_150),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_10),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_8),
.C(n_9),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_152),
.C(n_139),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g153 ( 
.A(n_143),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_134),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_156),
.C(n_152),
.Y(n_162)
);

OAI21x1_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_128),
.B(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_137),
.Y(n_159)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_163),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_148),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_166),
.A2(n_141),
.B(n_146),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_154),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_170),
.A3(n_129),
.B1(n_142),
.B2(n_155),
.C1(n_137),
.C2(n_8),
.Y(n_174)
);

OAI31xp33_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_145),
.A3(n_133),
.B(n_141),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_151),
.C(n_146),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_167),
.A2(n_166),
.B(n_131),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_172),
.B(n_173),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_174),
.Y(n_176)
);

MAJx2_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_169),
.C(n_168),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_176),
.Y(n_178)
);


endmodule