module real_jpeg_16823_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_SL g16 ( 
.A(n_0),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_18),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_1),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_2),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_3),
.A2(n_93),
.B1(n_96),
.B2(n_97),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_3),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_3),
.A2(n_96),
.B1(n_124),
.B2(n_127),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_3),
.A2(n_96),
.B1(n_137),
.B2(n_139),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_3),
.A2(n_96),
.B1(n_242),
.B2(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_4),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_4),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_4),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_4),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_4),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_5),
.A2(n_137),
.B1(n_283),
.B2(n_285),
.Y(n_282)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_5),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_6),
.A2(n_287),
.B1(n_289),
.B2(n_290),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_6),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_6),
.A2(n_289),
.B1(n_308),
.B2(n_311),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_6),
.A2(n_289),
.B1(n_412),
.B2(n_413),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_6),
.A2(n_289),
.B1(n_440),
.B2(n_441),
.Y(n_439)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g295 ( 
.A(n_7),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_8),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_8),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_8),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_8),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_8),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_9),
.Y(n_236)
);

BUFx8_ASAP7_75t_L g239 ( 
.A(n_9),
.Y(n_239)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_9),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_10),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_10),
.Y(n_216)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_10),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g248 ( 
.A(n_10),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_10),
.Y(n_261)
);

OAI32xp33_ASAP7_75t_L g28 ( 
.A1(n_11),
.A2(n_29),
.A3(n_32),
.B1(n_35),
.B2(n_41),
.Y(n_28)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_11),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_11),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_11),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_11),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_11),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_11),
.B(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_11),
.A2(n_188),
.B1(n_234),
.B2(n_237),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_12),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_13),
.A2(n_15),
.B(n_17),
.Y(n_14)
);

BUFx12f_ASAP7_75t_SL g15 ( 
.A(n_16),
.Y(n_15)
);

AOI21xp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_449),
.B(n_452),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_378),
.B(n_443),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AO221x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_274),
.B1(n_276),
.B2(n_371),
.C(n_377),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_221),
.B(n_273),
.Y(n_22)
);

AOI21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_197),
.B(n_220),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_145),
.B(n_196),
.Y(n_24)
);

NOR2xp67_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_131),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_26),
.B(n_131),
.Y(n_196)
);

XOR2x2_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_68),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_27),
.B(n_100),
.C(n_129),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_47),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_28),
.B(n_47),
.Y(n_200)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_40),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_36),
.A2(n_285),
.B1(n_302),
.B2(n_304),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_38),
.Y(n_312)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_39),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_40),
.B(n_106),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_40),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_41),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_42),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_79)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_56),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g134 ( 
.A1(n_48),
.A2(n_135),
.B1(n_136),
.B2(n_141),
.Y(n_134)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_49),
.B(n_57),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_50),
.A2(n_102),
.B(n_105),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AO22x2_ASAP7_75t_L g118 ( 
.A1(n_52),
.A2(n_114),
.B1(n_119),
.B2(n_121),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_52),
.Y(n_138)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_52),
.Y(n_140)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_52),
.Y(n_177)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_52),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_55),
.Y(n_165)
);

NOR2x1_ASAP7_75t_L g320 ( 
.A(n_56),
.B(n_286),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_63),
.Y(n_56)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_57),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_60),
.Y(n_182)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OA21x2_ASAP7_75t_L g183 ( 
.A1(n_64),
.A2(n_136),
.B(n_184),
.Y(n_183)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_67),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_100),
.B1(n_129),
.B2(n_130),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_69),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_69),
.A2(n_129),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_69),
.B(n_279),
.C(n_280),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_69),
.A2(n_129),
.B1(n_279),
.B2(n_329),
.Y(n_328)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_79),
.B1(n_85),
.B2(n_92),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g204 ( 
.A1(n_70),
.A2(n_79),
.B1(n_85),
.B2(n_92),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_70),
.A2(n_79),
.B(n_85),
.Y(n_342)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_70),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_70),
.B(n_79),
.Y(n_425)
);

NAND2x1p5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_79),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_77),
.Y(n_214)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_78),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_78),
.Y(n_267)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_85),
.Y(n_389)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_89),
.Y(n_414)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx2_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_99),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_100),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_100),
.A2(n_130),
.B1(n_148),
.B2(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_100),
.B(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_100),
.A2(n_130),
.B1(n_335),
.B2(n_363),
.Y(n_362)
);

AO22x2_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_108),
.B1(n_118),
.B2(n_123),
.Y(n_100)
);

AO22x1_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_108),
.B1(n_118),
.B2(n_123),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_101),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_101),
.B(n_299),
.Y(n_317)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI32xp33_ASAP7_75t_L g148 ( 
.A1(n_105),
.A2(n_149),
.A3(n_153),
.B1(n_155),
.B2(n_160),
.Y(n_148)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_108),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_108),
.Y(n_299)
);

NOR2x1p5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_118),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_113),
.B1(n_115),
.B2(n_116),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_112),
.Y(n_306)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_118),
.B(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_118),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_118),
.A2(n_299),
.B1(n_300),
.B2(n_307),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_120),
.Y(n_292)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_129),
.B(n_227),
.C(n_366),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.C(n_143),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_132),
.A2(n_133),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_132),
.B(n_200),
.C(n_202),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_132),
.A2(n_133),
.B1(n_281),
.B2(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_143),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_133),
.B(n_281),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_134),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_134),
.B(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_134),
.B(n_186),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_134),
.A2(n_167),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_135),
.A2(n_282),
.B1(n_286),
.B2(n_293),
.Y(n_281)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_144),
.A2(n_389),
.B1(n_390),
.B2(n_391),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_144),
.A2(n_390),
.B1(n_391),
.B2(n_411),
.Y(n_410)
);

AOI21x1_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_170),
.B(n_195),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_166),
.Y(n_146)
);

NOR2xp67_ASAP7_75t_SL g195 ( 
.A(n_147),
.B(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_167),
.B(n_258),
.Y(n_353)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21x1_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_190),
.B(n_194),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_185),
.B(n_189),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_183),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_177),
.Y(n_284)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_191),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_183),
.B(n_204),
.C(n_208),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_184),
.A2(n_282),
.B(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_188),
.B(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_192),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_219),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_219),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_202),
.B1(n_203),
.B2(n_218),
.Y(n_198)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_200),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_217),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_204),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_204),
.A2(n_298),
.B(n_313),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_204),
.B(n_298),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_204),
.B(n_279),
.C(n_353),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_204),
.A2(n_217),
.B1(n_279),
.B2(n_329),
.Y(n_359)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OA22x2_ASAP7_75t_L g232 ( 
.A1(n_210),
.A2(n_233),
.B1(n_240),
.B2(n_250),
.Y(n_232)
);

OAI21x1_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_241),
.B(n_246),
.Y(n_240)
);

OA22x2_ASAP7_75t_L g279 ( 
.A1(n_210),
.A2(n_233),
.B1(n_240),
.B2(n_250),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_210),
.B(n_240),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_210),
.A2(n_427),
.B(n_432),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_210),
.A2(n_427),
.B1(n_434),
.B2(n_439),
.Y(n_438)
);

OA22x2_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_210)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_211),
.Y(n_394)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_211),
.Y(n_397)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_222),
.B(n_223),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_254),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_224),
.B(n_255),
.C(n_256),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_231),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B(n_230),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_228),
.B(n_229),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_229),
.A2(n_301),
.B(n_317),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_231),
.A2(n_232),
.B1(n_341),
.B2(n_342),
.Y(n_348)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_232),
.Y(n_340)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_232),
.Y(n_366)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_233),
.Y(n_323)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_234),
.Y(n_429)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g242 ( 
.A(n_236),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_236),
.Y(n_441)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_240),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_241),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

INVx5_ASAP7_75t_L g440 ( 
.A(n_242),
.Y(n_440)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_268),
.B1(n_271),
.B2(n_272),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_269),
.A2(n_428),
.B1(n_430),
.B2(n_431),
.Y(n_427)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_354),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_343),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_326),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_277),
.B(n_326),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_296),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_278),
.B(n_297),
.C(n_314),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_279),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_279),
.A2(n_329),
.B1(n_407),
.B2(n_408),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_279),
.B(n_386),
.C(n_436),
.Y(n_435)
);

XNOR2x1_ASAP7_75t_L g327 ( 
.A(n_280),
.B(n_328),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_281),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_285),
.Y(n_303)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_285),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx12f_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_314),
.Y(n_296)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_302),
.A2(n_303),
.B1(n_392),
.B2(n_395),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

AND2x2_ASAP7_75t_SL g386 ( 
.A(n_307),
.B(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_313),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_313),
.A2(n_382),
.B1(n_398),
.B2(n_419),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_321),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g400 ( 
.A(n_315),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_318),
.Y(n_315)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_316),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_318),
.A2(n_319),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_319),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_319),
.A2(n_320),
.B1(n_322),
.B2(n_325),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_319),
.A2(n_325),
.B(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_323),
.B(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_324),
.B(n_451),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_330),
.C(n_333),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_327),
.B(n_330),
.Y(n_345)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_333),
.B(n_345),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_339),
.C(n_341),
.Y(n_333)
);

XNOR2x1_ASAP7_75t_L g347 ( 
.A(n_334),
.B(n_348),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_335),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_340),
.B(n_388),
.C(n_403),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_340),
.A2(n_383),
.B1(n_405),
.B2(n_406),
.Y(n_404)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_343),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_346),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g376 ( 
.A(n_344),
.B(n_346),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.C(n_352),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_350),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2x1_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_353),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_367),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_357),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_360),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_362),
.C(n_364),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_362),
.B1(n_364),
.B2(n_365),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_365),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_366),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_366),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_366),
.B(n_402),
.C(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_367),
.B(n_374),
.Y(n_373)
);

NAND2x1_ASAP7_75t_SL g367 ( 
.A(n_368),
.B(n_370),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_368),
.B(n_370),
.Y(n_372)
);

A2O1A1Ixp33_ASAP7_75t_L g371 ( 
.A1(n_372),
.A2(n_373),
.B(n_375),
.C(n_376),
.Y(n_371)
);

NAND3xp33_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_420),
.C(n_437),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_415),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_380),
.A2(n_445),
.B(n_446),
.Y(n_444)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_401),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_381),
.B(n_401),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_398),
.C(n_399),
.Y(n_381)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_382),
.Y(n_419)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_388),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_386),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_386),
.A2(n_403),
.B1(n_409),
.B2(n_410),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_395),
.Y(n_412)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_399),
.B(n_418),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_402),
.B(n_404),
.Y(n_401)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVxp33_ASAP7_75t_L g422 ( 
.A(n_406),
.Y(n_422)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_409),
.Y(n_436)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_411),
.B(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_417),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g445 ( 
.A(n_416),
.B(n_417),
.Y(n_445)
);

A2O1A1O1Ixp25_ASAP7_75t_L g443 ( 
.A1(n_420),
.A2(n_437),
.B(n_444),
.C(n_447),
.D(n_448),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_421),
.B(n_423),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_423),
.Y(n_447)
);

BUFx24_ASAP7_75t_SL g455 ( 
.A(n_423),
.Y(n_455)
);

FAx1_ASAP7_75t_SL g423 ( 
.A(n_424),
.B(n_426),
.CI(n_435),
.CON(n_423),
.SN(n_423)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_424),
.B(n_426),
.C(n_435),
.Y(n_442)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_430),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_442),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_438),
.B(n_442),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_438),
.B(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_438),
.B(n_450),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_439),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_453),
.Y(n_452)
);


endmodule