module real_jpeg_4510_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g116 ( 
.A(n_0),
.Y(n_116)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_1),
.A2(n_66),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_1),
.A2(n_66),
.B1(n_181),
.B2(n_184),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_1),
.A2(n_66),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_1),
.B(n_80),
.Y(n_242)
);

O2A1O1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_1),
.A2(n_81),
.B(n_259),
.C(n_261),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_1),
.B(n_170),
.C(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_1),
.B(n_153),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_1),
.B(n_38),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_1),
.B(n_172),
.Y(n_326)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_3),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_4),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_4),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_4),
.A2(n_94),
.B1(n_141),
.B2(n_144),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_4),
.A2(n_94),
.B1(n_274),
.B2(n_276),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_4),
.A2(n_94),
.B1(n_297),
.B2(n_299),
.Y(n_296)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_5),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_6),
.Y(n_192)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_7),
.Y(n_101)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_10),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_10),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_10),
.Y(n_97)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_10),
.Y(n_106)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_10),
.Y(n_158)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_11),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_11),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_32),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_12),
.A2(n_27),
.B1(n_184),
.B2(n_215),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_13),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_13),
.A2(n_49),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_13),
.A2(n_49),
.B1(n_82),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_13),
.A2(n_49),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_229),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_227),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_201),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_22),
.B(n_201),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_145),
.C(n_186),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_23),
.B(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_77),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_24),
.B(n_78),
.C(n_107),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_51),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_25),
.B(n_51),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_36),
.B(n_39),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_26),
.A2(n_188),
.B(n_189),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_30),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_31),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_32),
.Y(n_299)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_35),
.Y(n_176)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_35),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_36),
.Y(n_267)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_39),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_45),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_40),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_40),
.B(n_209),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_40),
.A2(n_209),
.B(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_40),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_43),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_44),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_45),
.B(n_190),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_47),
.Y(n_321)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

AO22x1_ASAP7_75t_SL g172 ( 
.A1(n_50),
.A2(n_173),
.B1(n_175),
.B2(n_177),
.Y(n_172)
);

AOI32xp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_58),
.A3(n_61),
.B1(n_64),
.B2(n_67),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_56),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_56),
.Y(n_143)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_57),
.Y(n_135)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_63),
.B(n_66),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_65),
.A2(n_66),
.B(n_157),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g261 ( 
.A1(n_66),
.A2(n_262),
.B(n_264),
.Y(n_261)
);

NAND2xp33_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_73),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AO22x2_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_81),
.B1(n_83),
.B2(n_86),
.Y(n_80)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_107),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_91),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_88),
.Y(n_79)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_80),
.B(n_92),
.Y(n_159)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_88),
.B(n_98),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_100),
.B1(n_102),
.B2(n_104),
.Y(n_99)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_98),
.Y(n_91)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_98),
.B(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_126),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_122),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_115),
.B1(n_117),
.B2(n_120),
.Y(n_110)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_113),
.Y(n_260)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_114),
.Y(n_263)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_116),
.Y(n_200)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_116),
.Y(n_275)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_118),
.Y(n_286)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_119),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_119),
.Y(n_278)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_SL g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_123),
.A2(n_127),
.B(n_153),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_123),
.B(n_127),
.Y(n_337)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_126),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_140),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_128),
.B(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_134),
.B1(n_136),
.B2(n_139),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_140),
.B(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_145),
.B(n_186),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_154),
.C(n_160),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_146),
.A2(n_160),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_146),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_152),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_150),
.B(n_153),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_152),
.B(n_337),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_154),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_159),
.Y(n_154)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_159),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_160),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_178),
.B(n_179),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_180),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_162),
.B(n_196),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_162),
.B(n_273),
.Y(n_272)
);

NOR2x1_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_172),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_166),
.B1(n_170),
.B2(n_171),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_169),
.Y(n_174)
);

INVx4_ASAP7_75t_SL g177 ( 
.A(n_170),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_172),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_172),
.B(n_273),
.Y(n_291)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_SL g175 ( 
.A(n_176),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_178),
.A2(n_214),
.B(n_218),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_178),
.B(n_179),
.Y(n_271)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_183),
.Y(n_265)
);

INVx11_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_193),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_193),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_189),
.B(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_189),
.B(n_295),
.Y(n_325)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_192),
.Y(n_313)
);

AND2x2_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_194),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_195),
.B(n_272),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_219),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_213),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_212),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_206),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_212),
.B(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_218),
.B(n_291),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_225),
.B2(n_226),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_223),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_247),
.B(n_349),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_245),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_231),
.B(n_245),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_236),
.C(n_238),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.C(n_243),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_255),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_243),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_244),
.B(n_311),
.Y(n_323)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_279),
.B(n_348),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_253),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_250),
.B(n_253),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.C(n_268),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_254),
.B(n_344),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_257),
.A2(n_268),
.B1(n_269),
.B2(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_257),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_266),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_258),
.A2(n_266),
.B1(n_339),
.B2(n_340),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_258),
.Y(n_340)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_266),
.Y(n_339)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_342),
.B(n_347),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_330),
.B(n_341),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_305),
.B(n_329),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_292),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_283),
.B(n_292),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_290),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_284),
.A2(n_285),
.B1(n_290),
.B2(n_308),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_290),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_300),
.Y(n_292)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_293),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_312),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_301),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_302),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_302),
.B(n_303),
.C(n_332),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_314),
.B(n_328),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_309),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_309),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_324),
.B(n_327),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_323),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_322),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_326),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_333),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_338),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_336),
.C(n_338),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_346),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_343),
.B(n_346),
.Y(n_347)
);


endmodule