module fake_jpeg_2242_n_60 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_60);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_44;
wire n_28;
wire n_26;
wire n_38;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_9),
.B(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_27),
.Y(n_32)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_1),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_22),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_21),
.B(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_19),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_34),
.Y(n_38)
);

OR2x2_ASAP7_75t_SL g34 ( 
.A(n_30),
.B(n_29),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_19),
.B1(n_21),
.B2(n_20),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_21),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_41),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_30),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_32),
.Y(n_44)
);

NOR4xp25_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_32),
.C(n_33),
.D(n_10),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_44),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_28),
.B1(n_20),
.B2(n_23),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_45),
.B(n_46),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_28),
.C(n_23),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_SL g50 ( 
.A(n_47),
.B(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_47),
.B(n_1),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_50),
.B(n_2),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_49),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_50),
.A2(n_16),
.B1(n_14),
.B2(n_11),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_3),
.B(n_4),
.Y(n_56)
);

FAx1_ASAP7_75t_SL g55 ( 
.A(n_53),
.B(n_54),
.CI(n_51),
.CON(n_55),
.SN(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_56),
.Y(n_57)
);

OAI31xp33_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_5),
.A3(n_6),
.B(n_7),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_58),
.B(n_9),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_7),
.C(n_8),
.Y(n_60)
);


endmodule