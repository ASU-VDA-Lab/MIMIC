module fake_jpeg_14737_n_392 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_392);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_392;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_41),
.B(n_45),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_13),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_43),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_15),
.B(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_51),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_59),
.Y(n_82)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_18),
.B(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_62),
.Y(n_86)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_31),
.B(n_0),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_31),
.B(n_1),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_69),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_73),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_65),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_20),
.B(n_1),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_28),
.B(n_2),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_79),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_38),
.B1(n_28),
.B2(n_37),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_87),
.A2(n_91),
.B(n_108),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_70),
.A2(n_30),
.B1(n_33),
.B2(n_24),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_41),
.B(n_23),
.Y(n_94)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_60),
.A2(n_30),
.B1(n_21),
.B2(n_33),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_96),
.A2(n_112),
.B1(n_114),
.B2(n_121),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_45),
.B(n_34),
.Y(n_97)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_97),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_34),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_104),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_52),
.B(n_40),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_40),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_118),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_55),
.A2(n_33),
.B1(n_24),
.B2(n_21),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_74),
.A2(n_24),
.B1(n_20),
.B2(n_16),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_71),
.A2(n_27),
.B1(n_23),
.B2(n_22),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_43),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_116),
.Y(n_155)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_49),
.B(n_27),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_51),
.A2(n_22),
.B1(n_16),
.B2(n_39),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_56),
.B(n_26),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_124),
.Y(n_159)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_44),
.Y(n_123)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_49),
.B(n_35),
.Y(n_124)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_59),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_128),
.B1(n_6),
.B2(n_7),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_59),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_130),
.Y(n_197)
);

BUFx4f_ASAP7_75t_SL g131 ( 
.A(n_81),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_131),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_80),
.B(n_64),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_133),
.B(n_164),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_100),
.A2(n_17),
.B1(n_6),
.B2(n_7),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_134),
.A2(n_142),
.B1(n_146),
.B2(n_167),
.Y(n_187)
);

INVx6_ASAP7_75t_SL g135 ( 
.A(n_93),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_135),
.B(n_138),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_82),
.B(n_5),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g207 ( 
.A1(n_136),
.A2(n_163),
.B(n_177),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_89),
.A2(n_67),
.B1(n_66),
.B2(n_50),
.Y(n_142)
);

BUFx24_ASAP7_75t_SL g143 ( 
.A(n_99),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_156),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_100),
.A2(n_101),
.B1(n_113),
.B2(n_89),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_147),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_148),
.Y(n_206)
);

INVx11_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_149),
.A2(n_150),
.B1(n_169),
.B2(n_171),
.Y(n_211)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_106),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_86),
.A2(n_53),
.B(n_47),
.C(n_46),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_179),
.B(n_116),
.C(n_103),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_160),
.B(n_173),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_110),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_161),
.Y(n_190)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_84),
.Y(n_162)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_88),
.B(n_8),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_105),
.B(n_35),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_165),
.B(n_166),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_119),
.B(n_128),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_101),
.A2(n_17),
.B1(n_9),
.B2(n_10),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_90),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_95),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_174),
.B1(n_77),
.B2(n_12),
.Y(n_204)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_78),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_172),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_35),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_95),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_87),
.B(n_11),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_111),
.B(n_19),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_114),
.B(n_19),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_92),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_180),
.B(n_188),
.C(n_195),
.Y(n_254)
);

AOI32xp33_ASAP7_75t_L g181 ( 
.A1(n_138),
.A2(n_125),
.A3(n_112),
.B1(n_91),
.B2(n_53),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_181),
.B(n_148),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_79),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_201),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_139),
.A2(n_177),
.B1(n_145),
.B2(n_179),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_186),
.A2(n_222),
.B1(n_161),
.B2(n_147),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_137),
.B(n_63),
.C(n_129),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_189),
.A2(n_144),
.B(n_131),
.Y(n_227)
);

AND2x4_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_85),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_193),
.A2(n_220),
.B(n_217),
.Y(n_247)
);

AO22x1_ASAP7_75t_L g194 ( 
.A1(n_145),
.A2(n_157),
.B1(n_90),
.B2(n_77),
.Y(n_194)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_194),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_35),
.C(n_19),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_202),
.Y(n_224)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_141),
.Y(n_200)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_78),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_151),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_123),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_210),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_204),
.A2(n_153),
.B1(n_171),
.B2(n_144),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_132),
.A2(n_127),
.B1(n_19),
.B2(n_26),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_205),
.A2(n_212),
.B1(n_214),
.B2(n_202),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_154),
.B(n_26),
.C(n_127),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_130),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_136),
.B(n_26),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_149),
.A2(n_26),
.B1(n_12),
.B2(n_11),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_152),
.Y(n_213)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_150),
.A2(n_26),
.B1(n_117),
.B2(n_169),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_136),
.B(n_175),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_140),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_131),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_216),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_175),
.A2(n_135),
.B1(n_165),
.B2(n_156),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_184),
.Y(n_223)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_223),
.Y(n_262)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_193),
.A2(n_176),
.B(n_158),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_226),
.A2(n_236),
.B(n_247),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_227),
.A2(n_194),
.B(n_209),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_229),
.A2(n_190),
.B1(n_219),
.B2(n_192),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_221),
.B(n_153),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_230),
.B(n_232),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_237),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_191),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_234),
.B(n_240),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_186),
.A2(n_130),
.B1(n_147),
.B2(n_140),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_235),
.A2(n_251),
.B1(n_260),
.B2(n_234),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_185),
.B(n_148),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_239),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_148),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_191),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_250),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_201),
.B(n_218),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_195),
.C(n_198),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_193),
.B(n_210),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_259),
.Y(n_280)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_213),
.Y(n_246)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_200),
.Y(n_248)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_193),
.A2(n_217),
.B(n_182),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_249),
.A2(n_258),
.B(n_197),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_206),
.B(n_215),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_252),
.B(n_253),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_190),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_184),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_255),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_208),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_256),
.B(n_257),
.Y(n_289)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_211),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_217),
.B(n_180),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_187),
.A2(n_194),
.B1(n_189),
.B2(n_207),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_261),
.A2(n_272),
.B(n_273),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_188),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_275),
.C(n_277),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_267),
.A2(n_278),
.B1(n_271),
.B2(n_276),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_270),
.B(n_264),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_233),
.A2(n_192),
.B(n_199),
.Y(n_272)
);

AOI32xp33_ASAP7_75t_L g273 ( 
.A1(n_237),
.A2(n_198),
.A3(n_196),
.B1(n_183),
.B2(n_197),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_274),
.A2(n_286),
.B(n_272),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_254),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_244),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_231),
.B(n_225),
.C(n_228),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_281),
.C(n_283),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_225),
.B(n_228),
.C(n_236),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_247),
.B(n_249),
.C(n_233),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_260),
.A2(n_257),
.B1(n_227),
.B2(n_251),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_284),
.A2(n_261),
.B1(n_283),
.B2(n_285),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_238),
.A2(n_239),
.B(n_258),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_287),
.A2(n_292),
.B1(n_288),
.B2(n_289),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_235),
.B(n_255),
.C(n_240),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_290),
.C(n_266),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_224),
.B(n_232),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_256),
.B(n_223),
.Y(n_291)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_291),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_253),
.A2(n_241),
.B1(n_248),
.B2(n_245),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_282),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_293),
.Y(n_328)
);

OA22x2_ASAP7_75t_L g294 ( 
.A1(n_286),
.A2(n_253),
.B1(n_242),
.B2(n_241),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_294),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_284),
.A2(n_245),
.B1(n_246),
.B2(n_269),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_295),
.A2(n_308),
.B(n_297),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_299),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_282),
.A2(n_276),
.B1(n_271),
.B2(n_262),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_300),
.A2(n_305),
.B1(n_307),
.B2(n_315),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_301),
.B(n_309),
.C(n_311),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_291),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_302),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_268),
.B(n_263),
.Y(n_303)
);

INVxp33_ASAP7_75t_L g330 ( 
.A(n_303),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_265),
.B(n_281),
.Y(n_306)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_306),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_279),
.B1(n_265),
.B2(n_270),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_264),
.B(n_275),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_262),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_310),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_312),
.A2(n_298),
.B1(n_293),
.B2(n_294),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_292),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_313),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_290),
.Y(n_314)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_314),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_274),
.A2(n_280),
.B1(n_269),
.B2(n_273),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_280),
.A2(n_233),
.B1(n_285),
.B2(n_261),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_317),
.B1(n_315),
.B2(n_307),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_277),
.B(n_267),
.Y(n_317)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_317),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_268),
.B(n_252),
.Y(n_318)
);

INVxp33_ASAP7_75t_L g338 ( 
.A(n_318),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_264),
.B(n_275),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_319),
.B(n_296),
.C(n_311),
.Y(n_336)
);

AOI21x1_ASAP7_75t_L g321 ( 
.A1(n_294),
.A2(n_308),
.B(n_295),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_321),
.A2(n_332),
.B(n_334),
.Y(n_352)
);

AO22x1_ASAP7_75t_L g322 ( 
.A1(n_294),
.A2(n_298),
.B1(n_316),
.B2(n_305),
.Y(n_322)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_322),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_324),
.B(n_325),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_325),
.A2(n_337),
.B1(n_321),
.B2(n_334),
.Y(n_351)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_306),
.Y(n_333)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_333),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_336),
.B(n_341),
.C(n_304),
.Y(n_343)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_299),
.Y(n_340)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_340),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_296),
.B(n_309),
.C(n_319),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_338),
.B(n_330),
.Y(n_342)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_342),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_343),
.B(n_341),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_326),
.B(n_304),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_345),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_347),
.A2(n_353),
.B1(n_329),
.B2(n_331),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_297),
.Y(n_349)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_349),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_301),
.C(n_336),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_350),
.B(n_355),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_351),
.B(n_354),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_320),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_339),
.A2(n_340),
.B(n_332),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_328),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_326),
.B(n_323),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_320),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_329),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_357),
.B(n_323),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_359),
.B(n_350),
.C(n_335),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_361),
.A2(n_363),
.B(n_358),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_354),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_362),
.B(n_346),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_364),
.B(n_368),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_346),
.B(n_327),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_370),
.B(n_372),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_360),
.A2(n_352),
.B(n_349),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_371),
.A2(n_376),
.B(n_358),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_359),
.B(n_343),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_373),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_367),
.B(n_331),
.C(n_347),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_374),
.B(n_375),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_362),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_380),
.A2(n_348),
.B(n_344),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_369),
.A2(n_365),
.B(n_353),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_381),
.A2(n_374),
.B(n_357),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_378),
.A2(n_356),
.B1(n_367),
.B2(n_366),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_382),
.B(n_383),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_384),
.B(n_351),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_385),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_387),
.Y(n_388)
);

NAND4xp25_ASAP7_75t_SL g389 ( 
.A(n_388),
.B(n_375),
.C(n_386),
.D(n_377),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_389),
.B(n_379),
.C(n_327),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_390),
.B(n_333),
.C(n_370),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_391),
.B(n_348),
.Y(n_392)
);


endmodule