module fake_netlist_1_11623_n_656 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_656);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_656;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
OR2x2_ASAP7_75t_L g78 ( .A(n_39), .B(n_69), .Y(n_78) );
CKINVDCx14_ASAP7_75t_R g79 ( .A(n_15), .Y(n_79) );
CKINVDCx14_ASAP7_75t_R g80 ( .A(n_48), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_10), .Y(n_81) );
INVxp33_ASAP7_75t_L g82 ( .A(n_68), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_5), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_65), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_26), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_23), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_75), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_4), .Y(n_88) );
INVx2_ASAP7_75t_SL g89 ( .A(n_70), .Y(n_89) );
BUFx3_ASAP7_75t_L g90 ( .A(n_72), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_29), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_45), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_27), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_76), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_8), .Y(n_95) );
INVx2_ASAP7_75t_SL g96 ( .A(n_3), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_18), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_44), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_34), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_38), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_52), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_21), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_33), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_77), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_12), .Y(n_105) );
OR2x2_ASAP7_75t_L g106 ( .A(n_4), .B(n_57), .Y(n_106) );
NOR2xp67_ASAP7_75t_L g107 ( .A(n_55), .B(n_11), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_71), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_49), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_74), .Y(n_110) );
INVxp33_ASAP7_75t_L g111 ( .A(n_66), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_64), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_51), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_35), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_14), .Y(n_115) );
INVxp67_ASAP7_75t_L g116 ( .A(n_28), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_20), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_60), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_7), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_61), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_2), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_79), .B(n_0), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_93), .Y(n_123) );
AND2x6_ASAP7_75t_L g124 ( .A(n_90), .B(n_25), .Y(n_124) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_117), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_125) );
AND2x4_ASAP7_75t_L g126 ( .A(n_96), .B(n_1), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_93), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_96), .B(n_3), .Y(n_129) );
OAI22xp5_ASAP7_75t_L g130 ( .A1(n_88), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_88), .B(n_6), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_99), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_84), .Y(n_133) );
AND2x6_ASAP7_75t_L g134 ( .A(n_90), .B(n_36), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_89), .B(n_8), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_109), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_121), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_85), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_117), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_109), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_86), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_87), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_121), .Y(n_145) );
OAI21x1_ASAP7_75t_L g146 ( .A1(n_110), .A2(n_37), .B(n_67), .Y(n_146) );
CKINVDCx16_ASAP7_75t_R g147 ( .A(n_114), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_100), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_89), .B(n_9), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_87), .Y(n_150) );
AND2x6_ASAP7_75t_L g151 ( .A(n_91), .B(n_32), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_94), .B(n_9), .Y(n_152) );
INVx2_ASAP7_75t_SL g153 ( .A(n_110), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_101), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_119), .B(n_10), .Y(n_155) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_119), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_121), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_91), .Y(n_158) );
BUFx3_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_131), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_145), .Y(n_161) );
OR2x2_ASAP7_75t_L g162 ( .A(n_147), .B(n_95), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_158), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_147), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_158), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_158), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_146), .Y(n_167) );
INVx4_ASAP7_75t_L g168 ( .A(n_124), .Y(n_168) );
INVx4_ASAP7_75t_L g169 ( .A(n_124), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_151), .Y(n_170) );
AND2x4_ASAP7_75t_SL g171 ( .A(n_140), .B(n_97), .Y(n_171) );
NAND2xp33_ASAP7_75t_L g172 ( .A(n_151), .B(n_101), .Y(n_172) );
INVx5_ASAP7_75t_L g173 ( .A(n_124), .Y(n_173) );
OR2x6_ASAP7_75t_L g174 ( .A(n_122), .B(n_106), .Y(n_174) );
AND2x6_ASAP7_75t_L g175 ( .A(n_131), .B(n_92), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_127), .B(n_82), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_123), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_146), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_127), .B(n_111), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_123), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_123), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_128), .Y(n_182) );
INVx5_ASAP7_75t_L g183 ( .A(n_124), .Y(n_183) );
INVx2_ASAP7_75t_SL g184 ( .A(n_156), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_133), .B(n_112), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_145), .Y(n_186) );
OR2x6_ASAP7_75t_L g187 ( .A(n_122), .B(n_106), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_128), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_133), .B(n_80), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_145), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_135), .B(n_95), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_128), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_126), .A2(n_105), .B1(n_83), .B2(n_115), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_137), .Y(n_194) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_154), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_145), .Y(n_196) );
INVx2_ASAP7_75t_SL g197 ( .A(n_126), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_126), .B(n_92), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_145), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_137), .Y(n_200) );
INVx4_ASAP7_75t_L g201 ( .A(n_124), .Y(n_201) );
NAND3xp33_ASAP7_75t_L g202 ( .A(n_126), .B(n_121), .C(n_112), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_163), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_163), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_175), .A2(n_198), .B1(n_197), .B2(n_187), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_175), .A2(n_131), .B1(n_151), .B2(n_124), .Y(n_206) );
CKINVDCx8_ASAP7_75t_R g207 ( .A(n_164), .Y(n_207) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_184), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_175), .A2(n_131), .B1(n_151), .B2(n_124), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_168), .Y(n_210) );
OR2x6_ASAP7_75t_L g211 ( .A(n_174), .B(n_130), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_184), .A2(n_155), .B1(n_136), .B2(n_149), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_165), .Y(n_213) );
NOR2xp33_ASAP7_75t_R g214 ( .A(n_164), .B(n_132), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_176), .B(n_139), .Y(n_215) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_189), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_189), .B(n_153), .Y(n_217) );
OAI22xp33_ASAP7_75t_L g218 ( .A1(n_174), .A2(n_125), .B1(n_148), .B2(n_81), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_165), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_166), .Y(n_220) );
OAI22xp33_ASAP7_75t_L g221 ( .A1(n_174), .A2(n_125), .B1(n_129), .B2(n_144), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_166), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_177), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_179), .B(n_135), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_177), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_171), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_175), .A2(n_151), .B1(n_134), .B2(n_139), .Y(n_227) );
INVxp67_ASAP7_75t_SL g228 ( .A(n_160), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_185), .B(n_150), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_174), .B(n_153), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_187), .B(n_142), .Y(n_231) );
INVx5_ASAP7_75t_L g232 ( .A(n_175), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_167), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_171), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_198), .B(n_143), .Y(n_235) );
INVx4_ASAP7_75t_L g236 ( .A(n_173), .Y(n_236) );
BUFx4f_ASAP7_75t_L g237 ( .A(n_175), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_162), .B(n_150), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_180), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_187), .B(n_143), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_180), .Y(n_241) );
INVx2_ASAP7_75t_SL g242 ( .A(n_173), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_167), .Y(n_243) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_168), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_168), .B(n_142), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_187), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_175), .A2(n_152), .B1(n_144), .B2(n_151), .Y(n_247) );
BUFx2_ASAP7_75t_L g248 ( .A(n_169), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_167), .Y(n_249) );
INVx4_ASAP7_75t_L g250 ( .A(n_173), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_169), .B(n_116), .Y(n_251) );
NAND2x1p5_ASAP7_75t_L g252 ( .A(n_169), .B(n_78), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_167), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_201), .B(n_78), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_181), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_205), .A2(n_198), .B1(n_160), .B2(n_197), .Y(n_256) );
AND2x6_ASAP7_75t_L g257 ( .A(n_231), .B(n_160), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_216), .Y(n_258) );
AOI21xp33_ASAP7_75t_L g259 ( .A1(n_247), .A2(n_172), .B(n_202), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g260 ( .A1(n_221), .A2(n_162), .B(n_195), .C(n_198), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_223), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_231), .A2(n_191), .B1(n_193), .B2(n_201), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_238), .A2(n_191), .B(n_200), .C(n_192), .Y(n_263) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_231), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_211), .A2(n_201), .B1(n_159), .B2(n_170), .Y(n_265) );
INVx3_ASAP7_75t_L g266 ( .A(n_203), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g267 ( .A1(n_215), .A2(n_200), .B(n_194), .C(n_192), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_234), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_229), .A2(n_194), .B(n_188), .C(n_182), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_L g270 ( .A1(n_224), .A2(n_188), .B(n_182), .C(n_181), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_208), .B(n_159), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_203), .Y(n_272) );
CKINVDCx11_ASAP7_75t_R g273 ( .A(n_234), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_246), .B(n_170), .Y(n_274) );
BUFx10_ASAP7_75t_L g275 ( .A(n_226), .Y(n_275) );
OR2x6_ASAP7_75t_L g276 ( .A(n_211), .B(n_167), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_223), .Y(n_277) );
BUFx6f_ASAP7_75t_L g278 ( .A(n_210), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_240), .B(n_178), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_240), .B(n_173), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g281 ( .A1(n_235), .A2(n_137), .B1(n_141), .B2(n_178), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_225), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_230), .B(n_173), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_217), .B(n_141), .Y(n_284) );
INVx2_ASAP7_75t_SL g285 ( .A(n_230), .Y(n_285) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_230), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_252), .A2(n_178), .B1(n_118), .B2(n_103), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_225), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_L g289 ( .A1(n_218), .A2(n_118), .B(n_98), .C(n_120), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_213), .A2(n_178), .B(n_107), .C(n_104), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_217), .B(n_121), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_226), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_204), .Y(n_293) );
A2O1A1Ixp33_ASAP7_75t_L g294 ( .A1(n_213), .A2(n_178), .B(n_108), .C(n_113), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_210), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_252), .A2(n_183), .B1(n_173), .B2(n_102), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_239), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_L g298 ( .A1(n_239), .A2(n_183), .B(n_138), .C(n_145), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_L g299 ( .A1(n_254), .A2(n_138), .B(n_196), .C(n_161), .Y(n_299) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_210), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_217), .B(n_183), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_204), .Y(n_302) );
OA21x2_ASAP7_75t_L g303 ( .A1(n_290), .A2(n_253), .B(n_249), .Y(n_303) );
AOI21xp33_ASAP7_75t_L g304 ( .A1(n_260), .A2(n_211), .B(n_212), .Y(n_304) );
OAI21x1_ASAP7_75t_L g305 ( .A1(n_281), .A2(n_249), .B(n_253), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_SL g306 ( .A1(n_269), .A2(n_241), .B(n_255), .C(n_219), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_258), .A2(n_211), .B1(n_252), .B2(n_237), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_291), .Y(n_308) );
OR2x6_ASAP7_75t_L g309 ( .A(n_264), .B(n_248), .Y(n_309) );
OAI21x1_ASAP7_75t_L g310 ( .A1(n_281), .A2(n_243), .B(n_233), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_261), .B(n_220), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_277), .Y(n_312) );
OAI21xp5_ASAP7_75t_L g313 ( .A1(n_279), .A2(n_206), .B(n_209), .Y(n_313) );
AOI21x1_ASAP7_75t_L g314 ( .A1(n_279), .A2(n_233), .B(n_243), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_259), .A2(n_183), .B(n_227), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_284), .Y(n_316) );
AO31x2_ASAP7_75t_L g317 ( .A1(n_294), .A2(n_255), .A3(n_241), .B(n_220), .Y(n_317) );
OA21x2_ASAP7_75t_L g318 ( .A1(n_259), .A2(n_222), .B(n_161), .Y(n_318) );
NAND2x1p5_ASAP7_75t_L g319 ( .A(n_266), .B(n_237), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_278), .Y(n_320) );
INVxp67_ASAP7_75t_SL g321 ( .A(n_286), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_301), .A2(n_183), .B(n_237), .Y(n_322) );
OAI21xp5_ASAP7_75t_L g323 ( .A1(n_267), .A2(n_228), .B(n_245), .Y(n_323) );
OA21x2_ASAP7_75t_L g324 ( .A1(n_298), .A2(n_196), .B(n_199), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_282), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_273), .Y(n_326) );
OAI21x1_ASAP7_75t_L g327 ( .A1(n_270), .A2(n_251), .B(n_199), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_288), .Y(n_328) );
OAI21x1_ASAP7_75t_L g329 ( .A1(n_287), .A2(n_138), .B(n_134), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_262), .A2(n_232), .B1(n_248), .B2(n_207), .Y(n_330) );
OAI21x1_ASAP7_75t_L g331 ( .A1(n_287), .A2(n_138), .B(n_134), .Y(n_331) );
NAND2x1p5_ASAP7_75t_L g332 ( .A(n_266), .B(n_232), .Y(n_332) );
OAI21x1_ASAP7_75t_L g333 ( .A1(n_299), .A2(n_134), .B(n_183), .Y(n_333) );
CKINVDCx8_ASAP7_75t_R g334 ( .A(n_268), .Y(n_334) );
OR2x6_ASAP7_75t_L g335 ( .A(n_276), .B(n_244), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_311), .B(n_297), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_312), .B(n_276), .Y(n_337) );
OAI221xp5_ASAP7_75t_L g338 ( .A1(n_304), .A2(n_289), .B1(n_207), .B2(n_292), .C(n_263), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_312), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_325), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_325), .Y(n_341) );
AOI222xp33_ASAP7_75t_L g342 ( .A1(n_316), .A2(n_256), .B1(n_257), .B2(n_285), .C1(n_275), .C2(n_293), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_307), .A2(n_276), .B1(n_257), .B2(n_256), .Y(n_343) );
INVx4_ASAP7_75t_L g344 ( .A(n_335), .Y(n_344) );
OR2x6_ASAP7_75t_L g345 ( .A(n_335), .B(n_302), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_311), .A2(n_272), .B1(n_302), .B2(n_296), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_328), .B(n_257), .Y(n_347) );
BUFx4f_ASAP7_75t_SL g348 ( .A(n_326), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_314), .Y(n_349) );
AND2x4_ASAP7_75t_L g350 ( .A(n_309), .B(n_300), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_314), .Y(n_351) );
OAI21x1_ASAP7_75t_L g352 ( .A1(n_305), .A2(n_296), .B(n_283), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_309), .A2(n_265), .B1(n_271), .B2(n_274), .Y(n_353) );
OAI21x1_ASAP7_75t_L g354 ( .A1(n_305), .A2(n_280), .B(n_295), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_306), .Y(n_355) );
OAI221xp5_ASAP7_75t_L g356 ( .A1(n_334), .A2(n_214), .B1(n_232), .B2(n_278), .C(n_300), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_309), .A2(n_232), .B1(n_295), .B2(n_278), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_315), .A2(n_210), .B(n_244), .Y(n_358) );
AOI21xp5_ASAP7_75t_L g359 ( .A1(n_318), .A2(n_210), .B(n_244), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_335), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_308), .B(n_257), .Y(n_361) );
OAI21x1_ASAP7_75t_L g362 ( .A1(n_310), .A2(n_300), .B(n_295), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_339), .Y(n_363) );
INVx3_ASAP7_75t_L g364 ( .A(n_350), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_336), .B(n_317), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_349), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_336), .B(n_317), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_339), .B(n_317), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_340), .B(n_317), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_345), .Y(n_370) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_362), .Y(n_371) );
INVx2_ASAP7_75t_SL g372 ( .A(n_350), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_340), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_349), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_349), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_351), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_341), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_341), .B(n_317), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_337), .B(n_313), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_342), .B(n_320), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_351), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_351), .Y(n_382) );
OAI22xp5_ASAP7_75t_SL g383 ( .A1(n_348), .A2(n_326), .B1(n_334), .B2(n_335), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_362), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_337), .B(n_321), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_350), .B(n_318), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_350), .B(n_318), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_354), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_355), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_346), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_357), .Y(n_391) );
AND2x2_ASAP7_75t_SL g392 ( .A(n_344), .B(n_318), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_365), .B(n_354), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_363), .B(n_342), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_366), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_383), .B(n_275), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_371), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_365), .B(n_346), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_367), .B(n_355), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_366), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_367), .B(n_360), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_368), .B(n_360), .Y(n_402) );
NAND4xp25_ASAP7_75t_L g403 ( .A(n_385), .B(n_338), .C(n_343), .D(n_347), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_368), .A2(n_347), .B1(n_361), .B2(n_353), .C(n_344), .Y(n_404) );
INVxp67_ASAP7_75t_SL g405 ( .A(n_381), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_368), .B(n_344), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_363), .B(n_344), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_369), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_369), .Y(n_409) );
INVx1_ASAP7_75t_SL g410 ( .A(n_381), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_369), .B(n_345), .Y(n_411) );
AO21x2_ASAP7_75t_L g412 ( .A1(n_388), .A2(n_359), .B(n_310), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_373), .B(n_361), .Y(n_413) );
OAI221xp5_ASAP7_75t_L g414 ( .A1(n_383), .A2(n_353), .B1(n_345), .B2(n_356), .C(n_330), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_378), .Y(n_415) );
INVx4_ASAP7_75t_L g416 ( .A(n_370), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_378), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_378), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_373), .B(n_345), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_377), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_385), .B(n_345), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_377), .B(n_352), .Y(n_422) );
AOI31xp33_ASAP7_75t_L g423 ( .A1(n_390), .A2(n_357), .A3(n_319), .B(n_332), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_382), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_391), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_386), .B(n_352), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_386), .B(n_303), .Y(n_427) );
OAI221xp5_ASAP7_75t_L g428 ( .A1(n_390), .A2(n_323), .B1(n_309), .B2(n_319), .C(n_303), .Y(n_428) );
NAND3xp33_ASAP7_75t_L g429 ( .A(n_389), .B(n_157), .C(n_303), .Y(n_429) );
INVxp67_ASAP7_75t_SL g430 ( .A(n_382), .Y(n_430) );
OAI31xp33_ASAP7_75t_L g431 ( .A1(n_380), .A2(n_319), .A3(n_332), .B(n_320), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_366), .Y(n_432) );
AND2x2_ASAP7_75t_SL g433 ( .A(n_370), .B(n_303), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_374), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_374), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_408), .B(n_386), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_410), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_395), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_408), .B(n_409), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_425), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_420), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_409), .B(n_379), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_415), .B(n_379), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_396), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_420), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_424), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_424), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_415), .B(n_387), .Y(n_448) );
AND2x4_ASAP7_75t_SL g449 ( .A(n_416), .B(n_364), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_417), .B(n_375), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_423), .B(n_392), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_407), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_413), .Y(n_453) );
NOR2xp67_ASAP7_75t_L g454 ( .A(n_416), .B(n_376), .Y(n_454) );
AND2x4_ASAP7_75t_L g455 ( .A(n_417), .B(n_387), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_410), .Y(n_456) );
NOR2x1_ASAP7_75t_L g457 ( .A(n_423), .B(n_364), .Y(n_457) );
NAND4xp25_ASAP7_75t_SL g458 ( .A(n_404), .B(n_380), .C(n_387), .D(n_376), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_418), .B(n_372), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_418), .B(n_374), .Y(n_460) );
OAI33xp33_ASAP7_75t_L g461 ( .A1(n_394), .A2(n_389), .A3(n_12), .B1(n_13), .B2(n_14), .B3(n_15), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_393), .B(n_392), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_401), .B(n_375), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_401), .B(n_375), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_406), .B(n_364), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_399), .B(n_372), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_399), .B(n_372), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_393), .B(n_392), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_395), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_405), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_430), .Y(n_471) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_403), .A2(n_364), .B1(n_157), .B2(n_388), .C(n_376), .Y(n_472) );
INVxp67_ASAP7_75t_SL g473 ( .A(n_395), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_419), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_419), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_402), .B(n_388), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_398), .B(n_384), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_402), .B(n_11), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_398), .B(n_13), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_432), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_432), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_426), .B(n_384), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_434), .Y(n_483) );
INVxp67_ASAP7_75t_SL g484 ( .A(n_400), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_426), .B(n_384), .Y(n_485) );
NAND2xp33_ASAP7_75t_L g486 ( .A(n_434), .B(n_371), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_427), .B(n_371), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_435), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_400), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_421), .B(n_16), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_406), .B(n_16), .Y(n_491) );
INVx1_ASAP7_75t_SL g492 ( .A(n_440), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_446), .Y(n_493) );
INVx1_ASAP7_75t_SL g494 ( .A(n_456), .Y(n_494) );
NAND2x1p5_ASAP7_75t_L g495 ( .A(n_454), .B(n_416), .Y(n_495) );
NOR2x1_ASAP7_75t_SL g496 ( .A(n_451), .B(n_416), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_447), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_461), .B(n_403), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_471), .B(n_411), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_441), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_463), .B(n_411), .Y(n_501) );
INVx2_ASAP7_75t_SL g502 ( .A(n_437), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_445), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_455), .B(n_397), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_439), .Y(n_505) );
XOR2x1_ASAP7_75t_L g506 ( .A(n_465), .B(n_435), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_439), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_455), .B(n_397), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_470), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_480), .Y(n_510) );
BUFx2_ASAP7_75t_L g511 ( .A(n_455), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_438), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_453), .B(n_427), .Y(n_513) );
INVx1_ASAP7_75t_SL g514 ( .A(n_449), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_474), .B(n_422), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_436), .B(n_422), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_475), .B(n_431), .Y(n_517) );
BUFx2_ASAP7_75t_L g518 ( .A(n_465), .Y(n_518) );
AOI21x1_ASAP7_75t_L g519 ( .A1(n_451), .A2(n_429), .B(n_400), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_452), .B(n_436), .Y(n_520) );
XNOR2x1_ASAP7_75t_L g521 ( .A(n_444), .B(n_17), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_448), .B(n_433), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_481), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_483), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_458), .A2(n_414), .B1(n_431), .B2(n_428), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_448), .B(n_433), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_488), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_438), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_444), .B(n_433), .Y(n_529) );
INVx3_ASAP7_75t_L g530 ( .A(n_449), .Y(n_530) );
AOI221xp5_ASAP7_75t_L g531 ( .A1(n_479), .A2(n_157), .B1(n_429), .B2(n_397), .C(n_371), .Y(n_531) );
NAND2x1_ASAP7_75t_L g532 ( .A(n_457), .B(n_397), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_442), .B(n_412), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_463), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_462), .B(n_412), .Y(n_535) );
NAND4xp25_ASAP7_75t_L g536 ( .A(n_490), .B(n_17), .C(n_18), .D(n_19), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_462), .B(n_412), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_443), .B(n_412), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_472), .A2(n_371), .B1(n_324), .B2(n_134), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_491), .B(n_19), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_477), .B(n_20), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_477), .B(n_371), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_464), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_469), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_469), .B(n_371), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_468), .B(n_157), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_464), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_459), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_498), .A2(n_465), .B1(n_468), .B2(n_478), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_509), .Y(n_550) );
INVx3_ASAP7_75t_L g551 ( .A(n_495), .Y(n_551) );
OAI222xp33_ASAP7_75t_L g552 ( .A1(n_514), .A2(n_466), .B1(n_467), .B2(n_450), .C1(n_460), .C2(n_476), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_511), .B(n_487), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_505), .B(n_485), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_525), .A2(n_476), .B1(n_460), .B2(n_450), .Y(n_555) );
OAI21xp33_ASAP7_75t_SL g556 ( .A1(n_529), .A2(n_473), .B(n_484), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_507), .B(n_485), .Y(n_557) );
NOR2xp67_ASAP7_75t_SL g558 ( .A(n_530), .B(n_320), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_531), .A2(n_486), .B(n_489), .Y(n_559) );
OAI221xp5_ASAP7_75t_L g560 ( .A1(n_498), .A2(n_525), .B1(n_521), .B2(n_536), .C(n_529), .Y(n_560) );
AOI222xp33_ASAP7_75t_L g561 ( .A1(n_540), .A2(n_482), .B1(n_487), .B2(n_486), .C1(n_489), .C2(n_157), .Y(n_561) );
INVxp67_ASAP7_75t_L g562 ( .A(n_502), .Y(n_562) );
NAND4xp25_ASAP7_75t_L g563 ( .A(n_540), .B(n_482), .C(n_358), .D(n_322), .Y(n_563) );
AOI32xp33_ASAP7_75t_L g564 ( .A1(n_521), .A2(n_331), .A3(n_329), .B1(n_333), .B2(n_327), .Y(n_564) );
A2O1A1Ixp33_ASAP7_75t_SL g565 ( .A1(n_546), .A2(n_157), .B(n_24), .C(n_30), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_548), .B(n_324), .Y(n_566) );
OAI21xp5_ASAP7_75t_L g567 ( .A1(n_494), .A2(n_329), .B(n_331), .Y(n_567) );
NOR2x1_ASAP7_75t_L g568 ( .A(n_530), .B(n_324), .Y(n_568) );
OAI21xp5_ASAP7_75t_SL g569 ( .A1(n_530), .A2(n_332), .B(n_190), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_534), .B(n_324), .Y(n_570) );
INVx1_ASAP7_75t_SL g571 ( .A(n_492), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_502), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_518), .B(n_22), .Y(n_573) );
INVxp67_ASAP7_75t_SL g574 ( .A(n_506), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_506), .Y(n_575) );
BUFx2_ASAP7_75t_L g576 ( .A(n_495), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_493), .Y(n_577) );
AOI21xp33_ASAP7_75t_L g578 ( .A1(n_541), .A2(n_31), .B(n_40), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_497), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_543), .B(n_327), .Y(n_580) );
INVx3_ASAP7_75t_L g581 ( .A(n_532), .Y(n_581) );
NOR4xp25_ASAP7_75t_L g582 ( .A(n_517), .B(n_41), .C(n_42), .D(n_43), .Y(n_582) );
INVxp67_ASAP7_75t_L g583 ( .A(n_533), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g584 ( .A1(n_496), .A2(n_134), .B1(n_333), .B2(n_232), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_547), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_500), .Y(n_586) );
NAND3xp33_ASAP7_75t_L g587 ( .A(n_538), .B(n_190), .C(n_186), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_516), .B(n_537), .Y(n_588) );
OA21x2_ASAP7_75t_L g589 ( .A1(n_545), .A2(n_190), .B(n_186), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_520), .A2(n_190), .B1(n_186), .B2(n_50), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_577), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_588), .B(n_535), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_579), .Y(n_593) );
INVxp67_ASAP7_75t_L g594 ( .A(n_572), .Y(n_594) );
BUFx2_ASAP7_75t_L g595 ( .A(n_556), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_586), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_555), .B(n_513), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_550), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_585), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_554), .Y(n_600) );
XNOR2x2_ASAP7_75t_L g601 ( .A(n_571), .B(n_499), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_583), .B(n_515), .Y(n_602) );
AOI21xp33_ASAP7_75t_L g603 ( .A1(n_560), .A2(n_503), .B(n_523), .Y(n_603) );
OAI21xp33_ASAP7_75t_L g604 ( .A1(n_583), .A2(n_522), .B(n_526), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_562), .B(n_501), .Y(n_605) );
OAI22xp33_ASAP7_75t_L g606 ( .A1(n_551), .A2(n_519), .B1(n_510), .B2(n_524), .Y(n_606) );
INVx1_ASAP7_75t_SL g607 ( .A(n_576), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_549), .A2(n_561), .B1(n_574), .B2(n_562), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_575), .Y(n_609) );
OR2x2_ASAP7_75t_L g610 ( .A(n_557), .B(n_542), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_553), .B(n_527), .Y(n_611) );
INVxp33_ASAP7_75t_SL g612 ( .A(n_558), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_580), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_566), .B(n_544), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_551), .B(n_508), .Y(n_615) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_552), .A2(n_508), .B1(n_504), .B2(n_528), .C(n_512), .Y(n_616) );
INVxp67_ASAP7_75t_L g617 ( .A(n_609), .Y(n_617) );
AOI221xp5_ASAP7_75t_L g618 ( .A1(n_603), .A2(n_552), .B1(n_563), .B2(n_582), .C(n_564), .Y(n_618) );
AO22x2_ASAP7_75t_L g619 ( .A1(n_607), .A2(n_581), .B1(n_569), .B2(n_559), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_595), .A2(n_581), .B1(n_504), .B2(n_508), .Y(n_620) );
OAI21xp5_ASAP7_75t_L g621 ( .A1(n_608), .A2(n_559), .B(n_584), .Y(n_621) );
AOI221xp5_ASAP7_75t_SL g622 ( .A1(n_616), .A2(n_573), .B1(n_590), .B2(n_567), .C(n_578), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g623 ( .A1(n_597), .A2(n_570), .B1(n_504), .B2(n_587), .C(n_544), .Y(n_623) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_601), .Y(n_624) );
INVxp67_ASAP7_75t_L g625 ( .A(n_591), .Y(n_625) );
OAI221xp5_ASAP7_75t_L g626 ( .A1(n_604), .A2(n_584), .B1(n_565), .B2(n_568), .C(n_539), .Y(n_626) );
INVx1_ASAP7_75t_SL g627 ( .A(n_612), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_612), .A2(n_528), .B1(n_512), .B2(n_545), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_594), .A2(n_539), .B1(n_190), .B2(n_186), .C(n_589), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_613), .B(n_589), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_594), .A2(n_186), .B1(n_47), .B2(n_53), .C(n_54), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_625), .Y(n_632) );
OAI211xp5_ASAP7_75t_L g633 ( .A1(n_624), .A2(n_615), .B(n_602), .C(n_605), .Y(n_633) );
NOR2xp33_ASAP7_75t_SL g634 ( .A(n_627), .B(n_606), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_619), .A2(n_600), .B1(n_593), .B2(n_596), .C(n_598), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_619), .A2(n_599), .B1(n_606), .B2(n_611), .C(n_615), .Y(n_636) );
OAI211xp5_ASAP7_75t_SL g637 ( .A1(n_617), .A2(n_610), .B(n_614), .C(n_592), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_630), .Y(n_638) );
AOI222xp33_ASAP7_75t_L g639 ( .A1(n_621), .A2(n_134), .B1(n_56), .B2(n_58), .C1(n_59), .C2(n_62), .Y(n_639) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_631), .Y(n_640) );
NAND4xp25_ASAP7_75t_L g641 ( .A(n_636), .B(n_618), .C(n_622), .D(n_620), .Y(n_641) );
AND2x4_ASAP7_75t_L g642 ( .A(n_632), .B(n_628), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_638), .B(n_623), .Y(n_643) );
OAI22xp33_ASAP7_75t_L g644 ( .A1(n_634), .A2(n_626), .B1(n_629), .B2(n_73), .Y(n_644) );
NAND3xp33_ASAP7_75t_SL g645 ( .A(n_635), .B(n_46), .C(n_63), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_642), .Y(n_646) );
NOR2x1_ASAP7_75t_L g647 ( .A(n_645), .B(n_633), .Y(n_647) );
INVx1_ASAP7_75t_SL g648 ( .A(n_643), .Y(n_648) );
OAI22x1_ASAP7_75t_L g649 ( .A1(n_648), .A2(n_641), .B1(n_644), .B2(n_640), .Y(n_649) );
OR2x2_ASAP7_75t_SL g650 ( .A(n_646), .B(n_640), .Y(n_650) );
AOI22xp5_ASAP7_75t_SL g651 ( .A1(n_649), .A2(n_647), .B1(n_639), .B2(n_637), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_650), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_652), .A2(n_236), .B1(n_250), .B2(n_244), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_653), .A2(n_651), .B1(n_250), .B2(n_236), .Y(n_654) );
OAI31xp33_ASAP7_75t_L g655 ( .A1(n_654), .A2(n_242), .A3(n_244), .B(n_236), .Y(n_655) );
AOI21xp33_ASAP7_75t_SL g656 ( .A1(n_655), .A2(n_242), .B(n_250), .Y(n_656) );
endmodule