module fake_jpeg_19802_n_185 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_185);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_31),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g32 ( 
.A(n_26),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_40),
.Y(n_46)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_30),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_47),
.B(n_53),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_26),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_60),
.Y(n_64)
);

CKINVDCx12_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_34),
.Y(n_65)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_29),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_21),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_65),
.Y(n_101)
);

OR2x2_ASAP7_75t_SL g63 ( 
.A(n_49),
.B(n_32),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_68),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_66),
.B(n_71),
.Y(n_93)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

OR2x4_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_32),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_20),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_72),
.B(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_74),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_31),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_0),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_38),
.B1(n_42),
.B2(n_36),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_55),
.B1(n_35),
.B2(n_19),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_20),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_38),
.B1(n_42),
.B2(n_36),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_79),
.A2(n_75),
.B1(n_72),
.B2(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_20),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_80),
.B(n_81),
.Y(n_106)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_16),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_85),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_45),
.A2(n_15),
.B(n_18),
.C(n_25),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_21),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_87),
.C(n_28),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_21),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_57),
.A2(n_19),
.B1(n_14),
.B2(n_35),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_79),
.B1(n_73),
.B2(n_67),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_96),
.A2(n_111),
.B1(n_112),
.B2(n_88),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_104),
.B1(n_107),
.B2(n_110),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_29),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_113),
.Y(n_117)
);

AO22x2_ASAP7_75t_L g100 ( 
.A1(n_63),
.A2(n_28),
.B1(n_22),
.B2(n_24),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_102),
.B(n_77),
.C(n_83),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_64),
.A2(n_23),
.B1(n_16),
.B2(n_25),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_68),
.A2(n_23),
.B1(n_27),
.B2(n_18),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_69),
.A2(n_22),
.B1(n_1),
.B2(n_4),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_22),
.B1(n_1),
.B2(n_5),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_85),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_118),
.C(n_127),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_87),
.C(n_86),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_92),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_120),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_84),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_81),
.B1(n_84),
.B2(n_70),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_130),
.B1(n_110),
.B2(n_111),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_87),
.B(n_86),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_113),
.B1(n_109),
.B2(n_108),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_92),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_128),
.Y(n_139)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_97),
.B(n_1),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_70),
.B(n_77),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_94),
.A2(n_5),
.B(n_6),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_132),
.Y(n_143)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_11),
.Y(n_132)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_144),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_132),
.A2(n_99),
.B1(n_96),
.B2(n_114),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_138),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_124),
.A2(n_95),
.B1(n_93),
.B2(n_105),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_109),
.B1(n_100),
.B2(n_106),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_100),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_145),
.A2(n_123),
.B1(n_121),
.B2(n_108),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_133),
.A2(n_116),
.B(n_128),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_148),
.A2(n_152),
.B(n_156),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_141),
.B(n_131),
.Y(n_149)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_135),
.A2(n_122),
.B(n_116),
.C(n_127),
.D(n_115),
.Y(n_150)
);

XNOR2x1_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_143),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_151),
.A2(n_142),
.B1(n_139),
.B2(n_144),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_126),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_118),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_155),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_123),
.C(n_91),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_123),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_163),
.Y(n_166)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

INVxp33_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_164),
.A2(n_150),
.B(n_159),
.Y(n_167)
);

NAND2xp33_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_138),
.Y(n_165)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_165),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_168),
.C(n_172),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_161),
.A2(n_155),
.B1(n_146),
.B2(n_143),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_157),
.A2(n_153),
.B(n_140),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_171),
.B(n_162),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_134),
.B(n_8),
.Y(n_172)
);

AOI322xp5_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_175),
.A3(n_166),
.B1(n_169),
.B2(n_172),
.C1(n_134),
.C2(n_12),
.Y(n_178)
);

AOI21x1_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_164),
.B(n_160),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_162),
.C(n_158),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_11),
.C(n_13),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_174),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_177),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_179),
.Y(n_181)
);

AOI21x1_ASAP7_75t_L g182 ( 
.A1(n_180),
.A2(n_7),
.B(n_9),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_181),
.C(n_9),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_183),
.A2(n_181),
.B(n_10),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_10),
.Y(n_185)
);


endmodule