module fake_netlist_6_3407_n_1084 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_256, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_255, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_107, n_10, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1084);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_256;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_255;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1084;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_1008;
wire n_465;
wire n_367;
wire n_680;
wire n_760;
wire n_741;
wire n_1027;
wire n_875;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_1079;
wire n_362;
wire n_341;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_898;
wire n_617;
wire n_698;
wire n_1074;
wire n_1032;
wire n_845;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_772;
wire n_656;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_1017;
wire n_1004;
wire n_953;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_757;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_981;
wire n_476;
wire n_880;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_584;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_689;
wire n_354;
wire n_799;
wire n_505;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_834;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_515;
wire n_434;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_598;
wire n_496;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

BUFx2_ASAP7_75t_L g257 ( 
.A(n_33),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_251),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_120),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_9),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_214),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_190),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_205),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_105),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_52),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_256),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_39),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_50),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_176),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_32),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_172),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_163),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_129),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_207),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_250),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_80),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_29),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_130),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_203),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_249),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_247),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_100),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_117),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_145),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_58),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_201),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_162),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_86),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_6),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_252),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_143),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_72),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_15),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_151),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_92),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_156),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_154),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_173),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_192),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_2),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_39),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_10),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_108),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_97),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_113),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_78),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_215),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_191),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_165),
.Y(n_310)
);

BUFx10_ASAP7_75t_L g311 ( 
.A(n_15),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_127),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_169),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_73),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_146),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_152),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_44),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_10),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_55),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_17),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_89),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_268),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_261),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_257),
.B(n_0),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_262),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_278),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_260),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_261),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_271),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_301),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_290),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_294),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_298),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_298),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_317),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_318),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_313),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_316),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_316),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_263),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_284),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_272),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_277),
.B(n_0),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_285),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_280),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_288),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_320),
.Y(n_348)
);

NOR2xp67_ASAP7_75t_L g349 ( 
.A(n_258),
.B(n_1),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_310),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_314),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_258),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_291),
.Y(n_353)
);

NOR2xp67_ASAP7_75t_L g354 ( 
.A(n_275),
.B(n_1),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_281),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_275),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_296),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_302),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_303),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_313),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_281),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_296),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_311),
.B(n_2),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_319),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_355),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_322),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_264),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_340),
.B(n_287),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_360),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_355),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_361),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_361),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_325),
.B(n_343),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_346),
.B(n_311),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_360),
.Y(n_375)
);

BUFx10_ASAP7_75t_L g376 ( 
.A(n_322),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_352),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_326),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_352),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_353),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_326),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_357),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_364),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_357),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_332),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_332),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_364),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_362),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_341),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_362),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_333),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_333),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_323),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_348),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_327),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_358),
.A2(n_344),
.B1(n_348),
.B2(n_324),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_328),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_327),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_359),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_356),
.B(n_274),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_334),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_342),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_330),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_329),
.Y(n_404)
);

INVx5_ASAP7_75t_L g405 ( 
.A(n_324),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_335),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_329),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_330),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_338),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_345),
.Y(n_410)
);

BUFx12f_ASAP7_75t_L g411 ( 
.A(n_363),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_347),
.B(n_319),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_350),
.B(n_321),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_373),
.B(n_363),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_389),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_405),
.B(n_281),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_389),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_367),
.B(n_368),
.Y(n_418)
);

INVx3_ASAP7_75t_R g419 ( 
.A(n_394),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_379),
.Y(n_420)
);

INVx4_ASAP7_75t_SL g421 ( 
.A(n_410),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_370),
.Y(n_422)
);

AND2x2_ASAP7_75t_SL g423 ( 
.A(n_394),
.B(n_281),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_379),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_389),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_396),
.A2(n_349),
.B1(n_354),
.B2(n_265),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_411),
.A2(n_266),
.B1(n_267),
.B2(n_259),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_402),
.Y(n_428)
);

BUFx10_ASAP7_75t_L g429 ( 
.A(n_378),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_405),
.B(n_282),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_402),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_402),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_405),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_405),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_411),
.Y(n_435)
);

OAI22xp33_ASAP7_75t_L g436 ( 
.A1(n_366),
.A2(n_303),
.B1(n_337),
.B2(n_351),
.Y(n_436)
);

INVx6_ASAP7_75t_L g437 ( 
.A(n_405),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_410),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_367),
.B(n_368),
.Y(n_439)
);

INVx5_ASAP7_75t_L g440 ( 
.A(n_379),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_370),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_405),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_370),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_410),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_400),
.B(n_269),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_400),
.B(n_282),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_372),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_369),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_400),
.B(n_282),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_372),
.Y(n_450)
);

AND2x6_ASAP7_75t_L g451 ( 
.A(n_412),
.B(n_282),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_380),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_372),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_365),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_410),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_400),
.B(n_270),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_410),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_365),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_371),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_410),
.B(n_289),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_379),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_403),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_397),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_401),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_379),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_413),
.B(n_273),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_406),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_393),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_371),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_412),
.B(n_331),
.Y(n_470)
);

NAND2x1p5_ASAP7_75t_L g471 ( 
.A(n_403),
.B(n_289),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_408),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_379),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_382),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_381),
.B(n_276),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_384),
.Y(n_476)
);

BUFx10_ASAP7_75t_L g477 ( 
.A(n_386),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_384),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_399),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_418),
.B(n_439),
.Y(n_480)
);

NOR3xp33_ASAP7_75t_L g481 ( 
.A(n_418),
.B(n_374),
.C(n_380),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_414),
.B(n_384),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_422),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_472),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_439),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_423),
.B(n_376),
.Y(n_486)
);

O2A1O1Ixp33_ASAP7_75t_L g487 ( 
.A1(n_446),
.A2(n_408),
.B(n_383),
.C(n_387),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_472),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_423),
.B(n_376),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_470),
.B(n_376),
.Y(n_490)
);

O2A1O1Ixp5_ASAP7_75t_L g491 ( 
.A1(n_446),
.A2(n_384),
.B(n_390),
.C(n_382),
.Y(n_491)
);

O2A1O1Ixp33_ASAP7_75t_L g492 ( 
.A1(n_449),
.A2(n_383),
.B(n_387),
.C(n_377),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_422),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_475),
.B(n_385),
.Y(n_494)
);

NAND2xp33_ASAP7_75t_L g495 ( 
.A(n_451),
.B(n_391),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_470),
.B(n_376),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_392),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_463),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_L g499 ( 
.A1(n_449),
.A2(n_289),
.B1(n_388),
.B2(n_377),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_452),
.B(n_375),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_415),
.B(n_409),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_478),
.B(n_382),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_462),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_470),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_417),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_478),
.B(n_425),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_428),
.B(n_279),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_431),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_478),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_432),
.B(n_390),
.Y(n_510)
);

NOR2xp67_ASAP7_75t_SL g511 ( 
.A(n_437),
.B(n_289),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_451),
.A2(n_388),
.B1(n_311),
.B2(n_336),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_445),
.B(n_283),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_451),
.A2(n_336),
.B1(n_331),
.B2(n_390),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_476),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_456),
.B(n_286),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_476),
.B(n_442),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_476),
.B(n_395),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_427),
.B(n_395),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_429),
.B(n_292),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_476),
.Y(n_521)
);

NOR2x1_ASAP7_75t_R g522 ( 
.A(n_463),
.B(n_293),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_436),
.B(n_295),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_435),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_442),
.B(n_395),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_426),
.B(n_297),
.Y(n_526)
);

O2A1O1Ixp5_ASAP7_75t_L g527 ( 
.A1(n_416),
.A2(n_404),
.B(n_407),
.C(n_398),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_416),
.A2(n_404),
.B(n_398),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_468),
.B(n_398),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_441),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_454),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_429),
.B(n_299),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_451),
.A2(n_304),
.B1(n_305),
.B2(n_300),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_420),
.B(n_404),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_444),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_464),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_429),
.B(n_306),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_477),
.B(n_307),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_454),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_451),
.A2(n_407),
.B1(n_309),
.B2(n_312),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_420),
.B(n_407),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_444),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_420),
.B(n_308),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_458),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_458),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_419),
.B(n_315),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_441),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_464),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_424),
.B(n_47),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_451),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_459),
.B(n_48),
.Y(n_551)
);

NOR2x1p5_ASAP7_75t_L g552 ( 
.A(n_467),
.B(n_3),
.Y(n_552)
);

A2O1A1Ixp33_ASAP7_75t_L g553 ( 
.A1(n_459),
.A2(n_6),
.B(n_4),
.C(n_5),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_494),
.B(n_448),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_509),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_529),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_497),
.Y(n_557)
);

A2O1A1Ixp33_ASAP7_75t_L g558 ( 
.A1(n_480),
.A2(n_469),
.B(n_474),
.C(n_460),
.Y(n_558)
);

OAI21xp33_ASAP7_75t_SL g559 ( 
.A1(n_550),
.A2(n_485),
.B(n_503),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_504),
.B(n_469),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_482),
.B(n_424),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_531),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_513),
.B(n_488),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_509),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_488),
.B(n_424),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_515),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_504),
.B(n_465),
.Y(n_567)
);

NOR3xp33_ASAP7_75t_SL g568 ( 
.A(n_523),
.B(n_467),
.C(n_460),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_536),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_539),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_544),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_515),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_505),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_484),
.B(n_465),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_498),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_505),
.B(n_508),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_519),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_R g578 ( 
.A(n_548),
.B(n_477),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_519),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_500),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_545),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_535),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_517),
.A2(n_434),
.B(n_433),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_483),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_524),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_535),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_501),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_510),
.Y(n_588)
);

HB1xp67_ASAP7_75t_SL g589 ( 
.A(n_481),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_551),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_493),
.Y(n_591)
);

NOR3xp33_ASAP7_75t_SL g592 ( 
.A(n_486),
.B(n_430),
.C(n_477),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_506),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_546),
.B(n_471),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_L g595 ( 
.A1(n_491),
.A2(n_430),
.B(n_438),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_521),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_535),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_551),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_507),
.B(n_465),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_522),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_SL g601 ( 
.A(n_489),
.B(n_444),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_532),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_502),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_530),
.Y(n_604)
);

INVxp67_ASAP7_75t_SL g605 ( 
.A(n_521),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_R g606 ( 
.A(n_520),
.B(n_49),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_535),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_547),
.Y(n_608)
);

AND3x2_ASAP7_75t_SL g609 ( 
.A(n_550),
.B(n_7),
.C(n_8),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_521),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_525),
.A2(n_434),
.B(n_433),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_492),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_521),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_499),
.B(n_473),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_552),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_542),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_487),
.Y(n_617)
);

AOI21xp33_ASAP7_75t_L g618 ( 
.A1(n_559),
.A2(n_526),
.B(n_495),
.Y(n_618)
);

INVx5_ASAP7_75t_L g619 ( 
.A(n_582),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_563),
.B(n_490),
.Y(n_620)
);

OAI21x1_ASAP7_75t_L g621 ( 
.A1(n_595),
.A2(n_527),
.B(n_491),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_586),
.Y(n_622)
);

INVxp67_ASAP7_75t_SL g623 ( 
.A(n_598),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_577),
.B(n_579),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_558),
.A2(n_527),
.B(n_528),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_582),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_571),
.Y(n_627)
);

OA21x2_ASAP7_75t_L g628 ( 
.A1(n_558),
.A2(n_518),
.B(n_534),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_569),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_L g630 ( 
.A1(n_561),
.A2(n_541),
.B(n_549),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_571),
.Y(n_631)
);

OAI21x1_ASAP7_75t_L g632 ( 
.A1(n_583),
.A2(n_543),
.B(n_457),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_560),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_582),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_599),
.A2(n_542),
.B(n_514),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_569),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_593),
.A2(n_542),
.B(n_514),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_603),
.A2(n_542),
.B(n_540),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_598),
.A2(n_499),
.B1(n_512),
.B2(n_540),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_588),
.B(n_481),
.Y(n_640)
);

OAI21x1_ASAP7_75t_L g641 ( 
.A1(n_566),
.A2(n_455),
.B(n_473),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_554),
.B(n_590),
.Y(n_642)
);

INVxp67_ASAP7_75t_SL g643 ( 
.A(n_582),
.Y(n_643)
);

AOI21x1_ASAP7_75t_L g644 ( 
.A1(n_567),
.A2(n_516),
.B(n_511),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_605),
.A2(n_496),
.B(n_444),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_586),
.A2(n_461),
.B(n_471),
.Y(n_646)
);

OAI21x1_ASAP7_75t_L g647 ( 
.A1(n_566),
.A2(n_473),
.B(n_474),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_557),
.B(n_556),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_585),
.Y(n_649)
);

NOR4xp25_ASAP7_75t_L g650 ( 
.A(n_609),
.B(n_553),
.C(n_512),
.D(n_538),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_586),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_585),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_616),
.A2(n_461),
.B(n_440),
.Y(n_653)
);

OAI21x1_ASAP7_75t_L g654 ( 
.A1(n_566),
.A2(n_447),
.B(n_443),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_597),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_573),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_560),
.Y(n_657)
);

A2O1A1Ixp33_ASAP7_75t_L g658 ( 
.A1(n_568),
.A2(n_537),
.B(n_533),
.C(n_443),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_560),
.Y(n_659)
);

OAI21x1_ASAP7_75t_L g660 ( 
.A1(n_572),
.A2(n_450),
.B(n_447),
.Y(n_660)
);

OAI21x1_ASAP7_75t_L g661 ( 
.A1(n_572),
.A2(n_453),
.B(n_450),
.Y(n_661)
);

OAI21x1_ASAP7_75t_L g662 ( 
.A1(n_572),
.A2(n_453),
.B(n_421),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_562),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_614),
.A2(n_617),
.B(n_612),
.Y(n_664)
);

OAI21x1_ASAP7_75t_L g665 ( 
.A1(n_611),
.A2(n_421),
.B(n_461),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_575),
.Y(n_666)
);

NOR2xp67_ASAP7_75t_L g667 ( 
.A(n_575),
.B(n_51),
.Y(n_667)
);

OAI21x1_ASAP7_75t_L g668 ( 
.A1(n_574),
.A2(n_564),
.B(n_555),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_587),
.B(n_7),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_576),
.B(n_461),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_578),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_594),
.B(n_437),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_L g673 ( 
.A1(n_609),
.A2(n_437),
.B1(n_440),
.B2(n_11),
.Y(n_673)
);

A2O1A1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_592),
.A2(n_440),
.B(n_11),
.C(n_8),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_616),
.A2(n_440),
.B(n_421),
.Y(n_675)
);

OAI21x1_ASAP7_75t_L g676 ( 
.A1(n_564),
.A2(n_421),
.B(n_440),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_L g677 ( 
.A1(n_584),
.A2(n_255),
.B(n_54),
.Y(n_677)
);

NAND2x1_ASAP7_75t_L g678 ( 
.A(n_597),
.B(n_53),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_666),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_663),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_656),
.Y(n_681)
);

AO31x2_ASAP7_75t_L g682 ( 
.A1(n_638),
.A2(n_581),
.A3(n_570),
.B(n_584),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_673),
.A2(n_606),
.B1(n_602),
.B2(n_601),
.Y(n_683)
);

A2O1A1Ixp33_ASAP7_75t_L g684 ( 
.A1(n_673),
.A2(n_601),
.B(n_602),
.C(n_555),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_627),
.Y(n_685)
);

BUFx4f_ASAP7_75t_L g686 ( 
.A(n_649),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_L g687 ( 
.A1(n_640),
.A2(n_565),
.B(n_604),
.Y(n_687)
);

AO21x2_ASAP7_75t_L g688 ( 
.A1(n_618),
.A2(n_606),
.B(n_591),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_631),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_642),
.B(n_589),
.Y(n_690)
);

OAI21x1_ASAP7_75t_L g691 ( 
.A1(n_641),
.A2(n_555),
.B(n_591),
.Y(n_691)
);

A2O1A1Ixp33_ASAP7_75t_L g692 ( 
.A1(n_640),
.A2(n_615),
.B(n_608),
.C(n_610),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_659),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_648),
.B(n_600),
.Y(n_694)
);

OAI21x1_ASAP7_75t_L g695 ( 
.A1(n_647),
.A2(n_608),
.B(n_596),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_652),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_618),
.A2(n_607),
.B(n_597),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_639),
.A2(n_580),
.B1(n_610),
.B2(n_596),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_651),
.B(n_578),
.Y(n_699)
);

CKINVDCx11_ASAP7_75t_R g700 ( 
.A(n_671),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_629),
.Y(n_701)
);

AOI22x1_ASAP7_75t_L g702 ( 
.A1(n_664),
.A2(n_596),
.B1(n_613),
.B2(n_610),
.Y(n_702)
);

OAI21x1_ASAP7_75t_L g703 ( 
.A1(n_668),
.A2(n_613),
.B(n_607),
.Y(n_703)
);

BUFx10_ASAP7_75t_L g704 ( 
.A(n_624),
.Y(n_704)
);

O2A1O1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_674),
.A2(n_580),
.B(n_613),
.C(n_13),
.Y(n_705)
);

NOR2x1_ASAP7_75t_R g706 ( 
.A(n_636),
.B(n_607),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_633),
.Y(n_707)
);

OAI21x1_ASAP7_75t_L g708 ( 
.A1(n_665),
.A2(n_57),
.B(n_56),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_657),
.B(n_59),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_654),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_SL g711 ( 
.A(n_671),
.B(n_60),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_624),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_660),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_669),
.Y(n_714)
);

AO21x2_ASAP7_75t_L g715 ( 
.A1(n_625),
.A2(n_62),
.B(n_61),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_670),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_661),
.Y(n_717)
);

OAI21x1_ASAP7_75t_L g718 ( 
.A1(n_632),
.A2(n_64),
.B(n_63),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_620),
.A2(n_623),
.B1(n_639),
.B2(n_637),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_SL g720 ( 
.A(n_651),
.B(n_9),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_664),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_650),
.B(n_12),
.Y(n_722)
);

OAI21x1_ASAP7_75t_L g723 ( 
.A1(n_662),
.A2(n_676),
.B(n_621),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_650),
.B(n_667),
.Y(n_724)
);

OAI21x1_ASAP7_75t_SL g725 ( 
.A1(n_677),
.A2(n_66),
.B(n_65),
.Y(n_725)
);

OAI21xp5_ASAP7_75t_L g726 ( 
.A1(n_635),
.A2(n_68),
.B(n_67),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_651),
.Y(n_727)
);

AOI22x1_ASAP7_75t_L g728 ( 
.A1(n_645),
.A2(n_153),
.B1(n_254),
.B2(n_253),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_677),
.A2(n_628),
.B1(n_625),
.B2(n_672),
.Y(n_729)
);

CKINVDCx12_ASAP7_75t_R g730 ( 
.A(n_619),
.Y(n_730)
);

OA21x2_ASAP7_75t_L g731 ( 
.A1(n_630),
.A2(n_12),
.B(n_13),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_626),
.Y(n_732)
);

A2O1A1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_658),
.A2(n_14),
.B(n_16),
.C(n_17),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_630),
.A2(n_70),
.B(n_69),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_690),
.B(n_643),
.Y(n_735)
);

NAND2xp33_ASAP7_75t_SL g736 ( 
.A(n_679),
.B(n_655),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_680),
.Y(n_737)
);

AOI221xp5_ASAP7_75t_L g738 ( 
.A1(n_733),
.A2(n_646),
.B1(n_678),
.B2(n_622),
.C(n_655),
.Y(n_738)
);

OAI211xp5_ASAP7_75t_SL g739 ( 
.A1(n_683),
.A2(n_622),
.B(n_653),
.C(n_675),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_712),
.B(n_655),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_685),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_712),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_686),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_727),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_700),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_700),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_707),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_690),
.A2(n_634),
.B1(n_626),
.B2(n_628),
.Y(n_748)
);

BUFx2_ASAP7_75t_L g749 ( 
.A(n_696),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_683),
.A2(n_619),
.B1(n_634),
.B2(n_626),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_716),
.B(n_619),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_L g752 ( 
.A1(n_698),
.A2(n_644),
.B1(n_16),
.B2(n_18),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_722),
.A2(n_14),
.B1(n_18),
.B2(n_19),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_681),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_689),
.Y(n_755)
);

INVx4_ASAP7_75t_SL g756 ( 
.A(n_709),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_714),
.B(n_19),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_721),
.B(n_20),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_720),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_SL g760 ( 
.A1(n_726),
.A2(n_74),
.B(n_71),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_686),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_727),
.B(n_75),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_720),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_707),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_701),
.Y(n_765)
);

AOI221xp5_ASAP7_75t_L g766 ( 
.A1(n_733),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.C(n_26),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_693),
.B(n_24),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_697),
.A2(n_77),
.B(n_76),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_709),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_693),
.B(n_25),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_732),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_709),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_705),
.B(n_79),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_682),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_682),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_704),
.B(n_27),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_724),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_682),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_L g779 ( 
.A1(n_711),
.A2(n_731),
.B1(n_687),
.B2(n_694),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_698),
.B(n_684),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_704),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_704),
.B(n_30),
.Y(n_782)
);

INVx1_ASAP7_75t_SL g783 ( 
.A(n_699),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_699),
.B(n_31),
.Y(n_784)
);

INVx8_ASAP7_75t_L g785 ( 
.A(n_730),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_682),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_719),
.A2(n_31),
.B(n_32),
.Y(n_787)
);

NAND2x1_ASAP7_75t_L g788 ( 
.A(n_725),
.B(n_81),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_684),
.B(n_692),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_692),
.B(n_33),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_729),
.A2(n_688),
.B(n_734),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_731),
.B(n_34),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_728),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_SL g794 ( 
.A1(n_731),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_702),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_773),
.A2(n_715),
.B1(n_688),
.B2(n_729),
.Y(n_796)
);

OAI211xp5_ASAP7_75t_SL g797 ( 
.A1(n_753),
.A2(n_710),
.B(n_713),
.C(n_717),
.Y(n_797)
);

OAI221xp5_ASAP7_75t_L g798 ( 
.A1(n_787),
.A2(n_710),
.B1(n_713),
.B2(n_717),
.C(n_715),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_735),
.B(n_706),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_773),
.A2(n_708),
.B1(n_718),
.B2(n_703),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_773),
.A2(n_691),
.B1(n_695),
.B2(n_723),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_766),
.A2(n_780),
.B1(n_753),
.B2(n_763),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_760),
.A2(n_35),
.B(n_36),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_783),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_804)
);

CKINVDCx14_ASAP7_75t_R g805 ( 
.A(n_745),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_791),
.A2(n_83),
.B(n_82),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_741),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_756),
.B(n_84),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_SL g809 ( 
.A1(n_780),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_755),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_766),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_737),
.Y(n_812)
);

AOI221xp5_ASAP7_75t_L g813 ( 
.A1(n_763),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.C(n_44),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_767),
.B(n_85),
.Y(n_814)
);

AO21x2_ASAP7_75t_L g815 ( 
.A1(n_791),
.A2(n_45),
.B(n_46),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_SL g816 ( 
.A1(n_752),
.A2(n_45),
.B1(n_46),
.B2(n_87),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_777),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_817)
);

AOI221xp5_ASAP7_75t_L g818 ( 
.A1(n_779),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.C(n_96),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_759),
.A2(n_98),
.B1(n_99),
.B2(n_101),
.Y(n_819)
);

OAI221xp5_ASAP7_75t_L g820 ( 
.A1(n_772),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.C(n_106),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_769),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_821)
);

INVx4_ASAP7_75t_L g822 ( 
.A(n_785),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_747),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_764),
.Y(n_824)
);

OAI21x1_ASAP7_75t_L g825 ( 
.A1(n_768),
.A2(n_111),
.B(n_112),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_784),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_826)
);

OAI21x1_ASAP7_75t_L g827 ( 
.A1(n_768),
.A2(n_118),
.B(n_119),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_769),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_794),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_794),
.A2(n_128),
.B1(n_131),
.B2(n_132),
.Y(n_830)
);

AOI221xp5_ASAP7_75t_SL g831 ( 
.A1(n_779),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.C(n_136),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_756),
.B(n_137),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_736),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_833)
);

AOI222xp33_ASAP7_75t_L g834 ( 
.A1(n_757),
.A2(n_754),
.B1(n_758),
.B2(n_792),
.C1(n_749),
.C2(n_789),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_771),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_761),
.A2(n_141),
.B1(n_142),
.B2(n_144),
.Y(n_836)
);

BUFx4f_ASAP7_75t_SL g837 ( 
.A(n_765),
.Y(n_837)
);

OAI22xp33_ASAP7_75t_L g838 ( 
.A1(n_790),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_SL g839 ( 
.A1(n_789),
.A2(n_150),
.B1(n_155),
.B2(n_157),
.Y(n_839)
);

OA21x2_ASAP7_75t_L g840 ( 
.A1(n_795),
.A2(n_158),
.B(n_159),
.Y(n_840)
);

OAI221xp5_ASAP7_75t_L g841 ( 
.A1(n_788),
.A2(n_160),
.B1(n_161),
.B2(n_164),
.C(n_166),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_776),
.A2(n_167),
.B1(n_168),
.B2(n_170),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_774),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_744),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_782),
.A2(n_171),
.B1(n_174),
.B2(n_175),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_770),
.B(n_177),
.Y(n_846)
);

AOI221xp5_ASAP7_75t_L g847 ( 
.A1(n_758),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.C(n_181),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_843),
.Y(n_848)
);

OR2x2_ASAP7_75t_L g849 ( 
.A(n_815),
.B(n_786),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_807),
.B(n_810),
.Y(n_850)
);

AOI222xp33_ASAP7_75t_L g851 ( 
.A1(n_802),
.A2(n_754),
.B1(n_756),
.B2(n_793),
.C1(n_743),
.C2(n_785),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_835),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_812),
.B(n_775),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_824),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_815),
.B(n_778),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_823),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_844),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_840),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_834),
.B(n_748),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_840),
.Y(n_860)
);

AOI221xp5_ASAP7_75t_L g861 ( 
.A1(n_813),
.A2(n_751),
.B1(n_742),
.B2(n_785),
.C(n_750),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_796),
.B(n_781),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_799),
.B(n_751),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_798),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_818),
.B(n_781),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_825),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_827),
.Y(n_867)
);

AND2x4_ASAP7_75t_SL g868 ( 
.A(n_808),
.B(n_740),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_818),
.B(n_744),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_800),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_797),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_806),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_808),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_831),
.B(n_762),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_832),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_832),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_797),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_814),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_801),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_806),
.B(n_762),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_803),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_846),
.B(n_740),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_839),
.B(n_738),
.Y(n_883)
);

NOR2x1_ASAP7_75t_SL g884 ( 
.A(n_822),
.B(n_738),
.Y(n_884)
);

BUFx2_ASAP7_75t_SL g885 ( 
.A(n_822),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_839),
.B(n_746),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_841),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_847),
.Y(n_888)
);

OR2x2_ASAP7_75t_L g889 ( 
.A(n_804),
.B(n_182),
.Y(n_889)
);

NOR2x1_ASAP7_75t_SL g890 ( 
.A(n_821),
.B(n_739),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_809),
.B(n_829),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_847),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_828),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_837),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_830),
.B(n_183),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_813),
.B(n_184),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_838),
.B(n_185),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_826),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_816),
.B(n_186),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_852),
.Y(n_900)
);

OAI31xp33_ASAP7_75t_L g901 ( 
.A1(n_881),
.A2(n_820),
.A3(n_811),
.B(n_836),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_848),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_852),
.Y(n_903)
);

OAI33xp33_ASAP7_75t_L g904 ( 
.A1(n_881),
.A2(n_739),
.A3(n_816),
.B1(n_805),
.B2(n_819),
.B3(n_817),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_848),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_849),
.B(n_833),
.Y(n_906)
);

AOI221x1_ASAP7_75t_L g907 ( 
.A1(n_888),
.A2(n_845),
.B1(n_842),
.B2(n_189),
.C(n_193),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_852),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_854),
.Y(n_909)
);

OAI21x1_ASAP7_75t_L g910 ( 
.A1(n_860),
.A2(n_187),
.B(n_188),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_849),
.B(n_194),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_857),
.B(n_195),
.Y(n_912)
);

AOI33xp33_ASAP7_75t_L g913 ( 
.A1(n_864),
.A2(n_196),
.A3(n_197),
.B1(n_198),
.B2(n_199),
.B3(n_200),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_854),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_850),
.B(n_202),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_854),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_850),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_863),
.B(n_204),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_856),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_856),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_856),
.Y(n_921)
);

AOI33xp33_ASAP7_75t_L g922 ( 
.A1(n_864),
.A2(n_206),
.A3(n_208),
.B1(n_209),
.B2(n_210),
.B3(n_211),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_853),
.Y(n_923)
);

OAI33xp33_ASAP7_75t_L g924 ( 
.A1(n_888),
.A2(n_212),
.A3(n_213),
.B1(n_216),
.B2(n_217),
.B3(n_218),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_894),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_859),
.B(n_219),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_892),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_853),
.Y(n_928)
);

OAI33xp33_ASAP7_75t_L g929 ( 
.A1(n_892),
.A2(n_223),
.A3(n_224),
.B1(n_225),
.B2(n_226),
.B3(n_227),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_860),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_860),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_923),
.B(n_870),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_919),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_928),
.B(n_879),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_909),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_925),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_917),
.B(n_870),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_925),
.B(n_870),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_903),
.B(n_879),
.Y(n_939)
);

XOR2x2_ASAP7_75t_L g940 ( 
.A(n_926),
.B(n_886),
.Y(n_940)
);

INVxp67_ASAP7_75t_SL g941 ( 
.A(n_920),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_909),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_911),
.B(n_859),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_914),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_914),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_930),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_903),
.B(n_862),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_920),
.B(n_858),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_916),
.B(n_862),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_930),
.B(n_866),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_911),
.B(n_872),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_916),
.B(n_855),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_908),
.Y(n_953)
);

BUFx2_ASAP7_75t_L g954 ( 
.A(n_908),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_921),
.B(n_858),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_921),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_931),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_902),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_931),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_958),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_947),
.B(n_949),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_947),
.B(n_900),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_958),
.Y(n_963)
);

INVxp67_ASAP7_75t_SL g964 ( 
.A(n_933),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_935),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_939),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_943),
.B(n_902),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_935),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_939),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_942),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_949),
.B(n_905),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_SL g972 ( 
.A(n_936),
.B(n_894),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_932),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_942),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_961),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_967),
.B(n_951),
.Y(n_976)
);

INVxp67_ASAP7_75t_L g977 ( 
.A(n_964),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_961),
.B(n_940),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_R g979 ( 
.A(n_972),
.B(n_886),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_962),
.B(n_938),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_973),
.B(n_940),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_962),
.B(n_938),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_971),
.B(n_937),
.Y(n_983)
);

AO21x1_ASAP7_75t_L g984 ( 
.A1(n_960),
.A2(n_955),
.B(n_934),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_971),
.B(n_937),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_960),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_966),
.B(n_894),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_987),
.B(n_969),
.Y(n_988)
);

OAI22xp33_ASAP7_75t_L g989 ( 
.A1(n_981),
.A2(n_906),
.B1(n_887),
.B2(n_898),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_986),
.Y(n_990)
);

AND2x2_ASAP7_75t_SL g991 ( 
.A(n_978),
.B(n_913),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_977),
.A2(n_904),
.B1(n_883),
.B2(n_891),
.Y(n_992)
);

OAI321xp33_ASAP7_75t_L g993 ( 
.A1(n_977),
.A2(n_883),
.A3(n_906),
.B1(n_899),
.B2(n_896),
.C(n_887),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_979),
.B(n_932),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_987),
.Y(n_995)
);

AOI221xp5_ASAP7_75t_L g996 ( 
.A1(n_979),
.A2(n_899),
.B1(n_924),
.B2(n_929),
.C(n_891),
.Y(n_996)
);

NAND3xp33_ASAP7_75t_SL g997 ( 
.A(n_992),
.B(n_984),
.C(n_901),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_995),
.Y(n_998)
);

OAI32xp33_ASAP7_75t_SL g999 ( 
.A1(n_991),
.A2(n_976),
.A3(n_975),
.B1(n_985),
.B2(n_963),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_990),
.Y(n_1000)
);

AOI32xp33_ASAP7_75t_L g1001 ( 
.A1(n_989),
.A2(n_993),
.A3(n_996),
.B1(n_994),
.B2(n_988),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_990),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_1000),
.Y(n_1003)
);

NAND2xp33_ASAP7_75t_SL g1004 ( 
.A(n_997),
.B(n_999),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_998),
.B(n_980),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_1002),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_1001),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_1003),
.B(n_982),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_1005),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_1006),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_1004),
.A2(n_1007),
.B(n_922),
.C(n_887),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_1003),
.B(n_963),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_1003),
.B(n_968),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_1007),
.B(n_983),
.Y(n_1014)
);

AOI222xp33_ASAP7_75t_L g1015 ( 
.A1(n_1011),
.A2(n_895),
.B1(n_874),
.B2(n_884),
.C1(n_918),
.C2(n_898),
.Y(n_1015)
);

NAND4xp25_ASAP7_75t_L g1016 ( 
.A(n_1014),
.B(n_907),
.C(n_851),
.D(n_861),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_1010),
.A2(n_907),
.B(n_912),
.Y(n_1017)
);

AOI211xp5_ASAP7_75t_SL g1018 ( 
.A1(n_1009),
.A2(n_889),
.B(n_927),
.C(n_897),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_1008),
.Y(n_1019)
);

OAI221xp5_ASAP7_75t_L g1020 ( 
.A1(n_1013),
.A2(n_1012),
.B1(n_851),
.B2(n_889),
.C(n_897),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_R g1021 ( 
.A(n_1019),
.B(n_228),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1020),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_1017),
.A2(n_895),
.B(n_898),
.C(n_874),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_1016),
.A2(n_915),
.B1(n_885),
.B2(n_965),
.Y(n_1024)
);

AOI221xp5_ASAP7_75t_L g1025 ( 
.A1(n_1015),
.A2(n_974),
.B1(n_965),
.B2(n_970),
.C(n_915),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_1018),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_R g1027 ( 
.A(n_1019),
.B(n_229),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_1019),
.A2(n_885),
.B1(n_974),
.B2(n_880),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_1026),
.B(n_1022),
.Y(n_1029)
);

NAND2x1p5_ASAP7_75t_L g1030 ( 
.A(n_1024),
.B(n_910),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_1025),
.A2(n_865),
.B1(n_869),
.B2(n_893),
.Y(n_1031)
);

NOR3x1_ASAP7_75t_L g1032 ( 
.A(n_1021),
.B(n_1027),
.C(n_1023),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_1028),
.B(n_941),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1026),
.Y(n_1034)
);

NAND4xp75_ASAP7_75t_L g1035 ( 
.A(n_1022),
.B(n_865),
.C(n_869),
.D(n_880),
.Y(n_1035)
);

NAND4xp75_ASAP7_75t_L g1036 ( 
.A(n_1022),
.B(n_952),
.C(n_893),
.D(n_882),
.Y(n_1036)
);

NAND4xp25_ASAP7_75t_L g1037 ( 
.A(n_1022),
.B(n_878),
.C(n_873),
.D(n_876),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_R g1038 ( 
.A(n_1026),
.B(n_230),
.Y(n_1038)
);

NOR3x1_ASAP7_75t_L g1039 ( 
.A(n_1022),
.B(n_910),
.C(n_954),
.Y(n_1039)
);

NAND3x1_ASAP7_75t_SL g1040 ( 
.A(n_1021),
.B(n_952),
.C(n_884),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1034),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_L g1042 ( 
.A(n_1029),
.B(n_878),
.C(n_875),
.Y(n_1042)
);

NAND3xp33_ASAP7_75t_SL g1043 ( 
.A(n_1038),
.B(n_876),
.C(n_875),
.Y(n_1043)
);

NAND4xp25_ASAP7_75t_SL g1044 ( 
.A(n_1031),
.B(n_876),
.C(n_875),
.D(n_873),
.Y(n_1044)
);

AOI21xp33_ASAP7_75t_SL g1045 ( 
.A1(n_1030),
.A2(n_231),
.B(n_232),
.Y(n_1045)
);

OA22x2_ASAP7_75t_L g1046 ( 
.A1(n_1033),
.A2(n_954),
.B1(n_953),
.B2(n_956),
.Y(n_1046)
);

OAI221xp5_ASAP7_75t_L g1047 ( 
.A1(n_1037),
.A2(n_873),
.B1(n_955),
.B2(n_878),
.C(n_948),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_1040),
.A2(n_866),
.B1(n_867),
.B2(n_871),
.Y(n_1048)
);

NAND3x1_ASAP7_75t_L g1049 ( 
.A(n_1032),
.B(n_957),
.C(n_956),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_1039),
.A2(n_944),
.B(n_945),
.C(n_877),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1035),
.B(n_944),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_L g1052 ( 
.A(n_1036),
.B(n_866),
.C(n_867),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_1034),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1034),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_1034),
.A2(n_867),
.B1(n_871),
.B2(n_877),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_1053),
.B(n_950),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_1041),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_1049),
.Y(n_1058)
);

NAND3xp33_ASAP7_75t_L g1059 ( 
.A(n_1054),
.B(n_948),
.C(n_945),
.Y(n_1059)
);

AND4x1_ASAP7_75t_L g1060 ( 
.A(n_1050),
.B(n_233),
.C(n_234),
.D(n_235),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_1046),
.B(n_957),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_1043),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_1045),
.A2(n_1051),
.B(n_1055),
.C(n_1052),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1058),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1057),
.B(n_1042),
.Y(n_1065)
);

XNOR2x1_ASAP7_75t_L g1066 ( 
.A(n_1062),
.B(n_1044),
.Y(n_1066)
);

OAI22x1_ASAP7_75t_L g1067 ( 
.A1(n_1060),
.A2(n_1048),
.B1(n_1047),
.B2(n_957),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_1063),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_1056),
.A2(n_950),
.B1(n_959),
.B2(n_946),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1064),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_1066),
.A2(n_1061),
.B(n_1059),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_SL g1072 ( 
.A1(n_1065),
.A2(n_890),
.B(n_946),
.Y(n_1072)
);

NAND3xp33_ASAP7_75t_L g1073 ( 
.A(n_1068),
.B(n_950),
.C(n_905),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1070),
.B(n_1067),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_1071),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1075),
.B(n_1074),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1074),
.A2(n_1072),
.B(n_1073),
.Y(n_1077)
);

AOI222xp33_ASAP7_75t_SL g1078 ( 
.A1(n_1075),
.A2(n_1069),
.B1(n_959),
.B2(n_239),
.C1(n_240),
.C2(n_241),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_1078),
.A2(n_950),
.B1(n_868),
.B2(n_855),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1076),
.A2(n_868),
.B1(n_890),
.B2(n_242),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_L g1081 ( 
.A1(n_1080),
.A2(n_1077),
.B1(n_868),
.B2(n_243),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_1079),
.Y(n_1082)
);

AOI221xp5_ASAP7_75t_L g1083 ( 
.A1(n_1082),
.A2(n_1081),
.B1(n_237),
.B2(n_244),
.C(n_245),
.Y(n_1083)
);

OAI31xp33_ASAP7_75t_L g1084 ( 
.A1(n_1083),
.A2(n_236),
.A3(n_246),
.B(n_248),
.Y(n_1084)
);


endmodule