module fake_aes_9368_n_633 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_633);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_633;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_599;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_73;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g73 ( .A(n_9), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_70), .Y(n_74) );
CKINVDCx20_ASAP7_75t_R g75 ( .A(n_2), .Y(n_75) );
INVx1_ASAP7_75t_SL g76 ( .A(n_18), .Y(n_76) );
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_61), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_24), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_38), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_15), .Y(n_80) );
INVxp67_ASAP7_75t_L g81 ( .A(n_68), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_7), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_17), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_32), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_15), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_46), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_6), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_0), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_65), .Y(n_89) );
NOR2xp67_ASAP7_75t_L g90 ( .A(n_51), .B(n_43), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_62), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_26), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_13), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_50), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_54), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_66), .Y(n_96) );
CKINVDCx14_ASAP7_75t_R g97 ( .A(n_36), .Y(n_97) );
CKINVDCx16_ASAP7_75t_R g98 ( .A(n_47), .Y(n_98) );
NOR2xp67_ASAP7_75t_L g99 ( .A(n_30), .B(n_60), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_28), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_11), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_22), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_49), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_53), .Y(n_104) );
INVx2_ASAP7_75t_SL g105 ( .A(n_0), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_67), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_20), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_71), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_16), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_6), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_23), .Y(n_111) );
BUFx2_ASAP7_75t_SL g112 ( .A(n_25), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_35), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_52), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_34), .Y(n_115) );
INVxp33_ASAP7_75t_SL g116 ( .A(n_64), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_10), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_87), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_79), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_87), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_79), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_74), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_96), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_96), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_78), .B(n_83), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_98), .B(n_1), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
BUFx2_ASAP7_75t_L g128 ( .A(n_73), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_105), .B(n_1), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_89), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_97), .B(n_2), .Y(n_131) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_95), .A2(n_33), .B(n_69), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_105), .B(n_3), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_117), .B(n_3), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_80), .B(n_4), .Y(n_135) );
BUFx3_ASAP7_75t_L g136 ( .A(n_100), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_104), .Y(n_137) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_73), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_106), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_93), .Y(n_140) );
BUFx2_ASAP7_75t_L g141 ( .A(n_93), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_107), .B(n_4), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_113), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_114), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_115), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_82), .Y(n_146) );
BUFx3_ASAP7_75t_L g147 ( .A(n_91), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_81), .B(n_5), .Y(n_148) );
NOR2xp33_ASAP7_75t_SL g149 ( .A(n_77), .B(n_72), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_85), .B(n_5), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_88), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_102), .B(n_7), .Y(n_152) );
OAI22xp5_ASAP7_75t_SL g153 ( .A1(n_75), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_110), .B(n_8), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_77), .B(n_11), .Y(n_155) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_75), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_92), .B(n_12), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_112), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_128), .B(n_92), .Y(n_159) );
AOI22xp33_ASAP7_75t_L g160 ( .A1(n_146), .A2(n_116), .B1(n_111), .B2(n_76), .Y(n_160) );
BUFx4f_ASAP7_75t_L g161 ( .A(n_131), .Y(n_161) );
INVx4_ASAP7_75t_L g162 ( .A(n_144), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_128), .B(n_109), .Y(n_163) );
INVx5_ASAP7_75t_L g164 ( .A(n_123), .Y(n_164) );
INVx2_ASAP7_75t_SL g165 ( .A(n_147), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_141), .B(n_109), .Y(n_166) );
INVx2_ASAP7_75t_SL g167 ( .A(n_141), .Y(n_167) );
INVx4_ASAP7_75t_SL g168 ( .A(n_136), .Y(n_168) );
INVx2_ASAP7_75t_SL g169 ( .A(n_147), .Y(n_169) );
AND2x6_ASAP7_75t_L g170 ( .A(n_131), .B(n_116), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_158), .B(n_108), .Y(n_171) );
NAND2xp33_ASAP7_75t_L g172 ( .A(n_158), .B(n_108), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_123), .Y(n_173) );
AND2x2_ASAP7_75t_SL g174 ( .A(n_149), .B(n_94), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_140), .B(n_138), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_147), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_129), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_123), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_140), .B(n_103), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_129), .Y(n_180) );
AND2x6_ASAP7_75t_L g181 ( .A(n_150), .B(n_94), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_123), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_123), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_133), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_133), .Y(n_185) );
INVx2_ASAP7_75t_SL g186 ( .A(n_157), .Y(n_186) );
INVx4_ASAP7_75t_L g187 ( .A(n_144), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_122), .B(n_103), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_146), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_157), .B(n_101), .Y(n_190) );
OAI22xp33_ASAP7_75t_L g191 ( .A1(n_134), .A2(n_101), .B1(n_86), .B2(n_90), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_146), .Y(n_192) );
INVx2_ASAP7_75t_SL g193 ( .A(n_136), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_122), .B(n_86), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_146), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_136), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_127), .B(n_99), .Y(n_197) );
HB1xp67_ASAP7_75t_SL g198 ( .A(n_156), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_127), .B(n_12), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_144), .B(n_137), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_123), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_124), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_150), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_154), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_124), .Y(n_205) );
OR2x2_ASAP7_75t_L g206 ( .A(n_151), .B(n_13), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_124), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_137), .B(n_14), .Y(n_208) );
AND2x6_ASAP7_75t_L g209 ( .A(n_154), .B(n_42), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_144), .B(n_41), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_192), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_177), .B(n_145), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_192), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_162), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_180), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_184), .B(n_126), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_162), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_161), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_185), .B(n_145), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_171), .B(n_179), .Y(n_220) );
BUFx2_ASAP7_75t_L g221 ( .A(n_161), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_203), .A2(n_125), .B(n_143), .C(n_130), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_176), .B(n_149), .Y(n_223) );
NOR2x1p5_ASAP7_75t_L g224 ( .A(n_175), .B(n_155), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_162), .B(n_143), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_187), .B(n_155), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_206), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_170), .A2(n_152), .B1(n_148), .B2(n_153), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_174), .A2(n_135), .B1(n_134), .B2(n_153), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_186), .B(n_135), .Y(n_230) );
BUFx3_ASAP7_75t_L g231 ( .A(n_176), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_188), .B(n_130), .Y(n_232) );
BUFx3_ASAP7_75t_L g233 ( .A(n_209), .Y(n_233) );
INVx4_ASAP7_75t_L g234 ( .A(n_187), .Y(n_234) );
INVx8_ASAP7_75t_L g235 ( .A(n_170), .Y(n_235) );
NAND2x1p5_ASAP7_75t_L g236 ( .A(n_187), .B(n_142), .Y(n_236) );
OR2x2_ASAP7_75t_L g237 ( .A(n_167), .B(n_151), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_189), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g239 ( .A1(n_174), .A2(n_139), .B1(n_130), .B2(n_151), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_204), .B(n_120), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_188), .B(n_139), .Y(n_241) );
BUFx8_ASAP7_75t_L g242 ( .A(n_181), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_171), .B(n_139), .Y(n_243) );
AND2x4_ASAP7_75t_L g244 ( .A(n_159), .B(n_120), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_178), .Y(n_245) );
INVxp67_ASAP7_75t_L g246 ( .A(n_198), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_163), .B(n_118), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_166), .B(n_118), .Y(n_248) );
NOR2xp67_ASAP7_75t_L g249 ( .A(n_197), .B(n_121), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_195), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_178), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_170), .B(n_121), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_168), .B(n_124), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_182), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_170), .B(n_121), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_170), .A2(n_119), .B1(n_124), .B2(n_132), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_194), .A2(n_160), .B1(n_191), .B2(n_190), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_172), .A2(n_119), .B(n_132), .C(n_14), .Y(n_258) );
NAND3xp33_ASAP7_75t_SL g259 ( .A(n_160), .B(n_119), .C(n_132), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_182), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_168), .B(n_124), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_209), .A2(n_132), .B1(n_21), .B2(n_27), .Y(n_262) );
INVxp67_ASAP7_75t_L g263 ( .A(n_194), .Y(n_263) );
NAND2xp33_ASAP7_75t_L g264 ( .A(n_209), .B(n_19), .Y(n_264) );
INVx5_ASAP7_75t_L g265 ( .A(n_209), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_193), .B(n_29), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_169), .B(n_31), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_215), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_212), .B(n_172), .Y(n_269) );
INVx2_ASAP7_75t_SL g270 ( .A(n_219), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_234), .B(n_168), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_226), .A2(n_193), .B(n_196), .Y(n_272) );
AOI22xp33_ASAP7_75t_SL g273 ( .A1(n_229), .A2(n_181), .B1(n_209), .B2(n_191), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_234), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_230), .B(n_181), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_233), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_226), .A2(n_165), .B(n_200), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_263), .B(n_181), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_225), .A2(n_165), .B(n_200), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_L g280 ( .A1(n_220), .A2(n_208), .B(n_199), .C(n_210), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_244), .B(n_181), .Y(n_281) );
O2A1O1Ixp33_ASAP7_75t_L g282 ( .A1(n_257), .A2(n_210), .B(n_183), .C(n_201), .Y(n_282) );
BUFx12f_ASAP7_75t_L g283 ( .A(n_242), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_263), .B(n_183), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_265), .B(n_164), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_265), .B(n_164), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_224), .Y(n_287) );
AND2x6_ASAP7_75t_L g288 ( .A(n_235), .B(n_205), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_235), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_225), .A2(n_207), .B(n_201), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_235), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_265), .B(n_164), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_216), .A2(n_164), .B1(n_173), .B2(n_207), .Y(n_293) );
AO21x1_ASAP7_75t_L g294 ( .A1(n_258), .A2(n_173), .B(n_205), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_259), .A2(n_205), .B(n_202), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_259), .A2(n_205), .B(n_202), .Y(n_296) );
O2A1O1Ixp33_ASAP7_75t_L g297 ( .A1(n_222), .A2(n_202), .B(n_39), .C(n_40), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_237), .Y(n_298) );
NOR3xp33_ASAP7_75t_SL g299 ( .A(n_239), .B(n_37), .C(n_44), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_244), .B(n_202), .Y(n_300) );
NAND3xp33_ASAP7_75t_SL g301 ( .A(n_228), .B(n_45), .C(n_48), .Y(n_301) );
INVx5_ASAP7_75t_L g302 ( .A(n_265), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_232), .A2(n_55), .B(n_56), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_216), .B(n_57), .Y(n_304) );
NOR2xp67_ASAP7_75t_L g305 ( .A(n_246), .B(n_63), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_231), .B(n_58), .Y(n_306) );
O2A1O1Ixp33_ASAP7_75t_L g307 ( .A1(n_247), .A2(n_59), .B(n_248), .C(n_227), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_220), .B(n_243), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_240), .A2(n_242), .B1(n_243), .B2(n_252), .Y(n_309) );
A2O1A1Ixp33_ASAP7_75t_L g310 ( .A1(n_258), .A2(n_241), .B(n_238), .C(n_250), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_240), .B(n_249), .Y(n_311) );
A2O1A1Ixp33_ASAP7_75t_L g312 ( .A1(n_255), .A2(n_256), .B(n_264), .C(n_267), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_214), .Y(n_313) );
BUFx12f_ASAP7_75t_L g314 ( .A(n_218), .Y(n_314) );
AO31x2_ASAP7_75t_L g315 ( .A1(n_294), .A2(n_267), .A3(n_266), .B(n_213), .Y(n_315) );
O2A1O1Ixp33_ASAP7_75t_L g316 ( .A1(n_308), .A2(n_246), .B(n_223), .C(n_236), .Y(n_316) );
A2O1A1Ixp33_ASAP7_75t_L g317 ( .A1(n_310), .A2(n_262), .B(n_211), .C(n_217), .Y(n_317) );
O2A1O1Ixp33_ASAP7_75t_SL g318 ( .A1(n_280), .A2(n_253), .B(n_261), .C(n_245), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_274), .Y(n_319) );
OAI22xp33_ASAP7_75t_L g320 ( .A1(n_270), .A2(n_221), .B1(n_236), .B2(n_261), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_SL g321 ( .A1(n_312), .A2(n_253), .B(n_251), .C(n_254), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_283), .Y(n_322) );
AO31x2_ASAP7_75t_L g323 ( .A1(n_295), .A2(n_260), .A3(n_262), .B(n_296), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_268), .Y(n_324) );
BUFx4_ASAP7_75t_SL g325 ( .A(n_314), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_273), .A2(n_269), .B1(n_298), .B2(n_311), .Y(n_326) );
OAI21xp5_ASAP7_75t_L g327 ( .A1(n_282), .A2(n_277), .B(n_307), .Y(n_327) );
OAI21x1_ASAP7_75t_L g328 ( .A1(n_290), .A2(n_303), .B(n_272), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_SL g329 ( .A1(n_306), .A2(n_301), .B(n_297), .C(n_286), .Y(n_329) );
INVx1_ASAP7_75t_SL g330 ( .A(n_287), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_279), .A2(n_300), .B(n_275), .Y(n_331) );
O2A1O1Ixp33_ASAP7_75t_L g332 ( .A1(n_281), .A2(n_278), .B(n_304), .C(n_284), .Y(n_332) );
O2A1O1Ixp33_ASAP7_75t_SL g333 ( .A1(n_285), .A2(n_292), .B(n_271), .C(n_313), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_289), .B(n_291), .Y(n_334) );
A2O1A1Ixp33_ASAP7_75t_L g335 ( .A1(n_299), .A2(n_305), .B(n_309), .C(n_293), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_302), .A2(n_274), .B(n_276), .Y(n_336) );
OAI21xp5_ASAP7_75t_L g337 ( .A1(n_302), .A2(n_288), .B(n_274), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_288), .A2(n_276), .B1(n_289), .B2(n_291), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_289), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_291), .B(n_276), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_L g341 ( .A1(n_288), .A2(n_263), .B(n_257), .C(n_308), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_302), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_288), .B(n_270), .Y(n_343) );
O2A1O1Ixp33_ASAP7_75t_L g344 ( .A1(n_308), .A2(n_263), .B(n_257), .C(n_229), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_328), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_344), .B(n_324), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_319), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_321), .A2(n_318), .B(n_327), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_319), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_341), .Y(n_350) );
AO31x2_ASAP7_75t_L g351 ( .A1(n_317), .A2(n_326), .A3(n_335), .B(n_331), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_343), .A2(n_320), .B1(n_338), .B2(n_332), .Y(n_352) );
AO31x2_ASAP7_75t_L g353 ( .A1(n_315), .A2(n_323), .A3(n_336), .B(n_340), .Y(n_353) );
CKINVDCx14_ASAP7_75t_R g354 ( .A(n_322), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_330), .B(n_343), .Y(n_355) );
NAND2x1p5_ASAP7_75t_L g356 ( .A(n_319), .B(n_334), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_325), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_316), .B(n_334), .Y(n_358) );
AO31x2_ASAP7_75t_L g359 ( .A1(n_315), .A2(n_323), .A3(n_329), .B(n_342), .Y(n_359) );
AOI22xp33_ASAP7_75t_SL g360 ( .A1(n_337), .A2(n_339), .B1(n_338), .B2(n_333), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_315), .Y(n_361) );
NOR2x1_ASAP7_75t_SL g362 ( .A(n_323), .B(n_265), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_344), .B(n_270), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_344), .B(n_270), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_344), .Y(n_365) );
OAI21x1_ASAP7_75t_L g366 ( .A1(n_328), .A2(n_296), .B(n_295), .Y(n_366) );
BUFx2_ASAP7_75t_L g367 ( .A(n_319), .Y(n_367) );
CKINVDCx20_ASAP7_75t_R g368 ( .A(n_322), .Y(n_368) );
BUFx3_ASAP7_75t_L g369 ( .A(n_319), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_344), .B(n_270), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_346), .B(n_365), .Y(n_371) );
INVx2_ASAP7_75t_SL g372 ( .A(n_369), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_346), .B(n_365), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_350), .B(n_369), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_345), .Y(n_375) );
OA21x2_ASAP7_75t_L g376 ( .A1(n_348), .A2(n_366), .B(n_345), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_366), .Y(n_377) );
BUFx2_ASAP7_75t_L g378 ( .A(n_361), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_364), .B(n_350), .Y(n_379) );
AO21x2_ASAP7_75t_L g380 ( .A1(n_362), .A2(n_370), .B(n_363), .Y(n_380) );
OAI22xp5_ASAP7_75t_SL g381 ( .A1(n_354), .A2(n_357), .B1(n_368), .B2(n_355), .Y(n_381) );
AO21x2_ASAP7_75t_L g382 ( .A1(n_362), .A2(n_358), .B(n_352), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_359), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_349), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_369), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_349), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_353), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_364), .B(n_351), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_353), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_353), .Y(n_390) );
OAI21xp5_ASAP7_75t_L g391 ( .A1(n_360), .A2(n_367), .B(n_356), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_359), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_351), .B(n_359), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_367), .A2(n_347), .B1(n_356), .B2(n_357), .Y(n_394) );
AOI21x1_ASAP7_75t_L g395 ( .A1(n_359), .A2(n_351), .B(n_353), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_353), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_359), .Y(n_397) );
INVx2_ASAP7_75t_SL g398 ( .A(n_347), .Y(n_398) );
OAI221xp5_ASAP7_75t_L g399 ( .A1(n_356), .A2(n_229), .B1(n_273), .B2(n_257), .C(n_263), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g400 ( .A1(n_347), .A2(n_344), .B(n_341), .Y(n_400) );
BUFx3_ASAP7_75t_L g401 ( .A(n_347), .Y(n_401) );
OA21x2_ASAP7_75t_L g402 ( .A1(n_351), .A2(n_348), .B(n_366), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_371), .B(n_351), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_371), .B(n_373), .Y(n_404) );
INVxp67_ASAP7_75t_SL g405 ( .A(n_375), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_371), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_378), .B(n_388), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_373), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_373), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_379), .Y(n_410) );
BUFx3_ASAP7_75t_L g411 ( .A(n_385), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_393), .B(n_388), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_375), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_375), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_379), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_399), .A2(n_378), .B1(n_379), .B2(n_374), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_387), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_393), .B(n_388), .Y(n_418) );
INVx4_ASAP7_75t_L g419 ( .A(n_385), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_393), .B(n_374), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_387), .Y(n_421) );
BUFx3_ASAP7_75t_L g422 ( .A(n_385), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_387), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_389), .Y(n_424) );
INVx3_ASAP7_75t_L g425 ( .A(n_376), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_377), .Y(n_426) );
OAI31xp33_ASAP7_75t_SL g427 ( .A1(n_399), .A2(n_391), .A3(n_400), .B(n_389), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_389), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_390), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_390), .B(n_396), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_378), .B(n_396), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_374), .B(n_397), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_383), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_384), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_374), .B(n_397), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_383), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_374), .B(n_392), .Y(n_437) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_376), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_374), .B(n_392), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_392), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_384), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_392), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_412), .B(n_402), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_404), .B(n_386), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_412), .B(n_402), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_432), .B(n_435), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_412), .B(n_402), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_404), .B(n_386), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_417), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_403), .B(n_402), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_417), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_403), .B(n_402), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_432), .B(n_402), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_434), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_421), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_426), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_406), .B(n_394), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_416), .A2(n_382), .B1(n_400), .B2(n_380), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_435), .B(n_395), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_407), .B(n_382), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_426), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_406), .B(n_394), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_408), .B(n_372), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_411), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_421), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_423), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_408), .B(n_372), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_409), .B(n_372), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_409), .B(n_381), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_410), .B(n_395), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_410), .B(n_385), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_415), .B(n_395), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_415), .B(n_382), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_423), .Y(n_474) );
INVx2_ASAP7_75t_SL g475 ( .A(n_411), .Y(n_475) );
NOR3xp33_ASAP7_75t_L g476 ( .A(n_431), .B(n_381), .C(n_391), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_418), .B(n_382), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_437), .B(n_382), .Y(n_478) );
INVx2_ASAP7_75t_SL g479 ( .A(n_411), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_434), .Y(n_480) );
INVx1_ASAP7_75t_SL g481 ( .A(n_422), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_424), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_424), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_418), .B(n_380), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_437), .B(n_380), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_439), .B(n_380), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_428), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_439), .B(n_380), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_407), .B(n_376), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_428), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_431), .B(n_376), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_420), .B(n_376), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_420), .B(n_401), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_430), .B(n_401), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_441), .B(n_398), .Y(n_495) );
INVxp67_ASAP7_75t_SL g496 ( .A(n_454), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_449), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_470), .B(n_430), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_449), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_451), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_451), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_470), .B(n_430), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_472), .B(n_429), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_455), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_455), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_444), .B(n_441), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_446), .B(n_419), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_446), .B(n_419), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_446), .B(n_419), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_448), .B(n_413), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_472), .B(n_429), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_446), .B(n_419), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_450), .B(n_427), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_465), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_480), .B(n_413), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_465), .Y(n_516) );
INVx1_ASAP7_75t_SL g517 ( .A(n_464), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_466), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_493), .B(n_422), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_493), .B(n_422), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_450), .B(n_427), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_443), .B(n_405), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_452), .B(n_436), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_466), .Y(n_524) );
NOR2x1p5_ASAP7_75t_L g525 ( .A(n_464), .B(n_425), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_474), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_456), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_443), .B(n_405), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_452), .B(n_436), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_445), .B(n_442), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_474), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_445), .B(n_442), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_494), .B(n_442), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_482), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_447), .B(n_440), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_494), .B(n_440), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_482), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_447), .B(n_414), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_489), .B(n_414), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_483), .Y(n_540) );
AND2x4_ASAP7_75t_SL g541 ( .A(n_475), .B(n_398), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_483), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_456), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_489), .B(n_414), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_529), .B(n_460), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_533), .B(n_459), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_529), .B(n_460), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_498), .B(n_484), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_513), .B(n_484), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_496), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_517), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_498), .B(n_491), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_513), .B(n_459), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_497), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_499), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_500), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_501), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_521), .B(n_477), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_517), .A2(n_469), .B1(n_476), .B2(n_479), .Y(n_559) );
INVxp67_ASAP7_75t_L g560 ( .A(n_521), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_536), .B(n_453), .Y(n_561) );
NOR2x1_ASAP7_75t_L g562 ( .A(n_525), .B(n_495), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_504), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_502), .B(n_477), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_502), .B(n_453), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_505), .Y(n_566) );
NOR2xp67_ASAP7_75t_SL g567 ( .A(n_507), .B(n_479), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_503), .B(n_473), .Y(n_568) );
INVxp67_ASAP7_75t_L g569 ( .A(n_515), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_503), .B(n_473), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_530), .B(n_478), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_514), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_530), .B(n_478), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_527), .Y(n_574) );
AOI221xp5_ASAP7_75t_L g575 ( .A1(n_511), .A2(n_458), .B1(n_462), .B2(n_457), .C(n_490), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_516), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_532), .B(n_478), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_511), .B(n_492), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_554), .Y(n_579) );
OAI21xp33_ASAP7_75t_L g580 ( .A1(n_560), .A2(n_523), .B(n_532), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_560), .B(n_506), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_555), .Y(n_582) );
AOI21xp33_ASAP7_75t_SL g583 ( .A1(n_559), .A2(n_508), .B(n_509), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_556), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_557), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_562), .A2(n_508), .B1(n_512), .B2(n_522), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_553), .B(n_535), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_563), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_549), .A2(n_558), .B1(n_575), .B2(n_551), .Y(n_589) );
OAI211xp5_ASAP7_75t_L g590 ( .A1(n_569), .A2(n_481), .B(n_475), .C(n_528), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_571), .B(n_520), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_566), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_571), .B(n_519), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_565), .B(n_535), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_565), .B(n_510), .Y(n_595) );
INVxp67_ASAP7_75t_SL g596 ( .A(n_574), .Y(n_596) );
OAI22xp33_ASAP7_75t_SL g597 ( .A1(n_569), .A2(n_538), .B1(n_544), .B2(n_539), .Y(n_597) );
AOI221xp5_ASAP7_75t_L g598 ( .A1(n_550), .A2(n_531), .B1(n_540), .B2(n_537), .C(n_534), .Y(n_598) );
O2A1O1Ixp33_ASAP7_75t_SL g599 ( .A1(n_552), .A2(n_491), .B(n_495), .C(n_471), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_579), .Y(n_600) );
AOI222xp33_ASAP7_75t_L g601 ( .A1(n_580), .A2(n_586), .B1(n_598), .B2(n_590), .C1(n_581), .C2(n_582), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_583), .B(n_577), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g603 ( .A1(n_589), .A2(n_567), .B1(n_545), .B2(n_547), .C(n_568), .Y(n_603) );
AOI221xp5_ASAP7_75t_L g604 ( .A1(n_597), .A2(n_573), .B1(n_577), .B2(n_564), .C(n_578), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_590), .A2(n_573), .B1(n_570), .B2(n_546), .Y(n_605) );
AOI322xp5_ASAP7_75t_L g606 ( .A1(n_594), .A2(n_546), .A3(n_561), .B1(n_576), .B2(n_572), .C1(n_485), .C2(n_488), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_587), .A2(n_548), .B1(n_561), .B2(n_541), .Y(n_607) );
OAI211xp5_ASAP7_75t_L g608 ( .A1(n_599), .A2(n_468), .B(n_467), .C(n_463), .Y(n_608) );
NOR2xp33_ASAP7_75t_SL g609 ( .A(n_596), .B(n_492), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_598), .A2(n_478), .B1(n_485), .B2(n_488), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_584), .Y(n_611) );
OAI21xp33_ASAP7_75t_L g612 ( .A1(n_595), .A2(n_574), .B(n_486), .Y(n_612) );
NAND2xp33_ASAP7_75t_SL g613 ( .A(n_602), .B(n_593), .Y(n_613) );
AOI21xp33_ASAP7_75t_SL g614 ( .A1(n_601), .A2(n_592), .B(n_588), .Y(n_614) );
OAI211xp5_ASAP7_75t_L g615 ( .A1(n_610), .A2(n_585), .B(n_591), .C(n_518), .Y(n_615) );
OAI211xp5_ASAP7_75t_L g616 ( .A1(n_603), .A2(n_524), .B(n_542), .C(n_526), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_600), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_607), .A2(n_486), .B1(n_490), .B2(n_487), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_604), .A2(n_487), .B1(n_543), .B2(n_425), .C(n_438), .Y(n_619) );
AOI211xp5_ASAP7_75t_L g620 ( .A1(n_614), .A2(n_608), .B(n_609), .C(n_612), .Y(n_620) );
OAI211xp5_ASAP7_75t_L g621 ( .A1(n_613), .A2(n_606), .B(n_605), .C(n_611), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_616), .B(n_425), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_617), .B(n_425), .Y(n_623) );
NOR3xp33_ASAP7_75t_L g624 ( .A(n_621), .B(n_615), .C(n_619), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_623), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_625), .Y(n_626) );
AND3x1_ASAP7_75t_L g627 ( .A(n_624), .B(n_620), .C(n_622), .Y(n_627) );
NOR2xp67_ASAP7_75t_L g628 ( .A(n_626), .B(n_618), .Y(n_628) );
INVx5_ASAP7_75t_L g629 ( .A(n_628), .Y(n_629) );
AOI21x1_ASAP7_75t_L g630 ( .A1(n_629), .A2(n_627), .B(n_461), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_630), .A2(n_629), .B1(n_401), .B2(n_438), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_631), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_632), .A2(n_438), .B1(n_440), .B2(n_433), .Y(n_633) );
endmodule