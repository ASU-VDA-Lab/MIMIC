module real_jpeg_25864_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_1),
.A2(n_55),
.B1(n_56),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_1),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_98),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_1),
.A2(n_27),
.B1(n_31),
.B2(n_98),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_2),
.A2(n_27),
.B1(n_31),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_2),
.A2(n_37),
.B1(n_55),
.B2(n_56),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_3),
.Y(n_94)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_6),
.A2(n_39),
.B1(n_40),
.B2(n_66),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_6),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_6),
.A2(n_66),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_6),
.A2(n_55),
.B1(n_56),
.B2(n_66),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_6),
.A2(n_27),
.B1(n_31),
.B2(n_66),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_7),
.A2(n_44),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_7),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_71),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_7),
.A2(n_55),
.B1(n_56),
.B2(n_71),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_7),
.A2(n_27),
.B1(n_31),
.B2(n_71),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_8),
.A2(n_27),
.B1(n_31),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_8),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_11),
.B(n_48),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_11),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_11),
.B(n_74),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_11),
.B(n_56),
.C(n_58),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_11),
.A2(n_39),
.B1(n_40),
.B2(n_110),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_11),
.B(n_67),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_11),
.A2(n_55),
.B1(n_56),
.B2(n_110),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_11),
.B(n_27),
.C(n_94),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_11),
.A2(n_26),
.B(n_201),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_13),
.A2(n_39),
.B1(n_40),
.B2(n_63),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_13),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_63),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_13),
.A2(n_55),
.B1(n_56),
.B2(n_63),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_13),
.A2(n_27),
.B1(n_31),
.B2(n_63),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_14),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_14),
.A2(n_32),
.B1(n_55),
.B2(n_56),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_15),
.A2(n_27),
.B1(n_31),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_15),
.Y(n_120)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_16),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_16),
.A2(n_25),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_139),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_138),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_113),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_21),
.B(n_113),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_82),
.C(n_100),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_22),
.B(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_23),
.B(n_52),
.C(n_68),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_38),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_24),
.B(n_38),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_33),
.B2(n_36),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_26),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_26),
.A2(n_85),
.B1(n_87),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_26),
.A2(n_30),
.B1(n_34),
.B2(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_26),
.B(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_26),
.A2(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_27),
.A2(n_31),
.B1(n_94),
.B2(n_95),
.Y(n_96)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_28),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_31),
.B(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_34),
.A2(n_214),
.B(n_222),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_36),
.Y(n_84)
);

AOI32xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.A3(n_45),
.B1(n_47),
.B2(n_50),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_40),
.B1(n_58),
.B2(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_39),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_74)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp33_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_46),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_40),
.B(n_164),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_43),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_81)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_47),
.Y(n_111)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_68),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_61),
.B(n_64),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_53),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_53),
.A2(n_64),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_60),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_54),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_54),
.A2(n_136),
.B(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_56),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_56),
.B(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_67),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_65),
.B(n_107),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_73),
.B(n_75),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_70),
.A2(n_74),
.B1(n_80),
.B2(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_77),
.Y(n_112)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_110),
.B(n_111),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_109),
.B(n_112),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_82),
.B(n_100),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_90),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_83),
.B(n_90),
.Y(n_137)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_89),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_89),
.B(n_110),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_96),
.B1(n_97),
.B2(n_99),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_91),
.A2(n_188),
.B(n_189),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_91),
.A2(n_189),
.B(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_92),
.A2(n_124),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_97),
.B(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_96),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_96),
.A2(n_103),
.B(n_174),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_96),
.B(n_110),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_99),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.C(n_108),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_101),
.A2(n_102),
.B1(n_105),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_104),
.B(n_124),
.Y(n_189)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_106),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_127),
.B2(n_128),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_121),
.B1(n_125),
.B2(n_126),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_118),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_137),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_243),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_158),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_156),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_143),
.B(n_156),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.C(n_149),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_144),
.A2(n_145),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_148),
.B(n_149),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_154),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_183),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_237),
.B(n_242),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_190),
.B(n_236),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_179),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_161),
.B(n_179),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_172),
.C(n_176),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_162),
.B(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_165),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B(n_170),
.Y(n_165)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_172),
.A2(n_176),
.B1(n_177),
.B2(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_172),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_175),
.Y(n_188)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_184),
.B2(n_185),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_180),
.B(n_186),
.C(n_187),
.Y(n_241)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_230),
.B(n_235),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_210),
.B(n_229),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_204),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_204),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_199),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_198),
.C(n_199),
.Y(n_234)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_200),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_208),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_218),
.B(n_228),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_216),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_216),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_223),
.B(n_227),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_221),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_234),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_241),
.Y(n_242)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);


endmodule