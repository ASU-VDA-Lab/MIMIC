module fake_jpeg_17004_n_292 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_292);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_292;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_20),
.B(n_7),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_41),
.Y(n_48)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g41 ( 
.A(n_25),
.B(n_0),
.CON(n_41),
.SN(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_29),
.Y(n_50)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_31),
.B1(n_33),
.B2(n_23),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_44),
.A2(n_49),
.B1(n_21),
.B2(n_24),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_31),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_63),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_31),
.B1(n_33),
.B2(n_23),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_51),
.B(n_18),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_0),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_17),
.B(n_23),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_33),
.B1(n_19),
.B2(n_26),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_40),
.B1(n_43),
.B2(n_38),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_38),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_64),
.B(n_72),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_65),
.B(n_95),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_67),
.A2(n_73),
.B1(n_87),
.B2(n_59),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_21),
.Y(n_107)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_43),
.B1(n_37),
.B2(n_38),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_74),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_17),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_77),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_17),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_0),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_83),
.B(n_19),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_37),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_32),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVxp33_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_46),
.A2(n_40),
.B1(n_19),
.B2(n_26),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_32),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_57),
.B1(n_59),
.B2(n_55),
.Y(n_108)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_26),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_53),
.B(n_30),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_44),
.Y(n_97)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

OA21x2_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_47),
.B(n_58),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_104),
.A2(n_107),
.B(n_118),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_35),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_68),
.C(n_69),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_108),
.A2(n_110),
.B1(n_57),
.B2(n_55),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_98),
.A2(n_30),
.B1(n_24),
.B2(n_22),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_70),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_117),
.Y(n_153)
);

NAND2x1_ASAP7_75t_SL g118 ( 
.A(n_84),
.B(n_27),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_66),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_125),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_66),
.B(n_61),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_77),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_127),
.B(n_135),
.C(n_139),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_101),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_145),
.Y(n_157)
);

OAI32xp33_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_76),
.A3(n_66),
.B1(n_87),
.B2(n_80),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_99),
.A3(n_104),
.B1(n_118),
.B2(n_123),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_126),
.A2(n_84),
.B1(n_80),
.B2(n_69),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_131),
.A2(n_116),
.B(n_27),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_70),
.Y(n_132)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_134),
.A2(n_156),
.B(n_122),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_78),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_78),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_138),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_42),
.C(n_56),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

AO22x1_ASAP7_75t_L g141 ( 
.A1(n_104),
.A2(n_71),
.B1(n_54),
.B2(n_61),
.Y(n_141)
);

AO22x1_ASAP7_75t_L g177 ( 
.A1(n_141),
.A2(n_59),
.B1(n_54),
.B2(n_116),
.Y(n_177)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_79),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_143),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_42),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_99),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_124),
.B(n_86),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_75),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_96),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_154),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_155),
.B1(n_54),
.B2(n_120),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_101),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_114),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_93),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_57),
.B1(n_90),
.B2(n_92),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_42),
.B(n_27),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_158),
.B(n_19),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_160),
.C(n_127),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_107),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_123),
.B(n_118),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_161),
.A2(n_170),
.B(n_171),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_153),
.A2(n_117),
.B1(n_107),
.B2(n_106),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_167),
.B1(n_174),
.B2(n_180),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_106),
.B1(n_90),
.B2(n_115),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_124),
.Y(n_168)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_122),
.Y(n_170)
);

AOI221xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_147),
.B1(n_129),
.B2(n_151),
.C(n_34),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_134),
.A2(n_139),
.B1(n_130),
.B2(n_141),
.Y(n_174)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_182),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_177),
.A2(n_155),
.B(n_152),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_26),
.Y(n_178)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_147),
.B1(n_156),
.B2(n_154),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_148),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_137),
.B1(n_85),
.B2(n_56),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_189),
.A2(n_194),
.B(n_177),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_195),
.C(n_200),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_42),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_170),
.A2(n_142),
.B1(n_140),
.B2(n_133),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_196),
.A2(n_205),
.B1(n_22),
.B2(n_29),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_186),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_209),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_163),
.B(n_168),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_198),
.B(n_199),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_164),
.B(n_133),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_128),
.C(n_137),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_202),
.A2(n_178),
.B(n_158),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_203),
.Y(n_216)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_85),
.B1(n_2),
.B2(n_3),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_34),
.C(n_28),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_208),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_157),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_34),
.C(n_28),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_210),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_187),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_223),
.B1(n_230),
.B2(n_22),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_186),
.Y(n_214)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_208),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_217),
.B(n_227),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_192),
.B(n_173),
.Y(n_219)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_191),
.A2(n_184),
.B1(n_172),
.B2(n_162),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_193),
.B(n_167),
.Y(n_221)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

A2O1A1Ixp33_ASAP7_75t_SL g224 ( 
.A1(n_191),
.A2(n_180),
.B(n_174),
.C(n_171),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_224),
.A2(n_226),
.B(n_196),
.Y(n_243)
);

AOI322xp5_ASAP7_75t_L g227 ( 
.A1(n_188),
.A2(n_160),
.A3(n_177),
.B1(n_181),
.B2(n_179),
.C1(n_22),
.C2(n_28),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_188),
.A2(n_181),
.B(n_179),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_228),
.A2(n_189),
.B(n_205),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_229),
.B(n_195),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_242),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_243),
.B(n_221),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_201),
.Y(n_233)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_216),
.A2(n_206),
.B1(n_202),
.B2(n_200),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_219),
.B1(n_224),
.B2(n_212),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_220),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_237),
.A2(n_224),
.B1(n_222),
.B2(n_225),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_190),
.C(n_207),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_244),
.C(n_245),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_228),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_206),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_203),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_246),
.A2(n_225),
.B1(n_213),
.B2(n_222),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_238),
.A2(n_224),
.B1(n_211),
.B2(n_213),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_247),
.A2(n_259),
.B1(n_1),
.B2(n_2),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_258),
.C(n_231),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

NAND4xp25_ASAP7_75t_SL g269 ( 
.A(n_250),
.B(n_9),
.C(n_14),
.D(n_5),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_253),
.B(n_1),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_226),
.B(n_214),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_9),
.B(n_14),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_243),
.A2(n_215),
.B(n_218),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_257),
.A2(n_237),
.B(n_245),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_215),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_238),
.A2(n_230),
.B1(n_9),
.B2(n_10),
.Y(n_259)
);

OAI221xp5_ASAP7_75t_L g260 ( 
.A1(n_255),
.A2(n_235),
.B1(n_236),
.B2(n_239),
.C(n_242),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_260),
.B(n_261),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_264),
.C(n_265),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_11),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_251),
.A2(n_8),
.B(n_14),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_269),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_270),
.C(n_259),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_254),
.A2(n_10),
.B(n_13),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_249),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_274),
.C(n_271),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_252),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_275),
.A2(n_276),
.B(n_277),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_252),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_254),
.Y(n_280)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_280),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_278),
.A2(n_256),
.B(n_10),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_281),
.A2(n_284),
.B(n_7),
.Y(n_288)
);

AO21x1_ASAP7_75t_L g287 ( 
.A1(n_282),
.A2(n_7),
.B(n_12),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_8),
.C(n_13),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_283),
.A2(n_279),
.B(n_6),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_278),
.A2(n_11),
.B(n_13),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_287),
.C(n_288),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_12),
.C(n_29),
.Y(n_290)
);

AO21x1_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_12),
.B(n_4),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_289),
.B1(n_3),
.B2(n_29),
.Y(n_292)
);


endmodule