module fake_netlist_6_763_n_252 (n_41, n_16, n_45, n_1, n_46, n_34, n_42, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_27, n_3, n_14, n_38, n_0, n_39, n_32, n_4, n_36, n_22, n_26, n_13, n_35, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_43, n_5, n_19, n_47, n_48, n_29, n_31, n_25, n_40, n_44, n_252);

input n_41;
input n_16;
input n_45;
input n_1;
input n_46;
input n_34;
input n_42;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_39;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_43;
input n_5;
input n_19;
input n_47;
input n_48;
input n_29;
input n_31;
input n_25;
input n_40;
input n_44;

output n_252;

wire n_52;
wire n_91;
wire n_119;
wire n_163;
wire n_146;
wire n_235;
wire n_193;
wire n_147;
wire n_191;
wire n_154;
wire n_88;
wire n_209;
wire n_98;
wire n_113;
wire n_63;
wire n_223;
wire n_73;
wire n_148;
wire n_199;
wire n_138;
wire n_161;
wire n_208;
wire n_68;
wire n_226;
wire n_228;
wire n_166;
wire n_184;
wire n_212;
wire n_50;
wire n_158;
wire n_49;
wire n_210;
wire n_217;
wire n_83;
wire n_216;
wire n_206;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_153;
wire n_168;
wire n_215;
wire n_125;
wire n_178;
wire n_247;
wire n_225;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_227;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_204;
wire n_245;
wire n_87;
wire n_195;
wire n_189;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_213;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_197;
wire n_137;
wire n_203;
wire n_142;
wire n_143;
wire n_207;
wire n_242;
wire n_180;
wire n_155;
wire n_62;
wire n_219;
wire n_75;
wire n_109;
wire n_150;
wire n_233;
wire n_122;
wire n_205;
wire n_140;
wire n_218;
wire n_70;
wire n_120;
wire n_234;
wire n_251;
wire n_214;
wire n_67;
wire n_82;
wire n_236;
wire n_246;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_237;
wire n_81;
wire n_59;
wire n_244;
wire n_181;
wire n_76;
wire n_182;
wire n_238;
wire n_124;
wire n_239;
wire n_55;
wire n_126;
wire n_202;
wire n_94;
wire n_108;
wire n_97;
wire n_58;
wire n_116;
wire n_211;
wire n_64;
wire n_220;
wire n_117;
wire n_118;
wire n_175;
wire n_224;
wire n_231;
wire n_65;
wire n_230;
wire n_93;
wire n_80;
wire n_141;
wire n_240;
wire n_135;
wire n_200;
wire n_196;
wire n_165;
wire n_139;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_222;
wire n_95;
wire n_179;
wire n_243;
wire n_248;
wire n_107;
wire n_71;
wire n_74;
wire n_229;
wire n_190;
wire n_123;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_249;
wire n_173;
wire n_201;
wire n_250;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_183;
wire n_232;
wire n_115;
wire n_69;
wire n_128;
wire n_241;
wire n_79;
wire n_194;
wire n_171;
wire n_192;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_56;
wire n_221;

INVx1_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

INVxp33_ASAP7_75t_SL g54 ( 
.A(n_41),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVxp33_ASAP7_75t_SL g56 ( 
.A(n_21),
.Y(n_56)
);

INVxp67_ASAP7_75t_SL g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_7),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_18),
.B(n_12),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_4),
.Y(n_70)
);

INVxp33_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_6),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_7),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_8),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_0),
.Y(n_87)
);

AND2x4_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_19),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_1),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

AND2x4_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_23),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_2),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_54),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

OA21x2_ASAP7_75t_L g98 ( 
.A1(n_67),
.A2(n_3),
.B(n_5),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_3),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_70),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_5),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_56),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_54),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_70),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_56),
.B1(n_53),
.B2(n_62),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_93),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_94),
.B(n_69),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_25),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_27),
.Y(n_120)
);

AND2x4_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_24),
.Y(n_121)
);

AND2x4_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_93),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_28),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_17),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_87),
.B(n_72),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

OR2x6_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_91),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_99),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_90),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_90),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_92),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_112),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

OR2x6_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_126),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_114),
.Y(n_147)
);

OR2x6_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_126),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_135),
.B(n_106),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_123),
.B(n_120),
.C(n_110),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

AND2x4_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_79),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_117),
.Y(n_155)
);

AND2x4_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_133),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_80),
.B1(n_89),
.B2(n_100),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_143),
.A2(n_128),
.B(n_131),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_138),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_144),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_129),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_124),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

AND2x4_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_141),
.Y(n_167)
);

AO21x2_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_119),
.B(n_95),
.Y(n_168)
);

AOI21x1_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_127),
.B(n_141),
.Y(n_169)
);

CKINVDCx11_ASAP7_75t_R g170 ( 
.A(n_161),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_132),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

OAI21x1_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_98),
.B(n_92),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_103),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_153),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_155),
.Y(n_184)
);

OA21x2_ASAP7_75t_L g185 ( 
.A1(n_175),
.A2(n_165),
.B(n_147),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_164),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_162),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_148),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_148),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_146),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_183),
.A2(n_146),
.B1(n_112),
.B2(n_157),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

OAI33xp33_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_157),
.A3(n_149),
.B1(n_171),
.B2(n_144),
.B3(n_179),
.Y(n_201)
);

AO21x2_ASAP7_75t_L g202 ( 
.A1(n_192),
.A2(n_168),
.B(n_175),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

AOI221xp5_ASAP7_75t_L g204 ( 
.A1(n_198),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.C(n_97),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

OA21x2_ASAP7_75t_L g206 ( 
.A1(n_193),
.A2(n_169),
.B(n_173),
.Y(n_206)
);

INVxp67_ASAP7_75t_SL g207 ( 
.A(n_189),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_199),
.Y(n_208)
);

AO21x2_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_168),
.B(n_169),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_146),
.Y(n_210)
);

INVxp67_ASAP7_75t_SL g211 ( 
.A(n_189),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_210),
.A2(n_188),
.B1(n_190),
.B2(n_187),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_208),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_190),
.Y(n_216)
);

OR2x6_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_197),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_207),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_202),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_202),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_213),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_202),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_223),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_216),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_219),
.A2(n_204),
.B1(n_208),
.B2(n_195),
.Y(n_228)
);

NAND2x1p5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_205),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_209),
.Y(n_230)
);

NOR3x1_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_224),
.C(n_221),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_222),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_226),
.Y(n_233)
);

NOR3x1_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_125),
.C(n_183),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_233),
.B(n_222),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_231),
.Y(n_236)
);

INVxp67_ASAP7_75t_SL g237 ( 
.A(n_236),
.Y(n_237)
);

NOR4xp25_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_232),
.C(n_204),
.D(n_234),
.Y(n_238)
);

OAI31xp33_ASAP7_75t_SL g239 ( 
.A1(n_236),
.A2(n_6),
.A3(n_8),
.B(n_9),
.Y(n_239)
);

AOI221xp5_ASAP7_75t_L g240 ( 
.A1(n_238),
.A2(n_101),
.B1(n_10),
.B2(n_229),
.C(n_167),
.Y(n_240)
);

OAI211xp5_ASAP7_75t_L g241 ( 
.A1(n_239),
.A2(n_98),
.B(n_101),
.C(n_196),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_98),
.B1(n_167),
.B2(n_203),
.Y(n_242)
);

NOR4xp25_ASAP7_75t_SL g243 ( 
.A(n_240),
.B(n_15),
.C(n_30),
.D(n_31),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_32),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_36),
.Y(n_245)
);

OAI211xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_205),
.B(n_145),
.C(n_185),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_242),
.Y(n_247)
);

NOR3xp33_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_244),
.C(n_246),
.Y(n_248)
);

AOI221xp5_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_145),
.B1(n_154),
.B2(n_46),
.C(n_47),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_185),
.B1(n_206),
.B2(n_145),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_248),
.Y(n_251)
);

AOI221xp5_ASAP7_75t_L g252 ( 
.A1(n_251),
.A2(n_250),
.B1(n_249),
.B2(n_154),
.C(n_111),
.Y(n_252)
);


endmodule