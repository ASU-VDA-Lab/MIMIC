module real_jpeg_32415_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_324;
wire n_86;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_0),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_1),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_1),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_1),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_1),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g206 ( 
.A(n_1),
.B(n_207),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_1),
.B(n_246),
.Y(n_245)
);

AND2x2_ASAP7_75t_SL g309 ( 
.A(n_1),
.B(n_209),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_1),
.B(n_343),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_3),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_3),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_3),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_3),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_3),
.B(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_4),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_4),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_5),
.B(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_5),
.B(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_5),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_5),
.B(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_6),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_6),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_7),
.Y(n_78)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_7),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_8),
.B(n_35),
.Y(n_34)
);

AND2x4_ASAP7_75t_L g164 ( 
.A(n_8),
.B(n_165),
.Y(n_164)
);

NAND2x1_ASAP7_75t_L g190 ( 
.A(n_8),
.B(n_191),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_8),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_8),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_8),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_8),
.B(n_377),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_8),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_9),
.B(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_9),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_9),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_9),
.B(n_94),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_9),
.B(n_275),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_9),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_9),
.B(n_357),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_9),
.B(n_170),
.Y(n_386)
);

AOI21xp33_ASAP7_75t_SL g18 ( 
.A1(n_10),
.A2(n_19),
.B(n_20),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_11),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_11),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_12),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_13),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_13),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_13),
.B(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_14),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_15),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_15),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_35),
.Y(n_43)
);

AND2x4_ASAP7_75t_SL g57 ( 
.A(n_16),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_16),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_16),
.B(n_77),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_16),
.B(n_100),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_16),
.B(n_258),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_16),
.B(n_261),
.Y(n_260)
);

AND2x2_ASAP7_75t_SL g292 ( 
.A(n_16),
.B(n_293),
.Y(n_292)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_17),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_17),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_17),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_17),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_17),
.B(n_221),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_325),
.B(n_430),
.C(n_441),
.Y(n_21)
);

INVxp33_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

O2A1O1Ixp33_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_224),
.B(n_277),
.C(n_324),
.Y(n_23)
);

AOI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_177),
.B(n_223),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_132),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_71),
.C(n_107),
.Y(n_26)
);

XOR2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_55),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_37),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_29),
.B(n_55),
.C(n_176),
.Y(n_175)
);

OA21x2_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_34),
.B(n_36),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_34),
.Y(n_36)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_32),
.Y(n_305)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_36),
.B(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_36),
.B(n_161),
.C(n_163),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_37),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_44),
.C(n_51),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_39),
.A2(n_219),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_40),
.A2(n_102),
.B1(n_105),
.B2(n_106),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_40),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_40),
.B(n_106),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_40),
.A2(n_105),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_40),
.B(n_43),
.Y(n_266)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_42),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_43),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_43),
.A2(n_256),
.B(n_263),
.Y(n_255)
);

OAI221xp5_ASAP7_75t_L g263 ( 
.A1(n_43),
.A2(n_257),
.B1(n_259),
.B2(n_260),
.C(n_262),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g289 ( 
.A(n_43),
.B(n_257),
.C(n_259),
.Y(n_289)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_50),
.Y(n_142)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_53),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_54),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_54),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_56),
.B(n_65),
.C(n_69),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_56),
.A2(n_57),
.B1(n_80),
.B2(n_359),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_56),
.A2(n_57),
.B1(n_153),
.B2(n_154),
.Y(n_384)
);

MAJx2_ASAP7_75t_L g387 ( 
.A(n_56),
.B(n_80),
.C(n_356),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_56),
.B(n_154),
.C(n_385),
.Y(n_409)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_65),
.B1(n_69),
.B2(n_70),
.Y(n_60)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_61),
.A2(n_69),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_68),
.Y(n_221)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_68),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_69),
.B(n_311),
.C(n_312),
.Y(n_310)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

MAJx2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_87),
.C(n_101),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_82),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_80),
.Y(n_74)
);

MAJx2_ASAP7_75t_L g130 ( 
.A(n_75),
.B(n_80),
.C(n_82),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_78),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_78),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_80),
.B(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_80),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_80),
.B(n_259),
.C(n_303),
.Y(n_362)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_93),
.C(n_97),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_126),
.B2(n_131),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_127),
.C(n_130),
.Y(n_134)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_114),
.Y(n_109)
);

MAJx2_ASAP7_75t_L g161 ( 
.A(n_110),
.B(n_116),
.C(n_120),
.Y(n_161)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_113),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_120),
.B2(n_121),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_124),
.Y(n_357)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_159),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_133),
.B(n_160),
.C(n_175),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_136),
.C(n_148),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_148),
.Y(n_135)
);

XNOR2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_147),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_143),
.Y(n_137)
);

NOR2xp67_ASAP7_75t_SL g185 ( 
.A(n_138),
.B(n_143),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_138),
.B(n_143),
.Y(n_186)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_185),
.B(n_186),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g215 ( 
.A(n_149),
.B(n_153),
.C(n_155),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_149),
.A2(n_150),
.B1(n_316),
.B2(n_320),
.Y(n_315)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_150),
.B(n_309),
.C(n_320),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

OA22x2_ASAP7_75t_L g410 ( 
.A1(n_153),
.A2(n_154),
.B1(n_411),
.B2(n_412),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_153),
.B(n_194),
.C(n_309),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_175),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_168),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_169),
.C(n_172),
.Y(n_197)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_222),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_178),
.B(n_222),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_200),
.B2(n_201),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_199),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_184),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_197),
.B2(n_198),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_190),
.Y(n_196)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g251 ( 
.A(n_194),
.B(n_196),
.C(n_198),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_194),
.A2(n_195),
.B1(n_308),
.B2(n_309),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_194),
.A2(n_195),
.B1(n_257),
.B2(n_262),
.Y(n_427)
);

NOR3xp33_ASAP7_75t_L g442 ( 
.A(n_194),
.B(n_262),
.C(n_342),
.Y(n_442)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_197),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_199),
.Y(n_233)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_214),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_239),
.C(n_240),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_208),
.C(n_212),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_208),
.B1(n_212),
.B2(n_213),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_206),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_206),
.A2(n_212),
.B1(n_336),
.B2(n_341),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_206),
.B(n_341),
.C(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_208),
.Y(n_213)
);

INVx4_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_215),
.Y(n_240)
);

INVxp67_ASAP7_75t_SL g239 ( 
.A(n_216),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NOR2xp67_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_231),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_225),
.A2(n_231),
.B1(n_278),
.B2(n_321),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.C(n_230),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_236),
.Y(n_231)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_232),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.C(n_235),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_254),
.Y(n_236)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_237),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_238),
.B(n_253),
.C(n_280),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_241)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_242),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_250),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_248),
.B2(n_249),
.Y(n_243)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_244),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_244),
.B(n_248),
.C(n_250),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_245),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_245),
.A2(n_248),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_245),
.A2(n_248),
.B1(n_375),
.B2(n_376),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_245),
.B(n_375),
.C(n_380),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_247),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_248),
.B(n_289),
.C(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_251),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_254),
.B(n_322),
.C(n_323),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_264),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_265),
.C(n_267),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_259),
.B1(n_260),
.B2(n_262),
.Y(n_256)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_257),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_259),
.A2(n_260),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_274),
.Y(n_269)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_270),
.Y(n_312)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_274),
.Y(n_311)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NOR2x1_ASAP7_75t_SL g324 ( 
.A(n_278),
.B(n_321),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_282),
.Y(n_278)
);

INVxp33_ASAP7_75t_SL g392 ( 
.A(n_279),
.Y(n_392)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_298),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_283),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

INVxp33_ASAP7_75t_SL g364 ( 
.A(n_284),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_297),
.Y(n_285)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_286),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_287),
.Y(n_365)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_292),
.Y(n_348)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_297),
.B(n_364),
.C(n_365),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_298),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_306),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

MAJx2_ASAP7_75t_L g351 ( 
.A(n_300),
.B(n_352),
.C(n_353),
.Y(n_351)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_314),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_313),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_308),
.A2(n_309),
.B1(n_314),
.B2(n_315),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_310),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_310),
.Y(n_353)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NOR3xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_396),
.C(n_421),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_388),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

OA21x2_ASAP7_75t_SL g433 ( 
.A1(n_328),
.A2(n_434),
.B(n_435),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_366),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_330),
.B(n_436),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_354),
.C(n_363),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_332),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_332),
.B(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_351),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_334),
.A2(n_347),
.B1(n_349),
.B2(n_350),
.Y(n_333)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_334),
.Y(n_349)
);

XOR2x2_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_342),
.Y(n_334)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_336),
.Y(n_341)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_342),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_342),
.B(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_345),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_346),
.Y(n_408)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_347),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_348),
.B(n_439),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_348),
.B(n_442),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_349),
.B(n_350),
.C(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_351),
.Y(n_368)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_354),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_360),
.Y(n_354)
);

MAJx2_ASAP7_75t_L g370 ( 
.A(n_355),
.B(n_361),
.C(n_362),
.Y(n_370)
);

XOR2x2_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_358),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_363),
.B(n_394),
.Y(n_393)
);

INVxp33_ASAP7_75t_SL g436 ( 
.A(n_366),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_369),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_367),
.B(n_419),
.C(n_420),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

INVxp33_ASAP7_75t_SL g419 ( 
.A(n_370),
.Y(n_419)
);

INVxp33_ASAP7_75t_SL g420 ( 
.A(n_371),
.Y(n_420)
);

XOR2x2_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_381),
.Y(n_371)
);

MAJx2_ASAP7_75t_L g416 ( 
.A(n_372),
.B(n_382),
.C(n_417),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_373),
.A2(n_374),
.B1(n_378),
.B2(n_380),
.Y(n_372)
);

INVxp33_ASAP7_75t_SL g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_378),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_387),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_383),
.A2(n_384),
.B1(n_385),
.B2(n_386),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_386),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_387),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_393),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_389),
.B(n_393),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.C(n_392),
.Y(n_389)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

OAI21xp33_ASAP7_75t_L g437 ( 
.A1(n_397),
.A2(n_422),
.B(n_432),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_418),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_398),
.B(n_418),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_415),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_401),
.B1(n_413),
.B2(n_414),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_400),
.B(n_413),
.C(n_416),
.Y(n_429)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

XNOR2x1_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_410),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_409),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_403),
.B(n_409),
.C(n_410),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx6_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_411),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_413),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_429),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_423),
.B(n_429),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_428),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_425),
.B(n_440),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_L g430 ( 
.A1(n_431),
.A2(n_433),
.B(n_437),
.C(n_438),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);


endmodule