module fake_jpeg_29472_n_530 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_530);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_530;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx5p33_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_15),
.B(n_4),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_51),
.B(n_15),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_55),
.B(n_59),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_56),
.A2(n_19),
.B1(n_26),
.B2(n_44),
.Y(n_154)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_14),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_16),
.B(n_25),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_61),
.B(n_65),
.Y(n_130)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_62),
.B(n_70),
.Y(n_111)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_63),
.Y(n_166)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_25),
.B(n_10),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_27),
.B(n_9),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_71),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_72),
.Y(n_169)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_76),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_78),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_27),
.B(n_9),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_79),
.B(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_84),
.Y(n_171)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_99),
.Y(n_125)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_87),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_16),
.B(n_8),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_95),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

INVxp67_ASAP7_75t_SL g98 ( 
.A(n_54),
.Y(n_98)
);

INVx5_ASAP7_75t_SL g164 ( 
.A(n_98),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_28),
.B(n_32),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_16),
.B(n_0),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_40),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_103),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_43),
.Y(n_105)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_28),
.B(n_0),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_106),
.B(n_19),
.Y(n_114)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_114),
.B(n_131),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_61),
.A2(n_32),
.B1(n_35),
.B2(n_39),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_117),
.A2(n_153),
.B1(n_154),
.B2(n_173),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_126),
.B(n_141),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_70),
.B(n_39),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_37),
.Y(n_134)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_42),
.Y(n_140)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_140),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_98),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_67),
.A2(n_40),
.B1(n_33),
.B2(n_50),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_146),
.A2(n_172),
.B1(n_54),
.B2(n_20),
.Y(n_177)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_57),
.Y(n_149)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_58),
.A2(n_21),
.B1(n_33),
.B2(n_26),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_67),
.B(n_48),
.Y(n_155)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_155),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_71),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_161),
.Y(n_224)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_162),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_56),
.A2(n_50),
.B(n_49),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_170),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_77),
.A2(n_91),
.B1(n_49),
.B2(n_50),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_69),
.A2(n_21),
.B1(n_26),
.B2(n_20),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_31),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_175),
.B(n_189),
.Y(n_228)
);

NAND2x1_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_21),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_176),
.B(n_219),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_177),
.A2(n_133),
.B1(n_159),
.B2(n_31),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_125),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_179),
.B(n_185),
.Y(n_229)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_110),
.Y(n_180)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_115),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_182),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_142),
.A2(n_87),
.B1(n_74),
.B2(n_101),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_183),
.A2(n_184),
.B1(n_221),
.B2(n_160),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_142),
.A2(n_88),
.B1(n_76),
.B2(n_96),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_137),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_164),
.A2(n_38),
.B1(n_89),
.B2(n_104),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_186),
.A2(n_208),
.B1(n_215),
.B2(n_216),
.Y(n_236)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_187),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_188),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_130),
.B(n_17),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_157),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_199),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_17),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_191),
.B(n_214),
.Y(n_244)
);

O2A1O1Ixp33_ASAP7_75t_SL g192 ( 
.A1(n_111),
.A2(n_21),
.B(n_54),
.C(n_89),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_192),
.A2(n_167),
.B1(n_160),
.B2(n_148),
.Y(n_262)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_194),
.Y(n_263)
);

OA22x2_ASAP7_75t_SL g195 ( 
.A1(n_151),
.A2(n_54),
.B1(n_21),
.B2(n_109),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_195),
.Y(n_259)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_136),
.Y(n_197)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_197),
.Y(n_264)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_144),
.Y(n_198)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_198),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_121),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_200),
.Y(n_227)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_115),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_202),
.Y(n_245)
);

INVx11_ASAP7_75t_L g203 ( 
.A(n_145),
.Y(n_203)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_203),
.Y(n_252)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_116),
.Y(n_204)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_204),
.Y(n_261)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_124),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_210),
.Y(n_239)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_207),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_164),
.A2(n_38),
.B1(n_48),
.B2(n_44),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_138),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_212),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_128),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_118),
.B(n_141),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_145),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_168),
.A2(n_42),
.B1(n_37),
.B2(n_35),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_158),
.B(n_53),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_159),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_171),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_218),
.B(n_161),
.Y(n_233)
);

AND2x2_ASAP7_75t_SL g219 ( 
.A(n_124),
.B(n_1),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_158),
.A2(n_95),
.B1(n_81),
.B2(n_78),
.Y(n_221)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_150),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_223),
.Y(n_242)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_127),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_225),
.Y(n_237)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_127),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_226),
.A2(n_120),
.B1(n_169),
.B2(n_129),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_233),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_234),
.Y(n_271)
);

AND2x6_ASAP7_75t_L g235 ( 
.A(n_174),
.B(n_172),
.Y(n_235)
);

A2O1A1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_235),
.A2(n_217),
.B(n_195),
.C(n_193),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_238),
.Y(n_279)
);

AOI22x1_ASAP7_75t_SL g241 ( 
.A1(n_176),
.A2(n_173),
.B1(n_153),
.B2(n_163),
.Y(n_241)
);

OAI21xp33_ASAP7_75t_SL g281 ( 
.A1(n_241),
.A2(n_165),
.B(n_201),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_247),
.A2(n_262),
.B1(n_224),
.B2(n_200),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_214),
.B(n_18),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_248),
.B(n_249),
.Y(n_275)
);

AOI21xp33_ASAP7_75t_L g249 ( 
.A1(n_189),
.A2(n_53),
.B(n_34),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_206),
.A2(n_166),
.B1(n_133),
.B2(n_120),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_250),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_191),
.A2(n_34),
.B(n_18),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_253),
.A2(n_220),
.B(n_178),
.Y(n_280)
);

INVx2_ASAP7_75t_R g254 ( 
.A(n_209),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_254),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_255),
.B(n_258),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_175),
.B(n_132),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_232),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_266),
.B(n_278),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_213),
.B1(n_195),
.B2(n_167),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_267),
.A2(n_269),
.B1(n_276),
.B2(n_284),
.Y(n_304)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_265),
.Y(n_268)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_213),
.B1(n_192),
.B2(n_209),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_270),
.A2(n_280),
.B(n_297),
.Y(n_313)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_264),
.Y(n_273)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_273),
.Y(n_305)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_240),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_274),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_241),
.A2(n_209),
.B1(n_219),
.B2(n_180),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_277),
.A2(n_281),
.B1(n_293),
.B2(n_295),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_232),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_222),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_248),
.C(n_258),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_254),
.A2(n_219),
.B1(n_181),
.B2(n_196),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_260),
.A2(n_187),
.B1(n_194),
.B2(n_113),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_229),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_285),
.B(n_287),
.Y(n_319)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_240),
.Y(n_286)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_229),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_260),
.A2(n_113),
.B1(n_223),
.B2(n_207),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_290),
.A2(n_256),
.B1(n_227),
.B2(n_237),
.Y(n_322)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_264),
.Y(n_291)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_291),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_260),
.A2(n_224),
.B(n_163),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_292),
.Y(n_323)
);

OAI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_235),
.A2(n_203),
.B1(n_225),
.B2(n_205),
.Y(n_293)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_244),
.B(n_143),
.C(n_119),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_294),
.B(n_276),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_255),
.A2(n_148),
.B1(n_215),
.B2(n_188),
.Y(n_295)
);

OAI21xp33_ASAP7_75t_SL g297 ( 
.A1(n_254),
.A2(n_226),
.B(n_204),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_228),
.B(n_197),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_228),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_273),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_299),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_307),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_266),
.B(n_253),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_308),
.B(n_325),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_269),
.A2(n_235),
.B1(n_236),
.B2(n_262),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_309),
.A2(n_322),
.B1(n_297),
.B2(n_304),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_233),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_310),
.B(n_315),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_281),
.A2(n_247),
.B1(n_239),
.B2(n_251),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_314),
.A2(n_328),
.B1(n_267),
.B2(n_290),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_239),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_291),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_316),
.Y(n_338)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_295),
.Y(n_317)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_317),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_288),
.B(n_251),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_321),
.Y(n_346)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_268),
.Y(n_320)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_320),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_288),
.B(n_242),
.Y(n_321)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_298),
.Y(n_326)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_326),
.Y(n_343)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_284),
.Y(n_327)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_327),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_277),
.A2(n_231),
.B1(n_227),
.B2(n_242),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_329),
.A2(n_341),
.B1(n_314),
.B2(n_328),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_313),
.A2(n_279),
.B(n_309),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_330),
.A2(n_320),
.B(n_311),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_334),
.A2(n_327),
.B1(n_322),
.B2(n_313),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_294),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_335),
.B(n_348),
.Y(n_359)
);

AO22x1_ASAP7_75t_SL g337 ( 
.A1(n_317),
.A2(n_293),
.B1(n_270),
.B2(n_294),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_337),
.B(n_301),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_302),
.B(n_282),
.C(n_292),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_353),
.C(n_357),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_304),
.A2(n_271),
.B1(n_289),
.B2(n_270),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_307),
.B(n_287),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_342),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_312),
.B(n_285),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_345),
.B(n_358),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_315),
.B(n_283),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_323),
.A2(n_296),
.B(n_289),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_349),
.A2(n_356),
.B(n_331),
.Y(n_369)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_321),
.Y(n_350)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_350),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_301),
.A2(n_278),
.B1(n_275),
.B2(n_280),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_351),
.A2(n_265),
.B1(n_257),
.B2(n_252),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_306),
.A2(n_307),
.B(n_312),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_352),
.A2(n_354),
.B(n_265),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_310),
.B(n_296),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_319),
.A2(n_275),
.B(n_245),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_324),
.Y(n_355)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_355),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_318),
.A2(n_261),
.B(n_245),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_261),
.C(n_237),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_319),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_358),
.B(n_299),
.Y(n_361)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_361),
.Y(n_392)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_346),
.Y(n_363)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_363),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_364),
.B(n_382),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_331),
.Y(n_365)
);

INVx13_ASAP7_75t_L g400 ( 
.A(n_365),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_344),
.B(n_316),
.Y(n_366)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_366),
.Y(n_399)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_346),
.Y(n_368)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_368),
.Y(n_417)
);

A2O1A1Ixp33_ASAP7_75t_SL g408 ( 
.A1(n_369),
.A2(n_337),
.B(n_340),
.C(n_355),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_370),
.A2(n_348),
.B1(n_347),
.B2(n_336),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_371),
.A2(n_372),
.B1(n_375),
.B2(n_381),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_334),
.A2(n_311),
.B1(n_305),
.B2(n_303),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_344),
.B(n_308),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_373),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_374),
.B(n_383),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_330),
.A2(n_305),
.B1(n_303),
.B2(n_324),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_350),
.B(n_324),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_379),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_333),
.B(n_230),
.C(n_243),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_386),
.C(n_357),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_338),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_343),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_380),
.B(n_384),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_347),
.A2(n_303),
.B1(n_300),
.B2(n_286),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_332),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_333),
.B(n_335),
.C(n_339),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_338),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_387),
.B(n_388),
.Y(n_410)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_343),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_354),
.B(n_243),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_389),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_390),
.A2(n_391),
.B1(n_412),
.B2(n_413),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_370),
.A2(n_336),
.B1(n_329),
.B2(n_341),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_395),
.B(n_407),
.C(n_359),
.Y(n_419)
);

BUFx24_ASAP7_75t_SL g401 ( 
.A(n_373),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_401),
.B(n_404),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_385),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_403),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_362),
.B(n_332),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_386),
.B(n_352),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_405),
.B(n_406),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_359),
.B(n_353),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_378),
.B(n_356),
.C(n_349),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_408),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_383),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_409),
.B(n_411),
.Y(n_435)
);

NOR3xp33_ASAP7_75t_L g411 ( 
.A(n_365),
.B(n_337),
.C(n_340),
.Y(n_411)
);

NOR4xp25_ASAP7_75t_L g412 ( 
.A(n_362),
.B(n_300),
.C(n_230),
.D(n_198),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_367),
.A2(n_300),
.B1(n_286),
.B2(n_274),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_376),
.B(n_252),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_414),
.B(n_361),
.Y(n_425)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_379),
.Y(n_418)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_418),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_419),
.B(n_433),
.C(n_230),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_410),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_420),
.B(n_442),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_406),
.B(n_359),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_421),
.B(n_424),
.Y(n_461)
);

OAI22x1_ASAP7_75t_L g423 ( 
.A1(n_408),
.A2(n_394),
.B1(n_374),
.B2(n_369),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_423),
.A2(n_429),
.B1(n_438),
.B2(n_384),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_405),
.B(n_376),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_425),
.B(n_431),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_395),
.B(n_414),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_426),
.B(n_430),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_416),
.A2(n_360),
.B1(n_389),
.B2(n_368),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_427),
.A2(n_400),
.B1(n_274),
.B2(n_231),
.Y(n_459)
);

NOR3xp33_ASAP7_75t_L g428 ( 
.A(n_397),
.B(n_387),
.C(n_366),
.Y(n_428)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_428),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_399),
.A2(n_392),
.B1(n_415),
.B2(n_398),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_407),
.B(n_364),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_390),
.B(n_371),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_393),
.B(n_375),
.C(n_360),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_417),
.A2(n_363),
.B1(n_388),
.B2(n_380),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_391),
.B(n_377),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_413),
.Y(n_455)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_410),
.Y(n_440)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_440),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_393),
.Y(n_442)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_437),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_446),
.B(n_449),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_457),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_432),
.A2(n_402),
.B1(n_417),
.B2(n_408),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_427),
.A2(n_372),
.B1(n_396),
.B2(n_418),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_450),
.B(n_460),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_430),
.B(n_396),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_451),
.B(n_452),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_426),
.B(n_408),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_441),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_453),
.B(n_257),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_455),
.B(n_458),
.Y(n_475)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_435),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_456),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_436),
.A2(n_385),
.B1(n_403),
.B2(n_400),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_421),
.B(n_381),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_459),
.A2(n_423),
.B1(n_433),
.B2(n_439),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_443),
.B(n_419),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_464),
.B(n_466),
.Y(n_480)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_454),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_443),
.B(n_425),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_467),
.B(n_476),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_460),
.B(n_424),
.C(n_422),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_468),
.B(n_472),
.C(n_473),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_455),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_444),
.A2(n_434),
.B(n_431),
.Y(n_470)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_470),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_452),
.B(n_422),
.C(n_441),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_447),
.B(n_231),
.C(n_246),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_447),
.B(n_263),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_451),
.B(n_263),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_477),
.B(n_461),
.Y(n_486)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_478),
.Y(n_491)
);

NOR2xp67_ASAP7_75t_L g479 ( 
.A(n_471),
.B(n_445),
.Y(n_479)
);

OAI211xp5_ASAP7_75t_SL g505 ( 
.A1(n_479),
.A2(n_62),
.B(n_20),
.C(n_3),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_481),
.B(n_489),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_465),
.A2(n_459),
.B1(n_458),
.B2(n_449),
.Y(n_482)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_482),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_469),
.A2(n_457),
.B(n_461),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_485),
.A2(n_493),
.B(n_482),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_486),
.B(n_487),
.Y(n_500)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_462),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_463),
.B(n_240),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_488),
.B(n_492),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_465),
.A2(n_257),
.B1(n_182),
.B2(n_246),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_211),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_472),
.A2(n_202),
.B(n_169),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_473),
.A2(n_152),
.B1(n_120),
.B2(n_3),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_494),
.B(n_491),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_480),
.B(n_484),
.C(n_483),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_496),
.B(n_502),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_481),
.B(n_474),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_497),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_498),
.B(n_507),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_485),
.A2(n_475),
.B(n_468),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_499),
.A2(n_504),
.B(n_1),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_484),
.B(n_475),
.Y(n_502)
);

AND2x6_ASAP7_75t_L g504 ( 
.A(n_487),
.B(n_85),
.Y(n_504)
);

AOI21x1_ASAP7_75t_L g511 ( 
.A1(n_505),
.A2(n_493),
.B(n_4),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_490),
.B(n_20),
.C(n_2),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_506),
.A2(n_1),
.B(n_3),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_503),
.B(n_489),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_509),
.B(n_510),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_511),
.A2(n_512),
.B(n_504),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_20),
.Y(n_512)
);

NOR2xp67_ASAP7_75t_SL g518 ( 
.A(n_513),
.B(n_499),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_516),
.B(n_518),
.Y(n_521)
);

NOR2x1_ASAP7_75t_L g519 ( 
.A(n_515),
.B(n_497),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_519),
.B(n_520),
.Y(n_523)
);

NOR2xp67_ASAP7_75t_SL g520 ( 
.A(n_508),
.B(n_514),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_517),
.B(n_495),
.C(n_512),
.Y(n_522)
);

NOR3xp33_ASAP7_75t_L g524 ( 
.A(n_522),
.B(n_501),
.C(n_495),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_524),
.A2(n_525),
.B(n_523),
.Y(n_526)
);

OAI311xp33_ASAP7_75t_L g525 ( 
.A1(n_521),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.C1(n_7),
.Y(n_525)
);

A2O1A1Ixp33_ASAP7_75t_SL g527 ( 
.A1(n_526),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_527),
.B(n_5),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_528),
.B(n_7),
.C(n_5),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_529),
.A2(n_5),
.B1(n_6),
.B2(n_365),
.Y(n_530)
);


endmodule