module real_jpeg_149_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_1),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_1),
.B(n_45),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_1),
.B(n_34),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_1),
.B(n_74),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_1),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_1),
.B(n_41),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_1),
.B(n_56),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_1),
.B(n_53),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_2),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_2),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_2),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_2),
.B(n_34),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_2),
.B(n_41),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_2),
.B(n_31),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_2),
.B(n_27),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g26 ( 
.A(n_4),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_4),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_4),
.B(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_4),
.B(n_45),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_4),
.B(n_74),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_8),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_8),
.B(n_41),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_8),
.B(n_31),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_8),
.B(n_34),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_10),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_10),
.B(n_45),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_10),
.B(n_74),
.Y(n_126)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_10),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_10),
.B(n_31),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_10),
.B(n_56),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_10),
.B(n_27),
.Y(n_274)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_11),
.B(n_34),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_11),
.B(n_27),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_11),
.B(n_56),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_11),
.B(n_41),
.Y(n_269)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_12),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_12),
.B(n_74),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_12),
.B(n_45),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_13),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_14),
.B(n_41),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_14),
.B(n_34),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_14),
.B(n_27),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_14),
.B(n_56),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_14),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_14),
.B(n_31),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_171),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_169),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_134),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_19),
.B(n_134),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_83),
.C(n_107),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_20),
.B(n_83),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_59),
.B2(n_60),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_21),
.B(n_61),
.C(n_76),
.Y(n_166)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.C(n_47),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_23),
.B(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_33),
.B2(n_35),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_26),
.B(n_30),
.C(n_33),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_26),
.B(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_26),
.A2(n_32),
.B1(n_181),
.B2(n_182),
.Y(n_237)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_29),
.A2(n_30),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_29),
.A2(n_30),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_30),
.B(n_102),
.C(n_104),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_30),
.B(n_278),
.Y(n_312)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_33),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g187 ( 
.A(n_34),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_36),
.B(n_47),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.C(n_43),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_37),
.B(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_38),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_38),
.B(n_115),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_40),
.A2(n_43),
.B1(n_44),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_40),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_40),
.A2(n_111),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_41),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_45),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_55),
.C(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_52),
.Y(n_57)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_55),
.Y(n_58)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_76),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_70),
.C(n_72),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_62),
.B(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.C(n_67),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_63),
.A2(n_67),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_63),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_64),
.B(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_64),
.B(n_164),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_64),
.B(n_68),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_66),
.A2(n_190),
.B1(n_191),
.B2(n_194),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_66),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_67),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_67),
.A2(n_87),
.B1(n_88),
.B2(n_192),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_133)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_82),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_78),
.A2(n_79),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_79),
.B(n_80),
.C(n_82),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_80),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_98),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_96),
.B2(n_97),
.Y(n_84)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_85),
.B(n_97),
.C(n_98),
.Y(n_155)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_95),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_87),
.A2(n_88),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_87),
.B(n_192),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_88),
.B(n_91),
.C(n_94),
.Y(n_145)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_104),
.B2(n_105),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_103),
.B(n_106),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_113),
.C(n_114),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_104),
.A2(n_105),
.B1(n_113),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_106),
.B(n_115),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_107),
.B(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_124),
.C(n_132),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_108),
.B(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.C(n_116),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_109),
.A2(n_116),
.B1(n_117),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_109),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_112),
.B(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_113),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_114),
.B(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_115),
.B(n_243),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_115),
.B(n_187),
.Y(n_271)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_120),
.C(n_122),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_118),
.A2(n_119),
.B1(n_122),
.B2(n_123),
.Y(n_179)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_120),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_132),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.C(n_129),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_129),
.B(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_129),
.A2(n_130),
.B(n_131),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_134)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_153),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_144),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_138),
.A2(n_139),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_184),
.C(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_142),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_149),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_165),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_201),
.B(n_334),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_199),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_173),
.B(n_199),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_197),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_174),
.B(n_197),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_176),
.B(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_188),
.C(n_195),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_177),
.B(n_207),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_183),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_178),
.B(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_180),
.B(n_183),
.Y(n_245)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_184),
.B(n_185),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_186),
.B(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_188),
.A2(n_189),
.B1(n_195),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_250),
.Y(n_201)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI21xp33_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_227),
.B(n_249),
.Y(n_203)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_204),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_225),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_205),
.B(n_225),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.C(n_222),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_222),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_217),
.C(n_219),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_210),
.A2(n_217),
.B1(n_218),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_210),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.C(n_215),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_211),
.A2(n_212),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_247),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_228),
.B(n_230),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_244),
.C(n_246),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_231),
.A2(n_232),
.B1(n_244),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_237),
.C(n_238),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_233),
.A2(n_234),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_237),
.B(n_238),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.C(n_242),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_241),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_242),
.B(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_244),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_246),
.B(n_329),
.Y(n_328)
);

NOR3xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_332),
.C(n_333),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_326),
.B(n_331),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_314),
.B(n_325),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_300),
.B(n_313),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_281),
.B(n_299),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_264),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_256),
.B(n_264),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_261),
.C(n_263),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_257),
.A2(n_258),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_258),
.A2(n_259),
.B(n_260),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_272),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_265),
.B(n_273),
.C(n_277),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_271),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_267),
.B(n_270),
.C(n_271),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_269),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_276),
.B1(n_277),
.B2(n_280),
.Y(n_272)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_273),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_280),
.A2(n_292),
.B(n_293),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_290),
.B(n_298),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_286),
.B(n_289),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_284),
.B(n_285),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_294),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_291),
.B(n_294),
.Y(n_298)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_301),
.B(n_302),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_308),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_307),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_307),
.C(n_308),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_312),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_311),
.C(n_312),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_315),
.B(n_316),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_320),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_321),
.C(n_322),
.Y(n_327)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_327),
.B(n_328),
.Y(n_331)
);


endmodule