module real_aes_11019_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_85;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_617;
wire n_139;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_87;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_95;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_265;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_283;
wire n_252;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
NAND2xp5_ASAP7_75t_L g592 ( .A(n_0), .B(n_59), .Y(n_592) );
AND2x2_ASAP7_75t_L g602 ( .A(n_0), .B(n_603), .Y(n_602) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_0), .Y(n_630) );
INVx1_ASAP7_75t_L g651 ( .A(n_0), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_1), .B(n_164), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_2), .B(n_126), .Y(n_207) );
INVx2_ASAP7_75t_L g535 ( .A(n_3), .Y(n_535) );
OR2x2_ASAP7_75t_L g561 ( .A(n_3), .B(n_533), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_4), .A2(n_40), .B1(n_569), .B2(n_573), .Y(n_568) );
INVx1_ASAP7_75t_L g660 ( .A(n_4), .Y(n_660) );
INVx1_ASAP7_75t_L g537 ( .A(n_5), .Y(n_537) );
BUFx2_ASAP7_75t_L g582 ( .A(n_5), .Y(n_582) );
BUFx2_ASAP7_75t_L g587 ( .A(n_5), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_6), .B(n_115), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_7), .B(n_107), .Y(n_256) );
NAND2x1p5_ASAP7_75t_L g196 ( .A(n_8), .B(n_107), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_9), .B(n_160), .Y(n_159) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_10), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_11), .A2(n_49), .B1(n_669), .B2(n_674), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_11), .A2(n_49), .B1(n_704), .B2(n_707), .Y(n_703) );
INVx1_ASAP7_75t_L g538 ( .A(n_12), .Y(n_538) );
AND2x2_ASAP7_75t_L g267 ( .A(n_13), .B(n_268), .Y(n_267) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_14), .Y(n_94) );
INVx1_ASAP7_75t_L g509 ( .A(n_15), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_16), .B(n_151), .Y(n_150) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_17), .A2(n_600), .B1(n_605), .B2(n_617), .C(n_632), .Y(n_599) );
AOI22xp33_ASAP7_75t_SL g700 ( .A1(n_17), .A2(n_77), .B1(n_701), .B2(n_702), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_18), .B(n_184), .Y(n_209) );
INVx1_ASAP7_75t_L g616 ( .A(n_19), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_19), .A2(n_61), .B1(n_694), .B2(n_697), .Y(n_693) );
NAND2xp33_ASAP7_75t_L g191 ( .A(n_20), .B(n_192), .Y(n_191) );
NAND2xp33_ASAP7_75t_L g254 ( .A(n_21), .B(n_192), .Y(n_254) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_22), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_23), .Y(n_114) );
INVx1_ASAP7_75t_L g719 ( .A(n_24), .Y(n_719) );
INVx1_ASAP7_75t_L g533 ( .A(n_25), .Y(n_533) );
INVx1_ASAP7_75t_L g686 ( .A(n_25), .Y(n_686) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_26), .B(n_147), .Y(n_195) );
OAI21x1_ASAP7_75t_L g109 ( .A1(n_27), .A2(n_52), .B(n_110), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_28), .A2(n_121), .B(n_273), .C(n_274), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_29), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_30), .B(n_119), .Y(n_141) );
NAND2xp33_ASAP7_75t_L g165 ( .A(n_31), .B(n_125), .Y(n_165) );
AND2x6_ASAP7_75t_L g84 ( .A(n_32), .B(n_85), .Y(n_84) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_32), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_32), .B(n_727), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_33), .B(n_118), .Y(n_181) );
AOI22xp33_ASAP7_75t_SL g741 ( .A1(n_34), .A2(n_517), .B1(n_518), .B2(n_742), .Y(n_741) );
CKINVDCx5p33_ASAP7_75t_R g742 ( .A(n_34), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_35), .B(n_253), .Y(n_252) );
NAND2xp33_ASAP7_75t_L g208 ( .A(n_36), .B(n_125), .Y(n_208) );
INVx1_ASAP7_75t_L g85 ( .A(n_37), .Y(n_85) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_37), .Y(n_727) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_38), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_39), .A2(n_715), .B1(n_716), .B2(n_717), .Y(n_714) );
CKINVDCx5p33_ASAP7_75t_R g715 ( .A(n_39), .Y(n_715) );
INVx1_ASAP7_75t_L g645 ( .A(n_40), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_41), .B(n_125), .Y(n_158) );
INVx1_ASAP7_75t_L g567 ( .A(n_42), .Y(n_567) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_43), .Y(n_512) );
INVx1_ASAP7_75t_L g562 ( .A(n_44), .Y(n_562) );
INVx1_ASAP7_75t_L g546 ( .A(n_45), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_46), .Y(n_139) );
AND2x2_ASAP7_75t_L g276 ( .A(n_47), .B(n_184), .Y(n_276) );
INVx1_ASAP7_75t_L g622 ( .A(n_48), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_48), .A2(n_55), .B1(n_688), .B2(n_691), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_50), .B(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g596 ( .A(n_51), .Y(n_596) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_53), .Y(n_194) );
NAND2xp33_ASAP7_75t_L g176 ( .A(n_54), .B(n_90), .Y(n_176) );
INVx1_ASAP7_75t_L g626 ( .A(n_55), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_56), .B(n_164), .Y(n_163) );
BUFx10_ASAP7_75t_L g736 ( .A(n_57), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_58), .B(n_89), .Y(n_250) );
INVx2_ASAP7_75t_L g603 ( .A(n_59), .Y(n_603) );
INVx1_ASAP7_75t_L g631 ( .A(n_59), .Y(n_631) );
NAND2xp33_ASAP7_75t_L g182 ( .A(n_60), .B(n_115), .Y(n_182) );
INVx1_ASAP7_75t_L g611 ( .A(n_61), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_62), .B(n_192), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_63), .Y(n_275) );
INVx2_ASAP7_75t_L g110 ( .A(n_64), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_65), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_66), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_67), .B(n_151), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_68), .Y(n_203) );
INVx1_ASAP7_75t_L g579 ( .A(n_69), .Y(n_579) );
INVx1_ASAP7_75t_L g266 ( .A(n_70), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_71), .Y(n_117) );
AND2x2_ASAP7_75t_L g131 ( .A(n_72), .B(n_107), .Y(n_131) );
INVx2_ASAP7_75t_L g597 ( .A(n_73), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_74), .B(n_184), .Y(n_183) );
BUFx3_ASAP7_75t_L g545 ( .A(n_75), .Y(n_545) );
INVx1_ASAP7_75t_L g572 ( .A(n_75), .Y(n_572) );
BUFx3_ASAP7_75t_L g528 ( .A(n_76), .Y(n_528) );
INVx1_ASAP7_75t_L g558 ( .A(n_76), .Y(n_558) );
OAI221xp5_ASAP7_75t_L g635 ( .A1(n_77), .A2(n_636), .B1(n_643), .B2(n_652), .C(n_661), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_95), .B(n_504), .Y(n_78) );
BUFx2_ASAP7_75t_SL g79 ( .A(n_80), .Y(n_79) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_86), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
AOI21xp5_ASAP7_75t_L g111 ( .A1(n_83), .A2(n_112), .B(n_122), .Y(n_111) );
INVx8_ASAP7_75t_L g149 ( .A(n_83), .Y(n_149) );
NOR2xp67_ASAP7_75t_L g261 ( .A(n_83), .B(n_262), .Y(n_261) );
INVx8_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
BUFx2_ASAP7_75t_L g166 ( .A(n_84), .Y(n_166) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_87), .Y(n_86) );
AO21x1_ASAP7_75t_L g756 ( .A1(n_87), .A2(n_757), .B(n_758), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g87 ( .A(n_88), .B(n_92), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g140 ( .A(n_89), .Y(n_140) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx2_ASAP7_75t_L g160 ( .A(n_90), .Y(n_160) );
INVx2_ASAP7_75t_L g178 ( .A(n_90), .Y(n_178) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_91), .Y(n_115) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_91), .Y(n_119) );
INVx2_ASAP7_75t_L g126 ( .A(n_91), .Y(n_126) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_91), .Y(n_129) );
INVx1_ASAP7_75t_L g270 ( .A(n_91), .Y(n_270) );
OAI21xp33_ASAP7_75t_L g122 ( .A1(n_92), .A2(n_123), .B(n_127), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_92), .A2(n_249), .B(n_250), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_93), .Y(n_92) );
INVx3_ASAP7_75t_L g148 ( .A(n_93), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_93), .A2(n_163), .B(n_165), .Y(n_162) );
BUFx2_ASAP7_75t_L g271 ( .A(n_93), .Y(n_271) );
BUFx12f_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx5_ASAP7_75t_L g121 ( .A(n_94), .Y(n_121) );
O2A1O1Ixp33_ASAP7_75t_L g138 ( .A1(n_94), .A2(n_139), .B(n_140), .C(n_141), .Y(n_138) );
INVx5_ASAP7_75t_L g161 ( .A(n_94), .Y(n_161) );
INVx2_ASAP7_75t_SL g95 ( .A(n_96), .Y(n_95) );
AND2x4_ASAP7_75t_L g96 ( .A(n_97), .B(n_403), .Y(n_96) );
NOR3xp33_ASAP7_75t_L g97 ( .A(n_98), .B(n_321), .C(n_354), .Y(n_97) );
OAI211xp5_ASAP7_75t_L g98 ( .A1(n_99), .A2(n_132), .B(n_241), .C(n_306), .Y(n_98) );
INVxp67_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g328 ( .A(n_104), .B(n_259), .Y(n_328) );
INVx2_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_105), .B(n_212), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_105), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g386 ( .A(n_105), .Y(n_386) );
AO21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_111), .B(n_131), .Y(n_105) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_106), .A2(n_111), .B(n_131), .Y(n_258) );
INVx3_ASAP7_75t_L g262 ( .A(n_106), .Y(n_262) );
INVx4_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx4f_ASAP7_75t_L g136 ( .A(n_107), .Y(n_136) );
INVx3_ASAP7_75t_L g155 ( .A(n_107), .Y(n_155) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_107), .A2(n_174), .B(n_183), .Y(n_173) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_107), .A2(n_174), .B(n_183), .Y(n_218) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_107), .A2(n_174), .B(n_183), .Y(n_240) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g152 ( .A(n_108), .Y(n_152) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g185 ( .A(n_109), .Y(n_185) );
OAI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_116), .B(n_120), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_114), .A2(n_718), .B1(n_719), .B2(n_720), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_114), .Y(n_720) );
INVx2_ASAP7_75t_L g145 ( .A(n_115), .Y(n_145) );
INVx2_ASAP7_75t_L g164 ( .A(n_115), .Y(n_164) );
INVx2_ASAP7_75t_SL g253 ( .A(n_115), .Y(n_253) );
NOR2xp67_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
INVx5_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
CKINVDCx6p67_ASAP7_75t_R g179 ( .A(n_121), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g147 ( .A(n_126), .Y(n_147) );
INVx2_ASAP7_75t_L g192 ( .A(n_126), .Y(n_192) );
NOR2xp33_ASAP7_75t_SL g127 ( .A(n_128), .B(n_130), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_128), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AOI311xp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_168), .A3(n_197), .B(n_210), .C(n_226), .Y(n_132) );
AND2x2_ASAP7_75t_L g283 ( .A(n_133), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g375 ( .A(n_133), .Y(n_375) );
BUFx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g337 ( .A(n_134), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_134), .B(n_171), .Y(n_489) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_153), .Y(n_134) );
AND2x2_ASAP7_75t_L g298 ( .A(n_135), .B(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g308 ( .A(n_135), .B(n_224), .Y(n_308) );
INVx1_ASAP7_75t_L g319 ( .A(n_135), .Y(n_319) );
OAI21x1_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_137), .B(n_150), .Y(n_135) );
OA21x2_ASAP7_75t_L g187 ( .A1(n_136), .A2(n_188), .B(n_196), .Y(n_187) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_136), .A2(n_201), .B(n_209), .Y(n_200) );
OAI21x1_ASAP7_75t_L g217 ( .A1(n_136), .A2(n_137), .B(n_150), .Y(n_217) );
OAI21x1_ASAP7_75t_L g223 ( .A1(n_136), .A2(n_188), .B(n_196), .Y(n_223) );
OAI21x1_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_142), .B(n_149), .Y(n_137) );
INVx1_ASAP7_75t_L g754 ( .A(n_139), .Y(n_754) );
O2A1O1Ixp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_146), .C(n_148), .Y(n_142) );
OAI22xp33_ASAP7_75t_L g752 ( .A1(n_143), .A2(n_517), .B1(n_518), .B2(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_143), .Y(n_753) );
O2A1O1Ixp5_ASAP7_75t_L g193 ( .A1(n_144), .A2(n_148), .B(n_194), .C(n_195), .Y(n_193) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
O2A1O1Ixp5_ASAP7_75t_L g202 ( .A1(n_148), .A2(n_203), .B(n_204), .C(n_205), .Y(n_202) );
OAI21x1_ASAP7_75t_L g174 ( .A1(n_149), .A2(n_175), .B(n_180), .Y(n_174) );
OAI21x1_ASAP7_75t_L g188 ( .A1(n_149), .A2(n_189), .B(n_193), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g201 ( .A1(n_149), .A2(n_202), .B(n_206), .Y(n_201) );
OAI21x1_ASAP7_75t_L g247 ( .A1(n_149), .A2(n_248), .B(n_251), .Y(n_247) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx2_ASAP7_75t_L g434 ( .A(n_153), .Y(n_434) );
OAI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_156), .B(n_167), .Y(n_153) );
OAI21x1_ASAP7_75t_L g225 ( .A1(n_154), .A2(n_156), .B(n_167), .Y(n_225) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_154), .A2(n_247), .B(n_256), .Y(n_246) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
OAI21x1_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_162), .B(n_166), .Y(n_156) );
AOI21x1_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_161), .Y(n_157) );
INVx1_ASAP7_75t_L g204 ( .A(n_160), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_161), .A2(n_181), .B(n_182), .Y(n_180) );
INVx1_ASAP7_75t_L g255 ( .A(n_161), .Y(n_255) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVxp67_ASAP7_75t_SL g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g449 ( .A(n_171), .Y(n_449) );
NAND2x1p5_ASAP7_75t_L g171 ( .A(n_172), .B(n_186), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
OR2x2_ASAP7_75t_L g340 ( .A(n_173), .B(n_299), .Y(n_340) );
AND2x2_ASAP7_75t_L g402 ( .A(n_173), .B(n_299), .Y(n_402) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_179), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_179), .A2(n_190), .B(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_179), .A2(n_207), .B(n_208), .Y(n_206) );
BUFx5_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g284 ( .A(n_186), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_186), .B(n_216), .Y(n_452) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g479 ( .A(n_187), .B(n_294), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_192), .B(n_275), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_194), .A2(n_714), .B1(n_721), .B2(n_722), .Y(n_713) );
INVx1_ASAP7_75t_L g721 ( .A(n_194), .Y(n_721) );
INVxp67_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x4_ASAP7_75t_L g367 ( .A(n_198), .B(n_368), .Y(n_367) );
AOI32xp33_ASAP7_75t_L g393 ( .A1(n_198), .A2(n_394), .A3(n_397), .B1(n_398), .B2(n_400), .Y(n_393) );
AND2x4_ASAP7_75t_L g493 ( .A(n_198), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_199), .B(n_282), .Y(n_334) );
OR2x2_ASAP7_75t_L g345 ( .A(n_199), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_199), .B(n_281), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_199), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g416 ( .A(n_199), .B(n_245), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_199), .B(n_368), .Y(n_484) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g212 ( .A(n_200), .Y(n_212) );
AND2x2_ASAP7_75t_L g312 ( .A(n_200), .B(n_258), .Y(n_312) );
NOR3xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_213), .C(n_219), .Y(n_210) );
INVx1_ASAP7_75t_L g237 ( .A(n_211), .Y(n_237) );
AND2x2_ASAP7_75t_L g461 ( .A(n_211), .B(n_328), .Y(n_461) );
AND2x2_ASAP7_75t_L g469 ( .A(n_211), .B(n_430), .Y(n_469) );
BUFx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
OR2x2_ASAP7_75t_L g325 ( .A(n_212), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g358 ( .A(n_212), .B(n_246), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_218), .Y(n_213) );
OAI211xp5_ASAP7_75t_SL g321 ( .A1(n_214), .A2(n_322), .B(n_329), .C(n_348), .Y(n_321) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
BUFx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g390 ( .A(n_216), .Y(n_390) );
AND2x4_ASAP7_75t_SL g442 ( .A(n_216), .B(n_293), .Y(n_442) );
NAND2x1_ASAP7_75t_L g474 ( .A(n_216), .B(n_377), .Y(n_474) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g231 ( .A(n_217), .Y(n_231) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_217), .Y(n_465) );
INVx2_ASAP7_75t_L g419 ( .A(n_218), .Y(n_419) );
INVx2_ASAP7_75t_L g430 ( .A(n_218), .Y(n_430) );
AND2x2_ASAP7_75t_L g498 ( .A(n_218), .B(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
OR2x2_ASAP7_75t_L g350 ( .A(n_220), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x4_ASAP7_75t_L g347 ( .A(n_221), .B(n_230), .Y(n_347) );
AND2x2_ASAP7_75t_L g388 ( .A(n_221), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_224), .Y(n_221) );
INVx2_ASAP7_75t_L g299 ( .A(n_222), .Y(n_299) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g235 ( .A(n_223), .B(n_224), .Y(n_235) );
INVx2_ASAP7_75t_L g294 ( .A(n_224), .Y(n_294) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NOR3xp33_ASAP7_75t_L g226 ( .A(n_227), .B(n_232), .C(n_236), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
BUFx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x4_ASAP7_75t_L g292 ( .A(n_230), .B(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AOI21xp33_ASAP7_75t_L g450 ( .A1(n_232), .A2(n_451), .B(n_453), .Y(n_450) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g427 ( .A(n_235), .B(n_239), .Y(n_427) );
NAND2xp33_ASAP7_75t_R g438 ( .A(n_235), .B(n_318), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NOR2xp67_ASAP7_75t_L g330 ( .A(n_239), .B(n_331), .Y(n_330) );
BUFx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx2_ASAP7_75t_SL g291 ( .A(n_240), .Y(n_291) );
INVx1_ASAP7_75t_L g351 ( .A(n_240), .Y(n_351) );
INVx1_ASAP7_75t_SL g396 ( .A(n_240), .Y(n_396) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_283), .B(n_285), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_277), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_257), .Y(n_243) );
OR2x2_ASAP7_75t_L g314 ( .A(n_244), .B(n_279), .Y(n_314) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g305 ( .A(n_246), .Y(n_305) );
AND2x2_ASAP7_75t_L g310 ( .A(n_246), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g326 ( .A(n_246), .Y(n_326) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_246), .Y(n_346) );
OR2x2_ASAP7_75t_L g369 ( .A(n_246), .B(n_258), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_254), .B(n_255), .Y(n_251) );
INVx2_ASAP7_75t_L g273 ( .A(n_253), .Y(n_273) );
AND2x2_ASAP7_75t_L g352 ( .A(n_257), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g423 ( .A(n_257), .Y(n_423) );
AND2x2_ASAP7_75t_L g443 ( .A(n_257), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g445 ( .A(n_257), .B(n_358), .Y(n_445) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
AND2x2_ASAP7_75t_L g458 ( .A(n_258), .B(n_411), .Y(n_458) );
INVx1_ASAP7_75t_L g311 ( .A(n_259), .Y(n_311) );
INVx1_ASAP7_75t_L g411 ( .A(n_259), .Y(n_411) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g282 ( .A(n_260), .Y(n_282) );
AOI21x1_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_263), .B(n_276), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_272), .Y(n_263) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_267), .B(n_271), .Y(n_264) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OAI32xp33_ASAP7_75t_L g467 ( .A1(n_277), .A2(n_468), .A3(n_470), .B1(n_471), .B2(n_473), .Y(n_467) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g287 ( .A(n_279), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g302 ( .A(n_282), .Y(n_302) );
INVxp67_ASAP7_75t_SL g344 ( .A(n_282), .Y(n_344) );
OR2x2_ASAP7_75t_L g432 ( .A(n_284), .B(n_433), .Y(n_432) );
OAI22xp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_288), .B1(n_295), .B2(n_300), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_289), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g324 ( .A(n_290), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g362 ( .A(n_291), .B(n_299), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_291), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g320 ( .A(n_292), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_292), .A2(n_383), .B1(n_388), .B2(n_391), .Y(n_382) );
AND2x2_ASAP7_75t_L g394 ( .A(n_292), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g297 ( .A(n_293), .Y(n_297) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_294), .B(n_299), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_295), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx1_ASAP7_75t_L g381 ( .A(n_298), .Y(n_381) );
INVx1_ASAP7_75t_L g377 ( .A(n_299), .Y(n_377) );
OAI22xp33_ASAP7_75t_L g496 ( .A1(n_300), .A2(n_497), .B1(n_501), .B2(n_502), .Y(n_496) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g415 ( .A(n_302), .Y(n_415) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g333 ( .A(n_304), .B(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g379 ( .A(n_304), .B(n_374), .Y(n_379) );
INVx1_ASAP7_75t_L g426 ( .A(n_305), .Y(n_426) );
A2O1A1Ixp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_309), .B(n_313), .C(n_315), .Y(n_306) );
NAND2x1_ASAP7_75t_SL g360 ( .A(n_307), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_307), .B(n_339), .Y(n_407) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND3xp33_ASAP7_75t_L g315 ( .A(n_308), .B(n_316), .C(n_320), .Y(n_315) );
OR2x6_ASAP7_75t_SL g418 ( .A(n_308), .B(n_419), .Y(n_418) );
INVx2_ASAP7_75t_SL g331 ( .A(n_309), .Y(n_331) );
AND2x4_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx1_ASAP7_75t_L g387 ( .A(n_310), .Y(n_387) );
AND2x2_ASAP7_75t_L g494 ( .A(n_310), .B(n_386), .Y(n_494) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AOI222xp33_ASAP7_75t_L g329 ( .A1(n_320), .A2(n_330), .B1(n_332), .B2(n_335), .C1(n_341), .C2(n_347), .Y(n_329) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NOR2x1_ASAP7_75t_L g323 ( .A(n_324), .B(n_327), .Y(n_323) );
INVx1_ASAP7_75t_L g353 ( .A(n_325), .Y(n_353) );
INVx1_ASAP7_75t_SL g399 ( .A(n_325), .Y(n_399) );
INVx1_ASAP7_75t_L g397 ( .A(n_327), .Y(n_397) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g398 ( .A(n_328), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g425 ( .A(n_328), .B(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g436 ( .A(n_328), .B(n_358), .Y(n_436) );
INVx2_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g392 ( .A(n_334), .Y(n_392) );
NOR2xp67_ASAP7_75t_SL g335 ( .A(n_336), .B(n_338), .Y(n_335) );
AND2x2_ASAP7_75t_L g455 ( .A(n_336), .B(n_395), .Y(n_455) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NOR2x1_ASAP7_75t_SL g412 ( .A(n_337), .B(n_362), .Y(n_412) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g466 ( .A(n_340), .Y(n_466) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_343), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g486 ( .A(n_343), .B(n_353), .Y(n_486) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g421 ( .A(n_345), .Y(n_421) );
OR2x2_ASAP7_75t_L g453 ( .A(n_345), .B(n_423), .Y(n_453) );
AND2x2_ASAP7_75t_L g429 ( .A(n_347), .B(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_352), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g451 ( .A(n_351), .B(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g473 ( .A(n_351), .B(n_474), .Y(n_473) );
OR2x2_ASAP7_75t_L g502 ( .A(n_351), .B(n_503), .Y(n_502) );
NAND4xp25_ASAP7_75t_L g354 ( .A(n_355), .B(n_370), .C(n_382), .D(n_393), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_359), .B1(n_363), .B2(n_365), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g408 ( .A(n_358), .B(n_409), .Y(n_408) );
NAND2xp67_ASAP7_75t_L g457 ( .A(n_358), .B(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AO21x1_ASAP7_75t_L g477 ( .A1(n_361), .A2(n_442), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_362), .Y(n_364) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g391 ( .A(n_368), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVxp67_ASAP7_75t_SL g372 ( .A(n_369), .Y(n_372) );
OR2x2_ASAP7_75t_L g462 ( .A(n_369), .B(n_410), .Y(n_462) );
AOI32xp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_375), .A3(n_376), .B1(n_378), .B2(n_380), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx1_ASAP7_75t_L g501 ( .A(n_372), .Y(n_501) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_378), .A2(n_400), .B1(n_477), .B2(n_480), .C(n_482), .Y(n_476) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
BUFx2_ASAP7_75t_SL g472 ( .A(n_386), .Y(n_472) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g448 ( .A(n_390), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g495 ( .A(n_398), .B(n_478), .Y(n_495) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NOR2x1_ASAP7_75t_L g403 ( .A(n_404), .B(n_475), .Y(n_403) );
NAND4xp25_ASAP7_75t_L g404 ( .A(n_405), .B(n_428), .C(n_439), .D(n_454), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_408), .B1(n_412), .B2(n_413), .C(n_417), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g428 ( .A1(n_408), .A2(n_429), .B(n_431), .Y(n_428) );
INVx1_ASAP7_75t_L g470 ( .A(n_409), .Y(n_470) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
OAI31xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_420), .A3(n_422), .B(n_424), .Y(n_417) );
NAND2xp33_ASAP7_75t_L g446 ( .A(n_418), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g478 ( .A(n_419), .B(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_419), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND2x1p5_ASAP7_75t_L g424 ( .A(n_425), .B(n_427), .Y(n_424) );
INVx1_ASAP7_75t_L g437 ( .A(n_425), .Y(n_437) );
INVx1_ASAP7_75t_L g444 ( .A(n_426), .Y(n_444) );
INVx1_ASAP7_75t_L g483 ( .A(n_427), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_430), .B(n_442), .Y(n_441) );
OAI22xp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_435), .B1(n_437), .B2(n_438), .Y(n_431) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_443), .B1(n_445), .B2(n_446), .C(n_450), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_442), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g492 ( .A(n_442), .Y(n_492) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B1(n_459), .B2(n_463), .C(n_467), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_457), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x4_ASAP7_75t_L g463 ( .A(n_464), .B(n_466), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVxp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_490), .Y(n_475) );
INVx2_ASAP7_75t_L g503 ( .A(n_479), .Y(n_503) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B1(n_485), .B2(n_487), .Y(n_482) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AOI211xp5_ASAP7_75t_SL g490 ( .A1(n_491), .A2(n_493), .B(n_495), .C(n_496), .Y(n_490) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OAI221xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_723), .B1(n_741), .B2(n_743), .C(n_747), .Y(n_504) );
XNOR2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_713), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_507), .A2(n_508), .B1(n_517), .B2(n_518), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B1(n_511), .B2(n_516), .Y(n_508) );
INVx1_ASAP7_75t_L g516 ( .A(n_509), .Y(n_516) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B1(n_514), .B2(n_515), .Y(n_511) );
INVx1_ASAP7_75t_L g515 ( .A(n_512), .Y(n_515) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NAND4xp75_ASAP7_75t_SL g519 ( .A(n_520), .B(n_578), .C(n_598), .D(n_681), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_553), .Y(n_520) );
AOI221xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_538), .B1(n_539), .B2(n_546), .C(n_547), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2x1p5_ASAP7_75t_L g523 ( .A(n_524), .B(n_529), .Y(n_523) );
INVx1_ASAP7_75t_L g734 ( .A(n_524), .Y(n_734) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g740 ( .A(n_525), .Y(n_740) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x4_ASAP7_75t_L g566 ( .A(n_527), .B(n_544), .Y(n_566) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g551 ( .A(n_528), .B(n_545), .Y(n_551) );
AND2x4_ASAP7_75t_L g571 ( .A(n_528), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
OR2x6_ASAP7_75t_L g540 ( .A(n_530), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g552 ( .A(n_530), .Y(n_552) );
NAND2x1p5_ASAP7_75t_L g530 ( .A(n_531), .B(n_536), .Y(n_530) );
AND2x2_ASAP7_75t_L g583 ( .A(n_531), .B(n_566), .Y(n_583) );
AND2x4_ASAP7_75t_L g739 ( .A(n_531), .B(n_740), .Y(n_739) );
AND2x4_ASAP7_75t_L g531 ( .A(n_532), .B(n_534), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x4_ASAP7_75t_L g712 ( .A(n_534), .B(n_686), .Y(n_712) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g685 ( .A(n_535), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g560 ( .A(n_537), .B(n_561), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_538), .A2(n_546), .B1(n_662), .B2(n_665), .Y(n_661) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x4_ASAP7_75t_L g557 ( .A(n_545), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_552), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx6f_ASAP7_75t_L g692 ( .A(n_551), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_562), .B1(n_563), .B2(n_567), .C(n_568), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_559), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_557), .Y(n_696) );
BUFx6f_ASAP7_75t_L g706 ( .A(n_557), .Y(n_706) );
INVx1_ASAP7_75t_L g577 ( .A(n_558), .Y(n_577) );
AND2x2_ASAP7_75t_L g563 ( .A(n_559), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OR2x6_ASAP7_75t_L g569 ( .A(n_560), .B(n_570), .Y(n_569) );
OR2x6_ASAP7_75t_L g573 ( .A(n_560), .B(n_574), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_562), .A2(n_653), .B1(n_656), .B2(n_660), .Y(n_652) );
INVx2_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g701 ( .A(n_565), .Y(n_701) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx6_ASAP7_75t_L g690 ( .A(n_566), .Y(n_690) );
OAI221xp5_ASAP7_75t_L g643 ( .A1(n_567), .A2(n_623), .B1(n_644), .B2(n_645), .C(n_646), .Y(n_643) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
BUFx6f_ASAP7_75t_L g699 ( .A(n_571), .Y(n_699) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_571), .Y(n_709) );
INVx1_ASAP7_75t_L g576 ( .A(n_572), .Y(n_576) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
OR2x6_ASAP7_75t_L g580 ( .A(n_581), .B(n_584), .Y(n_580) );
AND2x4_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
AND2x4_ASAP7_75t_L g711 ( .A(n_582), .B(n_712), .Y(n_711) );
NOR2xp67_ASAP7_75t_L g584 ( .A(n_585), .B(n_588), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OR2x6_ASAP7_75t_L g683 ( .A(n_586), .B(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx2_ASAP7_75t_L g680 ( .A(n_587), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_593), .Y(n_588) );
AND2x2_ASAP7_75t_L g662 ( .A(n_589), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x6_ASAP7_75t_L g632 ( .A(n_590), .B(n_633), .Y(n_632) );
OR2x6_ASAP7_75t_L g666 ( .A(n_590), .B(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
INVx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_595), .Y(n_604) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_596), .B(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g615 ( .A(n_596), .Y(n_615) );
INVx1_ASAP7_75t_L g620 ( .A(n_596), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_596), .B(n_597), .Y(n_625) );
INVx1_ASAP7_75t_L g664 ( .A(n_596), .Y(n_664) );
INVx1_ASAP7_75t_L g673 ( .A(n_596), .Y(n_673) );
INVx2_ASAP7_75t_L g610 ( .A(n_597), .Y(n_610) );
AND2x4_ASAP7_75t_L g614 ( .A(n_597), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g621 ( .A(n_597), .Y(n_621) );
INVx1_ASAP7_75t_L g642 ( .A(n_597), .Y(n_642) );
OAI31xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_635), .A3(n_668), .B(n_678), .Y(n_598) );
CKINVDCx6p67_ASAP7_75t_R g600 ( .A(n_601), .Y(n_600) );
AND2x4_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx2_ASAP7_75t_L g639 ( .A(n_602), .Y(n_639) );
AND2x2_ASAP7_75t_L g670 ( .A(n_602), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g650 ( .A(n_603), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_611), .B1(n_612), .B2(n_616), .Y(n_605) );
INVx2_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
BUFx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g655 ( .A(n_609), .Y(n_655) );
INVx1_ASAP7_75t_L g667 ( .A(n_610), .Y(n_667) );
AND2x4_ASAP7_75t_L g671 ( .A(n_610), .B(n_672), .Y(n_671) );
INVx2_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx3_ASAP7_75t_L g659 ( .A(n_614), .Y(n_659) );
INVx1_ASAP7_75t_L g677 ( .A(n_614), .Y(n_677) );
AND2x4_ASAP7_75t_L g641 ( .A(n_615), .B(n_642), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_622), .B1(n_623), .B2(n_626), .C(n_627), .Y(n_617) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
AND2x2_ASAP7_75t_L g634 ( .A(n_620), .B(n_621), .Y(n_634) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
BUFx2_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx3_ASAP7_75t_L g644 ( .A(n_634), .Y(n_644) );
INVx8_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x4_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
AND2x4_ASAP7_75t_L g675 ( .A(n_638), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
BUFx3_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2x1p5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
BUFx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx3_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
CKINVDCx11_ASAP7_75t_R g665 ( .A(n_666), .Y(n_665) );
INVx3_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx3_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
BUFx8_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AOI33xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_687), .A3(n_693), .B1(n_700), .B2(n_703), .B3(n_710), .Y(n_681) );
CKINVDCx5p33_ASAP7_75t_R g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_SL g732 ( .A(n_685), .Y(n_732) );
BUFx3_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
BUFx4f_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
BUFx3_ASAP7_75t_L g702 ( .A(n_692), .Y(n_702) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
BUFx4f_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g722 ( .A(n_714), .Y(n_722) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx8_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
CKINVDCx20_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OR2x6_ASAP7_75t_L g725 ( .A(n_726), .B(n_729), .Y(n_725) );
OR2x4_ASAP7_75t_L g751 ( .A(n_726), .B(n_730), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_727), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_SL g757 ( .A(n_727), .Y(n_757) );
INVx1_ASAP7_75t_L g746 ( .A(n_728), .Y(n_746) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AOI31xp33_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_733), .A3(n_735), .B(n_737), .Y(n_730) );
BUFx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx6_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVxp67_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_752), .B1(n_754), .B2(n_755), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx8_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
BUFx2_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
endmodule