module fake_netlist_1_212_n_818 (n_117, n_44, n_133, n_149, n_81, n_69, n_214, n_204, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_96, n_39, n_818);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_96;
input n_39;
output n_818;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_808;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_567;
wire n_809;
wire n_580;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_230;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_810;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_446;
wire n_420;
wire n_285;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_774;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_146), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_137), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_25), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_193), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_157), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_154), .Y(n_221) );
BUFx3_ASAP7_75t_L g222 ( .A(n_93), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_14), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_111), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_192), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_58), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_55), .Y(n_227) );
INVxp67_ASAP7_75t_SL g228 ( .A(n_96), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_191), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_8), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_77), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_12), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_93), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_134), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_160), .Y(n_235) );
CKINVDCx16_ASAP7_75t_R g236 ( .A(n_161), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_128), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_207), .Y(n_238) );
INVx1_ASAP7_75t_SL g239 ( .A(n_167), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_7), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_158), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_165), .Y(n_242) );
BUFx5_ASAP7_75t_L g243 ( .A(n_76), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_54), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_119), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_9), .Y(n_246) );
INVxp67_ASAP7_75t_SL g247 ( .A(n_107), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_79), .Y(n_248) );
CKINVDCx16_ASAP7_75t_R g249 ( .A(n_168), .Y(n_249) );
CKINVDCx16_ASAP7_75t_R g250 ( .A(n_164), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_78), .Y(n_251) );
BUFx3_ASAP7_75t_L g252 ( .A(n_38), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_210), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_138), .Y(n_254) );
CKINVDCx16_ASAP7_75t_R g255 ( .A(n_0), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_200), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_123), .Y(n_257) );
BUFx8_ASAP7_75t_SL g258 ( .A(n_47), .Y(n_258) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_145), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_142), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_122), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_150), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_124), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_215), .Y(n_264) );
BUFx3_ASAP7_75t_L g265 ( .A(n_186), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_176), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_60), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_163), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_209), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_6), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_136), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_169), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_174), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_80), .Y(n_274) );
NOR2xp67_ASAP7_75t_L g275 ( .A(n_198), .B(n_26), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_29), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_31), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_32), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_208), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_177), .Y(n_280) );
BUFx3_ASAP7_75t_L g281 ( .A(n_179), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_205), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_51), .Y(n_283) );
CKINVDCx14_ASAP7_75t_R g284 ( .A(n_144), .Y(n_284) );
CKINVDCx20_ASAP7_75t_R g285 ( .A(n_27), .Y(n_285) );
NOR2xp67_ASAP7_75t_L g286 ( .A(n_166), .B(n_183), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_82), .Y(n_287) );
INVxp67_ASAP7_75t_L g288 ( .A(n_63), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_202), .Y(n_289) );
INVx1_ASAP7_75t_SL g290 ( .A(n_132), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_97), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_141), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_69), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_159), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_173), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_199), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_94), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_139), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_133), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_115), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_34), .Y(n_301) );
CKINVDCx16_ASAP7_75t_R g302 ( .A(n_175), .Y(n_302) );
BUFx3_ASAP7_75t_L g303 ( .A(n_206), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_55), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_152), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_135), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_94), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g308 ( .A(n_98), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_130), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_187), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_87), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_38), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_185), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_184), .Y(n_314) );
XOR2xp5_ASAP7_75t_L g315 ( .A(n_156), .B(n_151), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_143), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_103), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_149), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_109), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_125), .Y(n_320) );
NOR2xp67_ASAP7_75t_L g321 ( .A(n_212), .B(n_120), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_13), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_127), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_121), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_56), .Y(n_325) );
BUFx2_ASAP7_75t_SL g326 ( .A(n_24), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_129), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_131), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_67), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_64), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_126), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_140), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_90), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_97), .Y(n_334) );
NOR2xp67_ASAP7_75t_L g335 ( .A(n_147), .B(n_178), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_243), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_243), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_268), .B(n_0), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_243), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_222), .B(n_1), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_243), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_320), .B(n_2), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_323), .B(n_2), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_243), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_218), .B(n_3), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_223), .B(n_4), .Y(n_346) );
AOI22xp5_ASAP7_75t_L g347 ( .A1(n_255), .A2(n_7), .B1(n_5), .B2(n_6), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_243), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_243), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_222), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_252), .B(n_5), .Y(n_351) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_265), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_220), .A2(n_10), .B1(n_8), .B2(n_9), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_230), .B(n_11), .Y(n_354) );
INVx4_ASAP7_75t_L g355 ( .A(n_265), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_281), .Y(n_356) );
AND2x6_ASAP7_75t_L g357 ( .A(n_281), .B(n_112), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_219), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_284), .B(n_11), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_284), .B(n_12), .Y(n_360) );
CKINVDCx11_ASAP7_75t_R g361 ( .A(n_226), .Y(n_361) );
CKINVDCx16_ASAP7_75t_R g362 ( .A(n_236), .Y(n_362) );
INVxp67_ASAP7_75t_L g363 ( .A(n_274), .Y(n_363) );
OA21x2_ASAP7_75t_L g364 ( .A1(n_219), .A2(n_114), .B(n_113), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_225), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_225), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_262), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_221), .B(n_14), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_249), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_270), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_262), .Y(n_371) );
BUFx8_ASAP7_75t_SL g372 ( .A(n_258), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_303), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_270), .Y(n_374) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_364), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g376 ( .A(n_363), .B(n_250), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_345), .A2(n_238), .B1(n_241), .B2(n_220), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_363), .B(n_259), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_336), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_355), .B(n_263), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_337), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_350), .B(n_263), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_373), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_340), .A2(n_246), .B1(n_251), .B2(n_240), .Y(n_384) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_340), .B(n_272), .Y(n_385) );
NAND2xp33_ASAP7_75t_L g386 ( .A(n_357), .B(n_216), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_336), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_336), .Y(n_388) );
INVx1_ASAP7_75t_SL g389 ( .A(n_359), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_337), .Y(n_390) );
INVx3_ASAP7_75t_L g391 ( .A(n_340), .Y(n_391) );
BUFx6f_ASAP7_75t_SL g392 ( .A(n_340), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_344), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_339), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_344), .Y(n_395) );
CKINVDCx14_ASAP7_75t_R g396 ( .A(n_369), .Y(n_396) );
INVx4_ASAP7_75t_L g397 ( .A(n_357), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_344), .Y(n_398) );
AND3x2_ASAP7_75t_L g399 ( .A(n_359), .B(n_247), .C(n_228), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_352), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_352), .Y(n_401) );
INVx2_ASAP7_75t_SL g402 ( .A(n_373), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_341), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_341), .Y(n_404) );
INVx4_ASAP7_75t_L g405 ( .A(n_357), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_348), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_350), .B(n_272), .Y(n_407) );
AND2x2_ASAP7_75t_SL g408 ( .A(n_351), .B(n_302), .Y(n_408) );
INVx3_ASAP7_75t_L g409 ( .A(n_351), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_348), .B(n_300), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_372), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_349), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_349), .B(n_300), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_378), .B(n_362), .Y(n_414) );
INVxp67_ASAP7_75t_L g415 ( .A(n_378), .Y(n_415) );
NAND2x1p5_ASAP7_75t_L g416 ( .A(n_408), .B(n_360), .Y(n_416) );
OAI21xp5_ASAP7_75t_L g417 ( .A1(n_381), .A2(n_364), .B(n_368), .Y(n_417) );
BUFx3_ASAP7_75t_L g418 ( .A(n_378), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_376), .B(n_362), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_389), .B(n_345), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_391), .B(n_360), .Y(n_421) );
INVx2_ASAP7_75t_SL g422 ( .A(n_408), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_411), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_391), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_384), .A2(n_342), .B1(n_343), .B2(n_338), .Y(n_425) );
NAND3xp33_ASAP7_75t_L g426 ( .A(n_384), .B(n_343), .C(n_347), .Y(n_426) );
AND2x6_ASAP7_75t_SL g427 ( .A(n_396), .B(n_361), .Y(n_427) );
AND2x2_ASAP7_75t_SL g428 ( .A(n_377), .B(n_347), .Y(n_428) );
O2A1O1Ixp33_ASAP7_75t_L g429 ( .A1(n_385), .A2(n_353), .B(n_354), .C(n_346), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_391), .Y(n_430) );
BUFx3_ASAP7_75t_L g431 ( .A(n_383), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_377), .B(n_227), .Y(n_432) );
INVx2_ASAP7_75t_SL g433 ( .A(n_399), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_397), .B(n_217), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_399), .B(n_409), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_409), .B(n_224), .Y(n_436) );
AND2x6_ASAP7_75t_L g437 ( .A(n_392), .B(n_303), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_392), .A2(n_353), .B1(n_241), .B2(n_257), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_402), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_390), .B(n_357), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_390), .B(n_357), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_394), .B(n_357), .Y(n_442) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_397), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_403), .B(n_235), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_382), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_382), .Y(n_446) );
INVx4_ASAP7_75t_L g447 ( .A(n_405), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_407), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_410), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_380), .B(n_231), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_380), .A2(n_266), .B1(n_257), .B2(n_233), .Y(n_451) );
INVx4_ASAP7_75t_L g452 ( .A(n_405), .Y(n_452) );
NOR3x1_ASAP7_75t_L g453 ( .A(n_410), .B(n_244), .C(n_226), .Y(n_453) );
BUFx8_ASAP7_75t_L g454 ( .A(n_375), .Y(n_454) );
NAND3xp33_ASAP7_75t_SL g455 ( .A(n_413), .B(n_266), .C(n_248), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_404), .B(n_310), .Y(n_456) );
NOR2xp67_ASAP7_75t_L g457 ( .A(n_400), .B(n_358), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_406), .B(n_313), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_412), .Y(n_459) );
AOI221xp5_ASAP7_75t_L g460 ( .A1(n_412), .A2(n_232), .B1(n_317), .B2(n_311), .C(n_233), .Y(n_460) );
AND2x6_ASAP7_75t_SL g461 ( .A(n_386), .B(n_278), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_379), .B(n_313), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_387), .B(n_324), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_387), .B(n_232), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_375), .A2(n_317), .B1(n_325), .B2(n_311), .Y(n_465) );
NOR2x1p5_ASAP7_75t_L g466 ( .A(n_375), .B(n_325), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_375), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g468 ( .A(n_455), .B(n_288), .C(n_329), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_445), .B(n_330), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_446), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_440), .A2(n_393), .B(n_388), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_415), .B(n_244), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_435), .B(n_291), .Y(n_473) );
BUFx2_ASAP7_75t_L g474 ( .A(n_416), .Y(n_474) );
OAI21xp5_ASAP7_75t_L g475 ( .A1(n_417), .A2(n_398), .B(n_395), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_441), .A2(n_398), .B(n_364), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_420), .A2(n_315), .B1(n_248), .B2(n_285), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_429), .A2(n_301), .B(n_307), .C(n_297), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_464), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_424), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_442), .A2(n_364), .B(n_400), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_442), .A2(n_364), .B(n_401), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_459), .A2(n_365), .B(n_366), .C(n_358), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_419), .B(n_267), .Y(n_484) );
AND2x4_ASAP7_75t_L g485 ( .A(n_435), .B(n_422), .Y(n_485) );
OR2x6_ASAP7_75t_L g486 ( .A(n_414), .B(n_326), .Y(n_486) );
NAND3xp33_ASAP7_75t_L g487 ( .A(n_425), .B(n_426), .C(n_465), .Y(n_487) );
AOI221xp5_ASAP7_75t_L g488 ( .A1(n_432), .A2(n_308), .B1(n_319), .B2(n_322), .C(n_312), .Y(n_488) );
BUFx3_ASAP7_75t_L g489 ( .A(n_423), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_430), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_433), .B(n_276), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_444), .B(n_277), .Y(n_492) );
OAI21xp33_ASAP7_75t_L g493 ( .A1(n_460), .A2(n_304), .B(n_293), .Y(n_493) );
AO32x2_ASAP7_75t_L g494 ( .A1(n_466), .A2(n_356), .A3(n_358), .B1(n_366), .B2(n_365), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_428), .A2(n_334), .B1(n_333), .B2(n_234), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_421), .A2(n_287), .B1(n_283), .B2(n_366), .Y(n_496) );
NAND2x1p5_ASAP7_75t_L g497 ( .A(n_431), .B(n_370), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_421), .A2(n_237), .B(n_229), .Y(n_498) );
INVx4_ASAP7_75t_L g499 ( .A(n_437), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_436), .A2(n_245), .B(n_242), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_458), .A2(n_371), .B1(n_367), .B2(n_374), .Y(n_501) );
INVxp67_ASAP7_75t_L g502 ( .A(n_458), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_450), .B(n_374), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_456), .B(n_367), .Y(n_504) );
OR2x6_ASAP7_75t_SL g505 ( .A(n_427), .B(n_453), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_462), .A2(n_371), .B1(n_254), .B2(n_256), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_463), .B(n_15), .Y(n_507) );
AOI33xp33_ASAP7_75t_L g508 ( .A1(n_449), .A2(n_282), .A3(n_253), .B1(n_260), .B2(n_261), .B3(n_264), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_434), .A2(n_271), .B(n_269), .Y(n_509) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_443), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_461), .B(n_239), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_457), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_439), .A2(n_280), .B(n_279), .Y(n_513) );
NAND2x1p5_ASAP7_75t_L g514 ( .A(n_447), .B(n_275), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_454), .B(n_273), .Y(n_515) );
AOI33xp33_ASAP7_75t_L g516 ( .A1(n_452), .A2(n_289), .A3(n_328), .B1(n_327), .B2(n_294), .B3(n_295), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_443), .A2(n_298), .B1(n_299), .B2(n_296), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_448), .A2(n_314), .B1(n_316), .B2(n_305), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_432), .B(n_16), .Y(n_519) );
AOI21xp33_ASAP7_75t_L g520 ( .A1(n_419), .A2(n_292), .B(n_290), .Y(n_520) );
OAI21x1_ASAP7_75t_L g521 ( .A1(n_417), .A2(n_318), .B(n_309), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_448), .Y(n_522) );
BUFx2_ASAP7_75t_L g523 ( .A(n_418), .Y(n_523) );
INVx1_ASAP7_75t_SL g524 ( .A(n_448), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_448), .B(n_306), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_459), .Y(n_526) );
AO32x2_ASAP7_75t_L g527 ( .A1(n_467), .A2(n_356), .A3(n_335), .B1(n_321), .B2(n_286), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_448), .B(n_332), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_448), .A2(n_331), .B1(n_356), .B2(n_18), .Y(n_529) );
OAI21xp33_ASAP7_75t_SL g530 ( .A1(n_445), .A2(n_331), .B(n_17), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_415), .A2(n_20), .B1(n_18), .B2(n_19), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_448), .A2(n_22), .B1(n_20), .B2(n_21), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_427), .Y(n_533) );
O2A1O1Ixp5_ASAP7_75t_SL g534 ( .A1(n_417), .A2(n_117), .B(n_118), .C(n_116), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_415), .B(n_21), .Y(n_535) );
INVxp67_ASAP7_75t_SL g536 ( .A(n_477), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_524), .B(n_23), .Y(n_537) );
AO32x2_ASAP7_75t_L g538 ( .A1(n_529), .A2(n_496), .A3(n_532), .B1(n_501), .B2(n_506), .Y(n_538) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_530), .A2(n_478), .B(n_502), .C(n_479), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_524), .B(n_26), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_470), .A2(n_29), .B1(n_27), .B2(n_28), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_522), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_528), .A2(n_31), .B1(n_28), .B2(n_30), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_523), .Y(n_544) );
AOI211x1_ASAP7_75t_L g545 ( .A1(n_487), .A2(n_34), .B(n_30), .C(n_33), .Y(n_545) );
AO31x2_ASAP7_75t_L g546 ( .A1(n_483), .A2(n_37), .A3(n_35), .B(n_36), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_484), .B(n_35), .Y(n_547) );
O2A1O1Ixp33_ASAP7_75t_L g548 ( .A1(n_503), .A2(n_39), .B(n_36), .C(n_37), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_526), .Y(n_549) );
AOI21xp33_ASAP7_75t_L g550 ( .A1(n_491), .A2(n_40), .B(n_41), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_472), .A2(n_43), .B1(n_41), .B2(n_42), .Y(n_551) );
AOI221x1_ASAP7_75t_L g552 ( .A1(n_487), .A2(n_42), .B1(n_44), .B2(n_45), .C(n_46), .Y(n_552) );
NAND3x1_ASAP7_75t_L g553 ( .A(n_505), .B(n_45), .C(n_47), .Y(n_553) );
INVxp67_ASAP7_75t_SL g554 ( .A(n_497), .Y(n_554) );
O2A1O1Ixp33_ASAP7_75t_L g555 ( .A1(n_519), .A2(n_48), .B(n_49), .C(n_50), .Y(n_555) );
INVx5_ASAP7_75t_SL g556 ( .A(n_486), .Y(n_556) );
NAND3xp33_ASAP7_75t_L g557 ( .A(n_520), .B(n_50), .C(n_52), .Y(n_557) );
NOR2x1_ASAP7_75t_R g558 ( .A(n_533), .B(n_52), .Y(n_558) );
INVx4_ASAP7_75t_L g559 ( .A(n_510), .Y(n_559) );
AO32x2_ASAP7_75t_L g560 ( .A1(n_517), .A2(n_53), .A3(n_54), .B1(n_56), .B2(n_57), .Y(n_560) );
AOI31xp67_ASAP7_75t_L g561 ( .A1(n_534), .A2(n_162), .A3(n_213), .B(n_211), .Y(n_561) );
BUFx3_ASAP7_75t_L g562 ( .A(n_486), .Y(n_562) );
BUFx3_ASAP7_75t_L g563 ( .A(n_497), .Y(n_563) );
O2A1O1Ixp33_ASAP7_75t_L g564 ( .A1(n_469), .A2(n_58), .B(n_59), .C(n_60), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_485), .B(n_61), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_480), .Y(n_566) );
OAI22x1_ASAP7_75t_L g567 ( .A1(n_495), .A2(n_62), .B1(n_63), .B2(n_64), .Y(n_567) );
AOI221x1_ASAP7_75t_L g568 ( .A1(n_468), .A2(n_65), .B1(n_66), .B2(n_67), .C(n_68), .Y(n_568) );
BUFx2_ASAP7_75t_L g569 ( .A(n_474), .Y(n_569) );
OR2x6_ASAP7_75t_L g570 ( .A(n_485), .B(n_68), .Y(n_570) );
AOI21xp33_ASAP7_75t_L g571 ( .A1(n_535), .A2(n_69), .B(n_70), .Y(n_571) );
A2O1A1Ixp33_ASAP7_75t_L g572 ( .A1(n_498), .A2(n_71), .B(n_72), .C(n_73), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_473), .B(n_71), .Y(n_573) );
AO31x2_ASAP7_75t_L g574 ( .A1(n_504), .A2(n_73), .A3(n_74), .B(n_75), .Y(n_574) );
AO31x2_ASAP7_75t_L g575 ( .A1(n_500), .A2(n_74), .A3(n_75), .B(n_76), .Y(n_575) );
BUFx2_ASAP7_75t_R g576 ( .A(n_515), .Y(n_576) );
AOI221xp5_ASAP7_75t_L g577 ( .A1(n_511), .A2(n_78), .B1(n_79), .B2(n_81), .C(n_82), .Y(n_577) );
NAND2xp33_ASAP7_75t_SL g578 ( .A(n_499), .B(n_83), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_490), .Y(n_579) );
AOI211x1_ASAP7_75t_L g580 ( .A1(n_492), .A2(n_84), .B(n_85), .C(n_86), .Y(n_580) );
AO32x2_ASAP7_75t_L g581 ( .A1(n_518), .A2(n_84), .A3(n_85), .B1(n_86), .B2(n_87), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_531), .Y(n_582) );
AO31x2_ASAP7_75t_L g583 ( .A1(n_527), .A2(n_88), .A3(n_89), .B(n_90), .Y(n_583) );
AO31x2_ASAP7_75t_L g584 ( .A1(n_527), .A2(n_91), .A3(n_92), .B(n_95), .Y(n_584) );
BUFx12f_ASAP7_75t_L g585 ( .A(n_514), .Y(n_585) );
NAND3xp33_ASAP7_75t_SL g586 ( .A(n_516), .B(n_98), .C(n_99), .Y(n_586) );
BUFx10_ASAP7_75t_L g587 ( .A(n_512), .Y(n_587) );
INVx3_ASAP7_75t_L g588 ( .A(n_514), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_525), .A2(n_99), .B1(n_100), .B2(n_101), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_493), .A2(n_100), .B1(n_101), .B2(n_102), .Y(n_590) );
AO31x2_ASAP7_75t_L g591 ( .A1(n_527), .A2(n_104), .A3(n_105), .B(n_106), .Y(n_591) );
NOR4xp25_ASAP7_75t_L g592 ( .A(n_508), .B(n_104), .C(n_105), .D(n_106), .Y(n_592) );
A2O1A1Ixp33_ASAP7_75t_L g593 ( .A1(n_507), .A2(n_107), .B(n_108), .C(n_109), .Y(n_593) );
AO31x2_ASAP7_75t_L g594 ( .A1(n_513), .A2(n_108), .A3(n_110), .B(n_148), .Y(n_594) );
OAI21x1_ASAP7_75t_L g595 ( .A1(n_509), .A2(n_153), .B(n_155), .Y(n_595) );
AO31x2_ASAP7_75t_L g596 ( .A1(n_494), .A2(n_170), .A3(n_171), .B(n_172), .Y(n_596) );
AO31x2_ASAP7_75t_L g597 ( .A1(n_494), .A2(n_180), .A3(n_181), .B(n_182), .Y(n_597) );
CKINVDCx16_ASAP7_75t_R g598 ( .A(n_494), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_470), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_524), .Y(n_600) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_488), .A2(n_188), .B1(n_189), .B2(n_190), .C(n_194), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_524), .Y(n_602) );
OAI21xp5_ASAP7_75t_L g603 ( .A1(n_521), .A2(n_195), .B(n_196), .Y(n_603) );
AOI21xp5_ASAP7_75t_SL g604 ( .A1(n_499), .A2(n_214), .B(n_201), .Y(n_604) );
AO31x2_ASAP7_75t_L g605 ( .A1(n_476), .A2(n_197), .A3(n_203), .B(n_204), .Y(n_605) );
O2A1O1Ixp33_ASAP7_75t_L g606 ( .A1(n_530), .A2(n_478), .B(n_415), .C(n_502), .Y(n_606) );
AO31x2_ASAP7_75t_L g607 ( .A1(n_476), .A2(n_483), .A3(n_481), .B(n_482), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_524), .B(n_448), .Y(n_608) );
BUFx3_ASAP7_75t_L g609 ( .A(n_489), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_524), .Y(n_610) );
OAI21xp5_ASAP7_75t_L g611 ( .A1(n_521), .A2(n_475), .B(n_471), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_524), .B(n_378), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_536), .B(n_582), .Y(n_613) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_554), .Y(n_614) );
A2O1A1Ixp33_ASAP7_75t_L g615 ( .A1(n_555), .A2(n_548), .B(n_564), .C(n_578), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_602), .B(n_610), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_607), .Y(n_617) );
INVx6_ASAP7_75t_L g618 ( .A(n_609), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_607), .Y(n_619) );
A2O1A1Ixp33_ASAP7_75t_L g620 ( .A1(n_601), .A2(n_593), .B(n_572), .C(n_547), .Y(n_620) );
OA21x2_ASAP7_75t_L g621 ( .A1(n_552), .A2(n_568), .B(n_595), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_549), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_544), .B(n_569), .Y(n_623) );
AO31x2_ASAP7_75t_L g624 ( .A1(n_567), .A2(n_543), .A3(n_541), .B(n_579), .Y(n_624) );
BUFx8_ASAP7_75t_L g625 ( .A(n_585), .Y(n_625) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_565), .Y(n_626) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_565), .Y(n_627) );
INVx3_ASAP7_75t_L g628 ( .A(n_559), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_570), .B(n_573), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_566), .Y(n_630) );
INVx8_ASAP7_75t_L g631 ( .A(n_570), .Y(n_631) );
AO21x2_ASAP7_75t_L g632 ( .A1(n_592), .A2(n_571), .B(n_557), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_537), .Y(n_633) );
OAI21x1_ASAP7_75t_L g634 ( .A1(n_604), .A2(n_588), .B(n_540), .Y(n_634) );
OA21x2_ASAP7_75t_L g635 ( .A1(n_590), .A2(n_550), .B(n_589), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_551), .Y(n_636) );
OA21x2_ASAP7_75t_L g637 ( .A1(n_561), .A2(n_605), .B(n_598), .Y(n_637) );
OA21x2_ASAP7_75t_L g638 ( .A1(n_577), .A2(n_596), .B(n_597), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_562), .B(n_576), .Y(n_639) );
AO21x2_ASAP7_75t_L g640 ( .A1(n_583), .A2(n_591), .B(n_584), .Y(n_640) );
OA21x2_ASAP7_75t_L g641 ( .A1(n_545), .A2(n_591), .B(n_584), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_556), .B(n_580), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_574), .Y(n_643) );
OR2x6_ASAP7_75t_L g644 ( .A(n_553), .B(n_558), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_574), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_574), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_581), .B(n_560), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_587), .B(n_538), .Y(n_648) );
INVx3_ASAP7_75t_L g649 ( .A(n_575), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_581), .Y(n_650) );
AND2x4_ASAP7_75t_L g651 ( .A(n_546), .B(n_594), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_560), .Y(n_652) );
AO21x2_ASAP7_75t_L g653 ( .A1(n_583), .A2(n_584), .B(n_591), .Y(n_653) );
NOR2xp33_ASAP7_75t_SL g654 ( .A(n_538), .B(n_594), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_542), .Y(n_655) );
NOR2x1_ASAP7_75t_SL g656 ( .A(n_570), .B(n_499), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_608), .B(n_524), .Y(n_657) );
OA21x2_ASAP7_75t_L g658 ( .A1(n_611), .A2(n_521), .B(n_603), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_612), .B(n_524), .Y(n_659) );
AOI21xp33_ASAP7_75t_L g660 ( .A1(n_606), .A2(n_539), .B(n_478), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_608), .A2(n_438), .B1(n_377), .B2(n_451), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_608), .B(n_524), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_582), .A2(n_428), .B1(n_586), .B2(n_536), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_608), .B(n_524), .Y(n_664) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_600), .Y(n_665) );
AO21x2_ASAP7_75t_L g666 ( .A1(n_611), .A2(n_603), .B(n_521), .Y(n_666) );
AND2x4_ASAP7_75t_L g667 ( .A(n_563), .B(n_554), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_536), .B(n_415), .Y(n_668) );
AO21x2_ASAP7_75t_L g669 ( .A1(n_611), .A2(n_603), .B(n_521), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_599), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_608), .B(n_524), .Y(n_671) );
O2A1O1Ixp33_ASAP7_75t_L g672 ( .A1(n_539), .A2(n_606), .B(n_593), .C(n_572), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_536), .B(n_415), .Y(n_673) );
AND2x4_ASAP7_75t_L g674 ( .A(n_563), .B(n_554), .Y(n_674) );
BUFx3_ASAP7_75t_L g675 ( .A(n_563), .Y(n_675) );
AO21x2_ASAP7_75t_L g676 ( .A1(n_611), .A2(n_603), .B(n_521), .Y(n_676) );
OA21x2_ASAP7_75t_L g677 ( .A1(n_611), .A2(n_521), .B(n_603), .Y(n_677) );
AND2x4_ASAP7_75t_L g678 ( .A(n_563), .B(n_554), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_608), .A2(n_438), .B1(n_377), .B2(n_451), .Y(n_679) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_600), .Y(n_680) );
AO21x2_ASAP7_75t_L g681 ( .A1(n_611), .A2(n_603), .B(n_521), .Y(n_681) );
BUFx3_ASAP7_75t_L g682 ( .A(n_563), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_613), .A2(n_679), .B1(n_661), .B2(n_673), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_617), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_619), .Y(n_685) );
BUFx3_ASAP7_75t_L g686 ( .A(n_625), .Y(n_686) );
INVxp67_ASAP7_75t_L g687 ( .A(n_625), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_655), .Y(n_688) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_614), .Y(n_689) );
BUFx2_ASAP7_75t_L g690 ( .A(n_614), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_616), .Y(n_691) );
OR2x2_ASAP7_75t_L g692 ( .A(n_657), .B(n_662), .Y(n_692) );
OR2x6_ASAP7_75t_L g693 ( .A(n_631), .B(n_626), .Y(n_693) );
OR2x6_ASAP7_75t_L g694 ( .A(n_631), .B(n_627), .Y(n_694) );
OR2x2_ASAP7_75t_L g695 ( .A(n_664), .B(n_671), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_670), .B(n_630), .Y(n_696) );
AO21x2_ASAP7_75t_L g697 ( .A1(n_643), .A2(n_646), .B(n_645), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_659), .B(n_622), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_636), .B(n_663), .Y(n_699) );
OR2x2_ASAP7_75t_L g700 ( .A(n_665), .B(n_680), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_647), .B(n_651), .Y(n_701) );
OR2x6_ASAP7_75t_L g702 ( .A(n_667), .B(n_674), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_651), .B(n_665), .Y(n_703) );
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_656), .A2(n_644), .B1(n_629), .B2(n_642), .Y(n_704) );
INVxp67_ASAP7_75t_L g705 ( .A(n_623), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_678), .B(n_641), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_668), .B(n_673), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_641), .B(n_633), .Y(n_708) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_675), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_641), .B(n_668), .Y(n_710) );
OR2x2_ASAP7_75t_L g711 ( .A(n_650), .B(n_652), .Y(n_711) );
OR2x2_ASAP7_75t_L g712 ( .A(n_648), .B(n_649), .Y(n_712) );
OR2x2_ASAP7_75t_L g713 ( .A(n_648), .B(n_649), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_624), .B(n_660), .Y(n_714) );
BUFx6f_ASAP7_75t_L g715 ( .A(n_682), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_640), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_653), .Y(n_717) );
OR2x6_ASAP7_75t_L g718 ( .A(n_672), .B(n_628), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_653), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_624), .B(n_654), .Y(n_720) );
OR2x2_ASAP7_75t_L g721 ( .A(n_632), .B(n_637), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_684), .Y(n_722) );
OR2x2_ASAP7_75t_L g723 ( .A(n_690), .B(n_703), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_701), .B(n_637), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_710), .B(n_638), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_710), .B(n_708), .Y(n_726) );
AND2x4_ASAP7_75t_L g727 ( .A(n_706), .B(n_634), .Y(n_727) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_689), .Y(n_728) );
AND2x4_ASAP7_75t_L g729 ( .A(n_706), .B(n_681), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_708), .B(n_638), .Y(n_730) );
AND2x2_ASAP7_75t_L g731 ( .A(n_714), .B(n_699), .Y(n_731) );
BUFx4f_ASAP7_75t_L g732 ( .A(n_702), .Y(n_732) );
AOI33xp33_ASAP7_75t_L g733 ( .A1(n_704), .A2(n_639), .A3(n_618), .B1(n_621), .B2(n_615), .B3(n_620), .Y(n_733) );
OR2x2_ASAP7_75t_L g734 ( .A(n_700), .B(n_669), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_688), .Y(n_735) );
OR2x2_ASAP7_75t_L g736 ( .A(n_700), .B(n_669), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_698), .B(n_666), .Y(n_737) );
OR2x2_ASAP7_75t_L g738 ( .A(n_692), .B(n_676), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_696), .B(n_677), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_695), .B(n_635), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_691), .Y(n_741) );
OR2x2_ASAP7_75t_L g742 ( .A(n_695), .B(n_621), .Y(n_742) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_709), .Y(n_743) );
INVxp67_ASAP7_75t_SL g744 ( .A(n_685), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_683), .B(n_635), .Y(n_745) );
INVxp67_ASAP7_75t_L g746 ( .A(n_686), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_711), .Y(n_747) );
AND2x2_ASAP7_75t_L g748 ( .A(n_720), .B(n_658), .Y(n_748) );
INVxp67_ASAP7_75t_SL g749 ( .A(n_744), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_746), .B(n_687), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_726), .B(n_712), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_747), .B(n_737), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_737), .B(n_711), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_731), .B(n_724), .Y(n_754) );
AND2x4_ASAP7_75t_L g755 ( .A(n_727), .B(n_716), .Y(n_755) );
AND2x4_ASAP7_75t_L g756 ( .A(n_727), .B(n_716), .Y(n_756) );
AND2x2_ASAP7_75t_L g757 ( .A(n_731), .B(n_713), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_725), .B(n_697), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_725), .B(n_697), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_739), .B(n_697), .Y(n_760) );
AND2x4_ASAP7_75t_L g761 ( .A(n_727), .B(n_717), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_730), .B(n_719), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_740), .B(n_718), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_722), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_742), .Y(n_765) );
INVxp67_ASAP7_75t_L g766 ( .A(n_743), .Y(n_766) );
OR2x2_ASAP7_75t_L g767 ( .A(n_723), .B(n_721), .Y(n_767) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_728), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_738), .Y(n_769) );
INVx4_ASAP7_75t_L g770 ( .A(n_732), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_738), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_768), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_764), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_766), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_752), .Y(n_775) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_749), .Y(n_776) );
AND2x2_ASAP7_75t_L g777 ( .A(n_754), .B(n_748), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_757), .B(n_741), .Y(n_778) );
OR2x2_ASAP7_75t_L g779 ( .A(n_751), .B(n_734), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_767), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_767), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_758), .B(n_729), .Y(n_782) );
OR2x2_ASAP7_75t_L g783 ( .A(n_753), .B(n_736), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_765), .Y(n_784) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_749), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_759), .B(n_735), .Y(n_786) );
NAND4xp25_ASAP7_75t_L g787 ( .A(n_750), .B(n_733), .C(n_707), .D(n_745), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_772), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_775), .B(n_760), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_780), .B(n_769), .Y(n_790) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_776), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_784), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_777), .B(n_762), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_781), .B(n_771), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_786), .B(n_774), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_787), .B(n_705), .Y(n_796) );
INVxp67_ASAP7_75t_L g797 ( .A(n_785), .Y(n_797) );
INVx2_ASAP7_75t_L g798 ( .A(n_773), .Y(n_798) );
OR2x2_ASAP7_75t_L g799 ( .A(n_779), .B(n_763), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_791), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_793), .B(n_782), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_796), .B(n_778), .Y(n_802) );
OR2x2_ASAP7_75t_L g803 ( .A(n_789), .B(n_783), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_798), .Y(n_804) );
BUFx2_ASAP7_75t_L g805 ( .A(n_797), .Y(n_805) );
AOI222xp33_ASAP7_75t_L g806 ( .A1(n_802), .A2(n_795), .B1(n_790), .B2(n_794), .C1(n_788), .C2(n_792), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_801), .B(n_805), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_800), .B(n_799), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_806), .B(n_807), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_809), .Y(n_810) );
OR2x2_ASAP7_75t_L g811 ( .A(n_810), .B(n_808), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_811), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g813 ( .A1(n_812), .A2(n_803), .B1(n_770), .B2(n_804), .Y(n_813) );
XNOR2x1_ASAP7_75t_L g814 ( .A(n_813), .B(n_693), .Y(n_814) );
OAI21xp5_ASAP7_75t_L g815 ( .A1(n_814), .A2(n_694), .B(n_693), .Y(n_815) );
OR2x2_ASAP7_75t_L g816 ( .A(n_815), .B(n_693), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g817 ( .A1(n_816), .A2(n_694), .B(n_715), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_817), .A2(n_756), .B1(n_755), .B2(n_761), .Y(n_818) );
endmodule