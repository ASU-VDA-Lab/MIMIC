module fake_netlist_1_10065_n_644 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_644);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_644;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g85 ( .A(n_84), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_54), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_70), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_77), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_62), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_51), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_61), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_56), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_17), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_74), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_17), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_41), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_52), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_65), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_60), .Y(n_99) );
HB1xp67_ASAP7_75t_L g100 ( .A(n_59), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_63), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_14), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_55), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_7), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_81), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_11), .Y(n_106) );
BUFx5_ASAP7_75t_L g107 ( .A(n_58), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_27), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_14), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_21), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_76), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_22), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_75), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_80), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_9), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_50), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_47), .Y(n_117) );
BUFx3_ASAP7_75t_L g118 ( .A(n_38), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_19), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_4), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_4), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_48), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_71), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_100), .B(n_0), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_85), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_106), .B(n_0), .Y(n_126) );
AND2x2_ASAP7_75t_SL g127 ( .A(n_87), .B(n_83), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_86), .Y(n_128) );
INVxp33_ASAP7_75t_SL g129 ( .A(n_106), .Y(n_129) );
NOR2x1_ASAP7_75t_L g130 ( .A(n_102), .B(n_33), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_88), .Y(n_131) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_87), .A2(n_32), .B(n_79), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_109), .B(n_1), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_89), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_91), .Y(n_135) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_94), .A2(n_31), .B(n_78), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_96), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_97), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_115), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_94), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_98), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_99), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_103), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_105), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_108), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_110), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_107), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_113), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_116), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_118), .B(n_1), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_118), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_117), .Y(n_152) );
BUFx2_ASAP7_75t_L g153 ( .A(n_150), .Y(n_153) );
BUFx10_ASAP7_75t_L g154 ( .A(n_150), .Y(n_154) );
INVx5_ASAP7_75t_L g155 ( .A(n_150), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_129), .B(n_123), .Y(n_156) );
INVxp67_ASAP7_75t_SL g157 ( .A(n_126), .Y(n_157) );
OR2x6_ASAP7_75t_L g158 ( .A(n_124), .B(n_121), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_147), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_125), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_147), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_125), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_140), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_127), .B(n_114), .Y(n_164) );
INVx4_ASAP7_75t_L g165 ( .A(n_150), .Y(n_165) );
BUFx3_ASAP7_75t_L g166 ( .A(n_151), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_127), .B(n_114), .Y(n_167) );
INVx1_ASAP7_75t_SL g168 ( .A(n_151), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_128), .B(n_123), .Y(n_169) );
HB1xp67_ASAP7_75t_L g170 ( .A(n_128), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_125), .Y(n_171) );
INVx2_ASAP7_75t_SL g172 ( .A(n_127), .Y(n_172) );
NAND3xp33_ASAP7_75t_L g173 ( .A(n_131), .B(n_122), .C(n_120), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_132), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_131), .B(n_119), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_134), .B(n_90), .Y(n_176) );
INVx4_ASAP7_75t_L g177 ( .A(n_132), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_133), .A2(n_104), .B1(n_93), .B2(n_95), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_134), .Y(n_179) );
OAI21xp33_ASAP7_75t_SL g180 ( .A1(n_135), .A2(n_152), .B(n_149), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_125), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_135), .A2(n_119), .B1(n_90), .B2(n_92), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_140), .Y(n_183) );
INVx5_ASAP7_75t_L g184 ( .A(n_125), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_140), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_140), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_125), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_170), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_157), .B(n_137), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_169), .B(n_137), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_183), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_159), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_176), .B(n_138), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_163), .Y(n_194) );
INVx5_ASAP7_75t_L g195 ( .A(n_154), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_163), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_185), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_179), .B(n_138), .Y(n_198) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_158), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_179), .B(n_141), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_180), .A2(n_152), .B(n_149), .C(n_148), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_175), .B(n_148), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_158), .B(n_165), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_168), .B(n_146), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_154), .B(n_92), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_153), .A2(n_132), .B(n_136), .Y(n_206) );
INVx4_ASAP7_75t_L g207 ( .A(n_165), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_159), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_172), .A2(n_146), .B1(n_145), .B2(n_144), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_158), .B(n_145), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_158), .B(n_144), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_161), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_153), .A2(n_136), .B(n_132), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_158), .B(n_165), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_183), .Y(n_215) );
NAND2x1p5_ASAP7_75t_L g216 ( .A(n_165), .B(n_136), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_178), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_154), .B(n_139), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_182), .B(n_143), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_172), .A2(n_143), .B1(n_142), .B2(n_141), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_155), .B(n_142), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_185), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_155), .B(n_139), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_156), .B(n_139), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_161), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_186), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_155), .B(n_112), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_154), .B(n_101), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_155), .B(n_111), .Y(n_229) );
OR2x2_ASAP7_75t_L g230 ( .A(n_178), .B(n_2), .Y(n_230) );
AO22x1_ASAP7_75t_L g231 ( .A1(n_155), .A2(n_130), .B1(n_85), .B2(n_136), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_155), .B(n_107), .Y(n_232) );
AOI21x1_ASAP7_75t_L g233 ( .A1(n_231), .A2(n_164), .B(n_167), .Y(n_233) );
NAND3xp33_ASAP7_75t_L g234 ( .A(n_209), .B(n_180), .C(n_173), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_230), .B(n_93), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_195), .Y(n_236) );
BUFx2_ASAP7_75t_L g237 ( .A(n_203), .Y(n_237) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_195), .Y(n_238) );
AO22x1_ASAP7_75t_L g239 ( .A1(n_217), .A2(n_95), .B1(n_174), .B2(n_177), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_195), .B(n_166), .Y(n_240) );
INVx3_ASAP7_75t_SL g241 ( .A(n_230), .Y(n_241) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_206), .A2(n_183), .B(n_186), .Y(n_242) );
BUFx2_ASAP7_75t_L g243 ( .A(n_203), .Y(n_243) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_213), .A2(n_173), .B(n_174), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_203), .A2(n_177), .B1(n_174), .B2(n_166), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_201), .A2(n_183), .B(n_166), .C(n_85), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_214), .B(n_174), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_212), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_190), .A2(n_85), .B(n_177), .C(n_181), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_189), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_188), .B(n_177), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_195), .Y(n_252) );
CKINVDCx8_ASAP7_75t_R g253 ( .A(n_217), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_214), .B(n_107), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g255 ( .A1(n_219), .A2(n_187), .B(n_181), .C(n_171), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_214), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_199), .B(n_2), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_193), .A2(n_187), .B(n_171), .C(n_162), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_195), .B(n_107), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_210), .B(n_107), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_218), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_207), .B(n_107), .Y(n_262) );
NOR2xp67_ASAP7_75t_L g263 ( .A(n_224), .B(n_3), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g264 ( .A1(n_220), .A2(n_184), .B1(n_162), .B2(n_6), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_211), .B(n_107), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_207), .B(n_184), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_212), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_218), .A2(n_184), .B1(n_160), .B2(n_6), .Y(n_268) );
NOR2xp33_ASAP7_75t_R g269 ( .A(n_207), .B(n_3), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_231), .A2(n_184), .B(n_160), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_198), .A2(n_200), .B(n_202), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_204), .B(n_5), .Y(n_272) );
OAI22x1_ASAP7_75t_L g273 ( .A1(n_216), .A2(n_5), .B1(n_7), .B2(n_8), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_225), .B(n_8), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_194), .A2(n_184), .B(n_160), .C(n_11), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_225), .B(n_9), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_251), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_250), .B(n_215), .Y(n_278) );
AO21x1_ASAP7_75t_L g279 ( .A1(n_264), .A2(n_216), .B(n_232), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_271), .A2(n_216), .B(n_223), .Y(n_280) );
OAI22xp33_ASAP7_75t_L g281 ( .A1(n_241), .A2(n_194), .B1(n_196), .B2(n_226), .Y(n_281) );
O2A1O1Ixp5_ASAP7_75t_SL g282 ( .A1(n_262), .A2(n_228), .B(n_205), .C(n_222), .Y(n_282) );
AO221x2_ASAP7_75t_L g283 ( .A1(n_239), .A2(n_10), .B1(n_12), .B2(n_13), .C(n_15), .Y(n_283) );
A2O1A1Ixp33_ASAP7_75t_L g284 ( .A1(n_234), .A2(n_197), .B(n_196), .C(n_226), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_249), .A2(n_221), .B(n_222), .Y(n_285) );
OAI21xp5_ASAP7_75t_L g286 ( .A1(n_247), .A2(n_197), .B(n_208), .Y(n_286) );
OAI21xp5_ASAP7_75t_L g287 ( .A1(n_247), .A2(n_208), .B(n_192), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_274), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_235), .B(n_192), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_272), .A2(n_191), .B1(n_227), .B2(n_229), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_237), .B(n_10), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_261), .B(n_12), .Y(n_292) );
AOI22xp33_ASAP7_75t_SL g293 ( .A1(n_269), .A2(n_13), .B1(n_15), .B2(n_16), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_236), .B(n_16), .Y(n_294) );
AO32x2_ASAP7_75t_L g295 ( .A1(n_264), .A2(n_160), .A3(n_20), .B1(n_23), .B2(n_24), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_253), .B(n_18), .Y(n_296) );
NOR2xp33_ASAP7_75t_SL g297 ( .A(n_236), .B(n_238), .Y(n_297) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_242), .A2(n_25), .B(n_26), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_L g299 ( .A1(n_246), .A2(n_184), .B(n_29), .C(n_30), .Y(n_299) );
BUFx2_ASAP7_75t_L g300 ( .A(n_236), .Y(n_300) );
NOR2xp67_ASAP7_75t_SL g301 ( .A(n_238), .B(n_28), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_251), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_274), .Y(n_303) );
O2A1O1Ixp33_ASAP7_75t_SL g304 ( .A1(n_275), .A2(n_34), .B(n_35), .C(n_36), .Y(n_304) );
OAI21x1_ASAP7_75t_L g305 ( .A1(n_270), .A2(n_37), .B(n_39), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_272), .A2(n_160), .B1(n_42), .B2(n_43), .Y(n_306) );
OAI21xp5_ASAP7_75t_L g307 ( .A1(n_245), .A2(n_40), .B(n_44), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_255), .A2(n_160), .B(n_46), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_243), .B(n_45), .Y(n_309) );
AO32x2_ASAP7_75t_L g310 ( .A1(n_244), .A2(n_49), .A3(n_53), .B1(n_57), .B2(n_64), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_288), .Y(n_311) );
AOI221xp5_ASAP7_75t_L g312 ( .A1(n_281), .A2(n_257), .B1(n_273), .B2(n_256), .C(n_254), .Y(n_312) );
O2A1O1Ixp33_ASAP7_75t_L g313 ( .A1(n_281), .A2(n_254), .B(n_276), .C(n_260), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_280), .A2(n_258), .B(n_270), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_303), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_289), .B(n_276), .Y(n_316) );
OAI21x1_ASAP7_75t_L g317 ( .A1(n_308), .A2(n_233), .B(n_265), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_284), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_280), .A2(n_244), .B(n_265), .Y(n_319) );
OR2x6_ASAP7_75t_L g320 ( .A(n_294), .B(n_238), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_292), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_290), .A2(n_248), .B1(n_267), .B2(n_263), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_278), .Y(n_323) );
A2O1A1Ixp33_ASAP7_75t_L g324 ( .A1(n_299), .A2(n_260), .B(n_268), .C(n_259), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_278), .B(n_252), .Y(n_325) );
INVx2_ASAP7_75t_SL g326 ( .A(n_300), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_291), .B(n_252), .Y(n_327) );
BUFx2_ASAP7_75t_SL g328 ( .A(n_294), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_277), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_287), .Y(n_330) );
AO21x2_ASAP7_75t_L g331 ( .A1(n_279), .A2(n_240), .B(n_266), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_286), .B(n_252), .Y(n_332) );
AO21x2_ASAP7_75t_L g333 ( .A1(n_308), .A2(n_66), .B(n_67), .Y(n_333) );
OAI21x1_ASAP7_75t_L g334 ( .A1(n_298), .A2(n_68), .B(n_69), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_302), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_295), .Y(n_336) );
NAND2x1p5_ASAP7_75t_L g337 ( .A(n_301), .B(n_82), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_326), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_315), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_315), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_311), .B(n_283), .Y(n_341) );
BUFx5_ASAP7_75t_L g342 ( .A(n_332), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_312), .A2(n_283), .B1(n_316), .B2(n_321), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_311), .B(n_293), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_332), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_336), .Y(n_346) );
BUFx2_ASAP7_75t_L g347 ( .A(n_320), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_320), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_335), .B(n_293), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_326), .Y(n_350) );
OA21x2_ASAP7_75t_L g351 ( .A1(n_336), .A2(n_285), .B(n_307), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_318), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_318), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_325), .Y(n_354) );
AO21x2_ASAP7_75t_L g355 ( .A1(n_314), .A2(n_285), .B(n_304), .Y(n_355) );
AOI211xp5_ASAP7_75t_SL g356 ( .A1(n_322), .A2(n_297), .B(n_296), .C(n_309), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_328), .B(n_306), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_331), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_331), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_335), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_323), .B(n_328), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_330), .B(n_306), .Y(n_362) );
OA21x2_ASAP7_75t_L g363 ( .A1(n_319), .A2(n_305), .B(n_310), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_330), .B(n_282), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_346), .Y(n_365) );
INVxp67_ASAP7_75t_SL g366 ( .A(n_358), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_345), .B(n_340), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_345), .B(n_331), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_346), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_342), .B(n_310), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_346), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_342), .B(n_310), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_339), .Y(n_373) );
NOR2x1_ASAP7_75t_L g374 ( .A(n_347), .B(n_320), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_358), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_358), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_359), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_342), .B(n_310), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_347), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_342), .B(n_295), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_339), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_340), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_353), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_353), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_342), .B(n_323), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_350), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_342), .B(n_353), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_352), .B(n_313), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_352), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_348), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_343), .A2(n_327), .B1(n_320), .B2(n_329), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_360), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_359), .Y(n_393) );
AO21x2_ASAP7_75t_L g394 ( .A1(n_364), .A2(n_317), .B(n_333), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_341), .B(n_333), .Y(n_395) );
BUFx2_ASAP7_75t_L g396 ( .A(n_342), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_359), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_360), .Y(n_398) );
INVx5_ASAP7_75t_L g399 ( .A(n_348), .Y(n_399) );
INVxp67_ASAP7_75t_L g400 ( .A(n_341), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_387), .B(n_342), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_387), .B(n_342), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_373), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_387), .B(n_342), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_373), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_368), .B(n_344), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_375), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_368), .B(n_344), .Y(n_408) );
INVx1_ASAP7_75t_SL g409 ( .A(n_386), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_386), .Y(n_410) );
INVx3_ASAP7_75t_L g411 ( .A(n_368), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_381), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_368), .B(n_349), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_367), .B(n_349), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_400), .B(n_364), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_375), .Y(n_416) );
BUFx2_ASAP7_75t_L g417 ( .A(n_396), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_381), .Y(n_418) );
INVx1_ASAP7_75t_SL g419 ( .A(n_396), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_379), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_400), .B(n_338), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_367), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_382), .B(n_362), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_365), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_392), .B(n_354), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_382), .Y(n_426) );
INVx8_ASAP7_75t_L g427 ( .A(n_399), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_392), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_365), .Y(n_429) );
AND2x4_ASAP7_75t_SL g430 ( .A(n_385), .B(n_361), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_398), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_398), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_375), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_380), .B(n_362), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_380), .B(n_351), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_369), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_380), .B(n_351), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_369), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_370), .B(n_351), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_395), .B(n_357), .Y(n_440) );
AND2x4_ASAP7_75t_L g441 ( .A(n_371), .B(n_361), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_389), .B(n_357), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_371), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_395), .B(n_351), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_370), .B(n_363), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_370), .B(n_363), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_389), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_372), .B(n_363), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_385), .B(n_356), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_379), .Y(n_450) );
NOR2x1p5_ASAP7_75t_L g451 ( .A(n_379), .B(n_356), .Y(n_451) );
INVx2_ASAP7_75t_SL g452 ( .A(n_399), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_407), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_422), .B(n_388), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_410), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_403), .Y(n_456) );
INVxp67_ASAP7_75t_L g457 ( .A(n_417), .Y(n_457) );
AOI21xp33_ASAP7_75t_SL g458 ( .A1(n_427), .A2(n_391), .B(n_378), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_403), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_407), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_405), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_405), .Y(n_462) );
INVx2_ASAP7_75t_SL g463 ( .A(n_427), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_452), .B(n_399), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_452), .B(n_399), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_411), .B(n_390), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_412), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_407), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_409), .B(n_388), .Y(n_469) );
NOR2xp33_ASAP7_75t_SL g470 ( .A(n_427), .B(n_399), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_414), .B(n_390), .Y(n_471) );
NOR2xp67_ASAP7_75t_SL g472 ( .A(n_417), .B(n_399), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_440), .B(n_390), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_430), .B(n_399), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_430), .B(n_378), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_434), .B(n_383), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_430), .B(n_372), .Y(n_477) );
INVx1_ASAP7_75t_SL g478 ( .A(n_419), .Y(n_478) );
INVxp67_ASAP7_75t_L g479 ( .A(n_415), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_434), .B(n_383), .Y(n_480) );
INVx2_ASAP7_75t_SL g481 ( .A(n_427), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_412), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_425), .B(n_384), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_418), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_440), .B(n_384), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_406), .B(n_374), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_423), .B(n_397), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_418), .Y(n_488) );
INVxp33_ASAP7_75t_L g489 ( .A(n_451), .Y(n_489) );
NAND2xp33_ASAP7_75t_L g490 ( .A(n_427), .B(n_374), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_416), .Y(n_491) );
INVx1_ASAP7_75t_SL g492 ( .A(n_420), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_426), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_442), .B(n_397), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_406), .B(n_397), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_408), .B(n_376), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_426), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_423), .B(n_393), .Y(n_498) );
INVx2_ASAP7_75t_SL g499 ( .A(n_450), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_416), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_428), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_428), .Y(n_502) );
NOR3xp33_ASAP7_75t_L g503 ( .A(n_421), .B(n_299), .C(n_324), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_408), .B(n_413), .Y(n_504) );
AND2x4_ASAP7_75t_L g505 ( .A(n_411), .B(n_393), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_416), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_413), .B(n_393), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_431), .B(n_377), .Y(n_508) );
BUFx2_ASAP7_75t_L g509 ( .A(n_441), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_401), .B(n_402), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_451), .A2(n_333), .B1(n_394), .B2(n_376), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_479), .B(n_415), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_510), .B(n_445), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_479), .B(n_446), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_495), .B(n_445), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_469), .B(n_446), .Y(n_516) );
NAND4xp25_ASAP7_75t_L g517 ( .A(n_511), .B(n_449), .C(n_411), .D(n_444), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_455), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_496), .B(n_411), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_504), .B(n_435), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_453), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_507), .B(n_435), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_454), .B(n_448), .Y(n_523) );
NOR2x1_ASAP7_75t_L g524 ( .A(n_464), .B(n_436), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_509), .B(n_441), .Y(n_525) );
NAND3xp33_ASAP7_75t_L g526 ( .A(n_511), .B(n_447), .C(n_432), .Y(n_526) );
NAND3xp33_ASAP7_75t_L g527 ( .A(n_457), .B(n_447), .C(n_432), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_456), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_486), .B(n_437), .Y(n_529) );
INVx1_ASAP7_75t_SL g530 ( .A(n_478), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_459), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_461), .Y(n_532) );
NAND2x1_ASAP7_75t_L g533 ( .A(n_472), .B(n_429), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_505), .B(n_437), .Y(n_534) );
OAI21xp5_ASAP7_75t_L g535 ( .A1(n_489), .A2(n_441), .B(n_438), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_462), .Y(n_536) );
OAI322xp33_ASAP7_75t_SL g537 ( .A1(n_476), .A2(n_431), .A3(n_436), .B1(n_438), .B2(n_443), .C1(n_424), .C2(n_429), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_505), .B(n_439), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_505), .B(n_439), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_467), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_453), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_475), .B(n_448), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_492), .B(n_441), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_482), .Y(n_544) );
INVx2_ASAP7_75t_SL g545 ( .A(n_499), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_484), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_477), .B(n_404), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_489), .B(n_443), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_499), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_488), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_460), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_480), .B(n_404), .Y(n_552) );
A2O1A1Ixp33_ASAP7_75t_L g553 ( .A1(n_463), .A2(n_402), .B(n_401), .C(n_424), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_493), .Y(n_554) );
AOI32xp33_ASAP7_75t_L g555 ( .A1(n_490), .A2(n_444), .A3(n_433), .B1(n_334), .B2(n_366), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_497), .Y(n_556) );
INVxp67_ASAP7_75t_L g557 ( .A(n_473), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_500), .B(n_433), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_460), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_485), .B(n_487), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_501), .Y(n_561) );
NAND4xp25_ASAP7_75t_L g562 ( .A(n_517), .B(n_458), .C(n_503), .D(n_470), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_523), .B(n_457), .Y(n_563) );
OAI22xp33_ASAP7_75t_SL g564 ( .A1(n_533), .A2(n_465), .B1(n_464), .B2(n_463), .Y(n_564) );
INVxp33_ASAP7_75t_L g565 ( .A(n_549), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_530), .B(n_483), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_552), .B(n_512), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_548), .A2(n_490), .B1(n_471), .B2(n_503), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_518), .B(n_502), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_555), .B(n_481), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_512), .Y(n_571) );
AO21x1_ASAP7_75t_L g572 ( .A1(n_533), .A2(n_465), .B(n_474), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_560), .B(n_498), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_552), .B(n_494), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_560), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_553), .A2(n_543), .B1(n_525), .B2(n_557), .Y(n_576) );
INVxp33_ASAP7_75t_L g577 ( .A(n_524), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_528), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_520), .B(n_500), .Y(n_579) );
NAND2xp33_ASAP7_75t_L g580 ( .A(n_553), .B(n_466), .Y(n_580) );
AOI221xp5_ASAP7_75t_L g581 ( .A1(n_537), .A2(n_508), .B1(n_466), .B2(n_491), .C(n_468), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_520), .B(n_506), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_513), .B(n_506), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_531), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_532), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_536), .Y(n_586) );
NOR2xp33_ASAP7_75t_SL g587 ( .A(n_545), .B(n_466), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_540), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_525), .A2(n_491), .B1(n_468), .B2(n_433), .Y(n_589) );
OAI221xp5_ASAP7_75t_SL g590 ( .A1(n_526), .A2(n_366), .B1(n_377), .B2(n_376), .C(n_295), .Y(n_590) );
OAI32xp33_ASAP7_75t_L g591 ( .A1(n_545), .A2(n_337), .A3(n_377), .B1(n_295), .B2(n_394), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_558), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_514), .B(n_394), .Y(n_593) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_558), .Y(n_594) );
AOI321xp33_ASAP7_75t_L g595 ( .A1(n_570), .A2(n_525), .A3(n_516), .B1(n_534), .B2(n_539), .C(n_538), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_575), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_573), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_562), .A2(n_535), .B1(n_534), .B2(n_539), .Y(n_598) );
NOR2x1_ASAP7_75t_L g599 ( .A(n_580), .B(n_527), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_564), .A2(n_538), .B(n_519), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_576), .A2(n_519), .B1(n_529), .B2(n_547), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_594), .B(n_513), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_568), .A2(n_529), .B1(n_547), .B2(n_542), .Y(n_603) );
OAI211xp5_ASAP7_75t_L g604 ( .A1(n_581), .A2(n_566), .B(n_590), .C(n_591), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_571), .Y(n_605) );
XOR2xp5_ASAP7_75t_L g606 ( .A(n_565), .B(n_561), .Y(n_606) );
OAI21xp33_ASAP7_75t_SL g607 ( .A1(n_577), .A2(n_542), .B(n_515), .Y(n_607) );
OAI211xp5_ASAP7_75t_L g608 ( .A1(n_590), .A2(n_556), .B(n_554), .C(n_550), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_587), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_567), .B(n_515), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_569), .A2(n_546), .B1(n_544), .B2(n_522), .C(n_551), .Y(n_611) );
OAI21xp5_ASAP7_75t_L g612 ( .A1(n_594), .A2(n_522), .B(n_559), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_578), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_572), .B(n_559), .Y(n_614) );
AOI31xp33_ASAP7_75t_L g615 ( .A1(n_599), .A2(n_579), .A3(n_563), .B(n_593), .Y(n_615) );
NAND2xp33_ASAP7_75t_R g616 ( .A(n_600), .B(n_583), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_611), .B(n_569), .Y(n_617) );
NOR2xp33_ASAP7_75t_R g618 ( .A(n_609), .B(n_588), .Y(n_618) );
NOR2x1_ASAP7_75t_L g619 ( .A(n_614), .B(n_586), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_604), .A2(n_607), .B1(n_608), .B2(n_609), .C(n_596), .Y(n_620) );
AO221x1_ASAP7_75t_L g621 ( .A1(n_595), .A2(n_585), .B1(n_584), .B2(n_592), .C(n_589), .Y(n_621) );
OAI221xp5_ASAP7_75t_L g622 ( .A1(n_598), .A2(n_574), .B1(n_582), .B2(n_551), .C(n_541), .Y(n_622) );
NAND3xp33_ASAP7_75t_SL g623 ( .A(n_601), .B(n_337), .C(n_521), .Y(n_623) );
O2A1O1Ixp33_ASAP7_75t_L g624 ( .A1(n_612), .A2(n_541), .B(n_521), .C(n_337), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_606), .Y(n_625) );
NAND4xp75_ASAP7_75t_L g626 ( .A(n_620), .B(n_603), .C(n_605), .D(n_597), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_625), .B(n_613), .Y(n_627) );
OAI211xp5_ASAP7_75t_L g628 ( .A1(n_618), .A2(n_602), .B(n_610), .C(n_363), .Y(n_628) );
OAI211xp5_ASAP7_75t_L g629 ( .A1(n_619), .A2(n_334), .B(n_317), .C(n_394), .Y(n_629) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_617), .Y(n_630) );
AOI211xp5_ASAP7_75t_SL g631 ( .A1(n_615), .A2(n_355), .B(n_72), .C(n_73), .Y(n_631) );
BUFx2_ASAP7_75t_L g632 ( .A(n_627), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_630), .Y(n_633) );
NOR2xp67_ASAP7_75t_L g634 ( .A(n_628), .B(n_622), .Y(n_634) );
NOR5xp2_ASAP7_75t_L g635 ( .A(n_626), .B(n_621), .C(n_616), .D(n_624), .E(n_623), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_633), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_632), .B(n_629), .Y(n_637) );
BUFx2_ASAP7_75t_L g638 ( .A(n_636), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_637), .Y(n_639) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_639), .Y(n_640) );
OAI21xp5_ASAP7_75t_L g641 ( .A1(n_640), .A2(n_638), .B(n_632), .Y(n_641) );
OAI21xp5_ASAP7_75t_L g642 ( .A1(n_641), .A2(n_634), .B(n_635), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_642), .A2(n_631), .B(n_355), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_643), .A2(n_355), .B(n_642), .Y(n_644) );
endmodule