module fake_jpeg_20446_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_35),
.Y(n_42)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_15),
.B(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_14),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_41),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_30),
.B1(n_29),
.B2(n_15),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_44),
.B1(n_40),
.B2(n_18),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_30),
.B1(n_29),
.B2(n_21),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_52),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_22),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_22),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_58),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_30),
.B1(n_29),
.B2(n_34),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_52),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_70),
.B1(n_72),
.B2(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_71),
.Y(n_96)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_68),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_23),
.B1(n_27),
.B2(n_24),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_78),
.B1(n_47),
.B2(n_45),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_38),
.B1(n_32),
.B2(n_40),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_47),
.B1(n_51),
.B2(n_45),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_40),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_28),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_27),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_38),
.B1(n_32),
.B2(n_23),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_18),
.B1(n_24),
.B2(n_25),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_74),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_31),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_18),
.B1(n_25),
.B2(n_31),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_41),
.B1(n_36),
.B2(n_22),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_17),
.B1(n_19),
.B2(n_3),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_28),
.B1(n_26),
.B2(n_17),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_41),
.B(n_28),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_51),
.Y(n_80)
);

AO22x1_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_50),
.B1(n_26),
.B2(n_17),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_81),
.A2(n_83),
.B1(n_91),
.B2(n_97),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_73),
.A2(n_47),
.B1(n_51),
.B2(n_45),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_86),
.A2(n_61),
.B1(n_71),
.B2(n_62),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_67),
.C(n_79),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_57),
.A2(n_50),
.B1(n_41),
.B2(n_22),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_58),
.A2(n_50),
.B1(n_28),
.B2(n_19),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_66),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_57),
.A2(n_50),
.B1(n_19),
.B2(n_26),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_76),
.B1(n_72),
.B2(n_70),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_60),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_55),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_97),
.B1(n_87),
.B2(n_98),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_63),
.C(n_69),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_68),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_112),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_74),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_110),
.B(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

INVxp67_ASAP7_75t_SL g113 ( 
.A(n_84),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_124),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_64),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_6),
.B(n_7),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_88),
.B(n_99),
.Y(n_136)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_119),
.B(n_121),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_89),
.B(n_75),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_90),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_87),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_125),
.A2(n_84),
.B1(n_94),
.B2(n_102),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_133),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_118),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_93),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_115),
.A2(n_98),
.B1(n_95),
.B2(n_101),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_137),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_88),
.B1(n_86),
.B2(n_95),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_2),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_144),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_141),
.A2(n_119),
.B1(n_104),
.B2(n_116),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_7),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_7),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_148),
.Y(n_162)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_149),
.B(n_158),
.Y(n_167)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_L g171 ( 
.A1(n_153),
.A2(n_132),
.B1(n_128),
.B2(n_134),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_112),
.C(n_122),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_139),
.C(n_143),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_156),
.B(n_141),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_120),
.B(n_108),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_142),
.A2(n_120),
.B1(n_108),
.B2(n_123),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_159),
.A2(n_138),
.B1(n_123),
.B2(n_133),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_157),
.A2(n_136),
.B1(n_129),
.B2(n_138),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_163),
.B1(n_164),
.B2(n_171),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_157),
.A2(n_126),
.B1(n_137),
.B2(n_131),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_165),
.A2(n_153),
.B1(n_155),
.B2(n_150),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_159),
.C(n_152),
.Y(n_177)
);

AOI321xp33_ASAP7_75t_L g169 ( 
.A1(n_147),
.A2(n_143),
.A3(n_107),
.B1(n_144),
.B2(n_126),
.C(n_127),
.Y(n_169)
);

OAI322xp33_ASAP7_75t_L g180 ( 
.A1(n_169),
.A2(n_117),
.A3(n_118),
.B1(n_145),
.B2(n_150),
.C1(n_12),
.C2(n_8),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_154),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_172),
.B(n_177),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_167),
.B(n_152),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_174),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_147),
.C(n_151),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_175),
.A2(n_180),
.B(n_165),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_151),
.C(n_156),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_176),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_162),
.B(n_158),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_170),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_179),
.A2(n_168),
.B1(n_162),
.B2(n_170),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_184),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_187),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_168),
.B(n_169),
.Y(n_187)
);

NAND4xp25_ASAP7_75t_SL g188 ( 
.A(n_184),
.B(n_183),
.C(n_10),
.D(n_11),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_190),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_172),
.C(n_176),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_182),
.A2(n_117),
.B1(n_10),
.B2(n_11),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_191),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_117),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_195),
.C(n_196),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_192),
.B(n_188),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_194),
.A2(n_189),
.B(n_190),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_196),
.B(n_13),
.C(n_14),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_200),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_199),
.B1(n_9),
.B2(n_14),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_9),
.Y(n_203)
);


endmodule