module fake_jpeg_2921_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_0),
.B(n_2),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_19),
.Y(n_24)
);

INVx3_ASAP7_75t_SL g17 ( 
.A(n_7),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_17),
.B(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_9),
.B(n_6),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_22),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_10),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_3),
.C(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_1),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_16),
.A2(n_11),
.B1(n_7),
.B2(n_13),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_26),
.B(n_21),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_20),
.A2(n_12),
.B1(n_8),
.B2(n_7),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_23),
.C(n_22),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_36),
.B(n_38),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_39),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_24),
.C(n_27),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_43),
.C(n_15),
.Y(n_47)
);

AO22x1_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_17),
.B1(n_12),
.B2(n_8),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_44),
.B(n_41),
.C(n_17),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_35),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_34),
.B1(n_26),
.B2(n_8),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_47),
.B(n_40),
.Y(n_48)
);

OAI21x1_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_45),
.B(n_49),
.Y(n_50)
);

BUFx24_ASAP7_75t_SL g51 ( 
.A(n_50),
.Y(n_51)
);


endmodule