module fake_jpeg_26917_n_153 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_23),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_22),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_5),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_2),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_13),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_66),
.Y(n_82)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_0),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_69),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_76),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_60),
.B1(n_48),
.B2(n_47),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_85),
.B1(n_53),
.B2(n_2),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_47),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_71),
.A2(n_60),
.B1(n_55),
.B2(n_52),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_1),
.B(n_3),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_56),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_53),
.B1(n_61),
.B2(n_57),
.Y(n_85)
);

FAx1_ASAP7_75t_SL g88 ( 
.A(n_82),
.B(n_62),
.CI(n_54),
.CON(n_88),
.SN(n_88)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_90),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_59),
.B(n_58),
.C(n_45),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_43),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_46),
.B(n_50),
.C(n_51),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_96),
.B1(n_97),
.B2(n_99),
.Y(n_107)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_21),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_1),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_100),
.A2(n_101),
.B1(n_4),
.B2(n_5),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

AO22x1_ASAP7_75t_SL g102 ( 
.A1(n_93),
.A2(n_72),
.B1(n_77),
.B2(n_78),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_102),
.A2(n_87),
.B1(n_89),
.B2(n_92),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_98),
.A2(n_25),
.B1(n_42),
.B2(n_41),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_98),
.B1(n_86),
.B2(n_95),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_104),
.A2(n_103),
.B1(n_110),
.B2(n_106),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_119),
.B1(n_9),
.B2(n_10),
.Y(n_132)
);

NOR2x1_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_88),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_113),
.B1(n_7),
.B2(n_8),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_107),
.Y(n_114)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_110),
.A2(n_4),
.B(n_6),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_9),
.B(n_10),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_109),
.B(n_6),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_116),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_108),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_113),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_124),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_112),
.A2(n_104),
.B(n_105),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_123),
.B(n_130),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_129),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_31),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_27),
.Y(n_131)
);

AOI221xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.C(n_14),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_32),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_124),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_135),
.B(n_137),
.Y(n_144)
);

AOI322xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_37),
.A3(n_16),
.B1(n_18),
.B2(n_20),
.C1(n_24),
.C2(n_34),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_141),
.A2(n_142),
.B1(n_136),
.B2(n_128),
.Y(n_143)
);

OAI31xp33_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_15),
.A3(n_35),
.B(n_38),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

NOR2xp67_ASAP7_75t_SL g146 ( 
.A(n_145),
.B(n_144),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_146),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_143),
.C(n_138),
.Y(n_148)
);

AOI21x1_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_141),
.B(n_140),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_149),
.A2(n_120),
.B1(n_121),
.B2(n_139),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_126),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_140),
.C(n_39),
.Y(n_152)
);

BUFx24_ASAP7_75t_SL g153 ( 
.A(n_152),
.Y(n_153)
);


endmodule