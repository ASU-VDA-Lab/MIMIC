module fake_ibex_1488_n_1370 (n_151, n_147, n_85, n_167, n_128, n_208, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_61, n_201, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_215, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_213, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_214, n_79, n_81, n_35, n_159, n_202, n_158, n_211, n_218, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_184, n_31, n_56, n_23, n_146, n_91, n_207, n_54, n_19, n_1370);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_61;
input n_201;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_215;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_213;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_214;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_158;
input n_211;
input n_218;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_207;
input n_54;
input n_19;

output n_1370;

wire n_1084;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_280;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_242;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_235;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_230;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_793;
wire n_937;
wire n_234;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_573;
wire n_359;
wire n_433;
wire n_262;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_369;
wire n_1301;
wire n_257;
wire n_869;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_562;
wire n_564;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1108;
wire n_382;
wire n_1239;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_1281;
wire n_695;
wire n_639;
wire n_1332;
wire n_482;
wire n_282;
wire n_870;
wire n_1298;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_252;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_241;
wire n_231;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_256;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1015;
wire n_663;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_258;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1318;
wire n_421;
wire n_738;
wire n_1217;
wire n_236;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_840;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1364;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_267;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_413;
wire n_1069;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_998;
wire n_1115;
wire n_801;
wire n_1046;
wire n_882;
wire n_942;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_444;
wire n_986;
wire n_495;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_227;
wire n_1087;
wire n_757;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_318;
wire n_291;
wire n_268;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_997;
wire n_891;
wire n_303;
wire n_717;
wire n_1357;
wire n_668;
wire n_871;
wire n_266;
wire n_1339;
wire n_485;
wire n_1315;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_460;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1048;
wire n_774;
wire n_588;
wire n_1251;
wire n_1247;
wire n_528;
wire n_260;
wire n_836;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_920;
wire n_664;
wire n_1067;
wire n_255;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1331;
wire n_1223;
wire n_1349;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_226;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1367;
wire n_1291;
wire n_317;
wire n_326;
wire n_270;
wire n_1340;
wire n_259;
wire n_276;
wire n_339;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_251;
wire n_1112;
wire n_1267;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_224;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1188;
wire n_261;
wire n_742;
wire n_1191;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_269;
wire n_570;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_246;
wire n_922;
wire n_851;
wire n_993;
wire n_253;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_1169;
wire n_245;
wire n_571;
wire n_229;
wire n_648;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_804;
wire n_484;
wire n_480;
wire n_1057;
wire n_354;
wire n_516;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_248;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_277;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_247;
wire n_237;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1221;
wire n_284;
wire n_1047;
wire n_792;
wire n_1314;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_232;
wire n_1050;
wire n_599;
wire n_1060;
wire n_756;
wire n_1257;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1362;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_1330;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_249;
wire n_478;
wire n_239;
wire n_336;
wire n_861;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_828;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_698;
wire n_1061;
wire n_682;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_265;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_243;
wire n_228;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_244;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1074;
wire n_759;
wire n_953;
wire n_1180;
wire n_536;
wire n_1220;
wire n_467;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_263;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_735;
wire n_305;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1033;
wire n_627;
wire n_990;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_653;
wire n_1205;
wire n_238;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_225;
wire n_511;
wire n_381;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_233;
wire n_414;
wire n_378;
wire n_952;
wire n_264;
wire n_1145;
wire n_537;
wire n_1113;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_240;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_254;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_271;
wire n_984;
wire n_394;
wire n_364;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_90),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_17),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_10),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_184),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_97),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_10),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_147),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_76),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_86),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_208),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_174),
.Y(n_234)
);

BUFx2_ASAP7_75t_SL g235 ( 
.A(n_218),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_26),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_45),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_165),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_20),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_163),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_150),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_138),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_58),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_162),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_139),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_79),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_34),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_131),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_190),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_175),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_18),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_105),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_196),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_59),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_122),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_119),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_113),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_158),
.B(n_53),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_15),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_202),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_117),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_99),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_168),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_200),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_126),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_114),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_170),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_194),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_82),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_57),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_107),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_187),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_95),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_21),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_65),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_153),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_55),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_124),
.Y(n_279)
);

INVxp33_ASAP7_75t_SL g280 ( 
.A(n_60),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_48),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_179),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_188),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_71),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_152),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_210),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_171),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_211),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_92),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_157),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_75),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_32),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_21),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_195),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_32),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_161),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_120),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_178),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_77),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_106),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_146),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_183),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_35),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_136),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_7),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_30),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_207),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_5),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_15),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_217),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_1),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_38),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_111),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_155),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_156),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g316 ( 
.A(n_13),
.Y(n_316)
);

BUFx10_ASAP7_75t_L g317 ( 
.A(n_198),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_204),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_101),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_41),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_130),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_160),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_176),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_80),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_35),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_23),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_48),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_203),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_103),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_4),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_201),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_182),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_100),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_33),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_186),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_129),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_38),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_145),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_109),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_180),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_193),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_177),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_16),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_11),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_43),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_199),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_140),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_197),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_189),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_47),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_54),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_132),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_173),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_191),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_50),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_137),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_26),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_11),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_54),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_154),
.Y(n_360)
);

NOR2xp67_ASAP7_75t_L g361 ( 
.A(n_69),
.B(n_46),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_185),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_20),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_133),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_222),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_151),
.Y(n_366)
);

BUFx10_ASAP7_75t_L g367 ( 
.A(n_59),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_128),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_33),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_53),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_72),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_159),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_135),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_39),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_115),
.B(n_64),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_205),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_215),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_167),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_116),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_34),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_209),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_172),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_144),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_7),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_102),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_118),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_81),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_104),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_66),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_123),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_206),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_L g392 ( 
.A(n_83),
.B(n_70),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_84),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_143),
.Y(n_394)
);

BUFx8_ASAP7_75t_SL g395 ( 
.A(n_142),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_58),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_192),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_17),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_96),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_64),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_62),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_98),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_316),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_250),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_250),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_305),
.B(n_0),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_395),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_367),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_316),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_395),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_0),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_292),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_266),
.Y(n_413)
);

BUFx8_ASAP7_75t_L g414 ( 
.A(n_256),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_321),
.Y(n_415)
);

BUFx8_ASAP7_75t_L g416 ( 
.A(n_318),
.Y(n_416)
);

OAI22x1_ASAP7_75t_L g417 ( 
.A1(n_355),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_396),
.B(n_2),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g419 ( 
.A(n_367),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_316),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_250),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_344),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_250),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_245),
.Y(n_424)
);

OA21x2_ASAP7_75t_L g425 ( 
.A1(n_298),
.A2(n_74),
.B(n_73),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_260),
.B(n_3),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_253),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_316),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_391),
.B(n_5),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_253),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_253),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_367),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_267),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_433)
);

CKINVDCx11_ASAP7_75t_R g434 ( 
.A(n_303),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_401),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_260),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_253),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_245),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_293),
.Y(n_439)
);

OAI22x1_ASAP7_75t_SL g440 ( 
.A1(n_303),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_257),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_316),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_316),
.Y(n_443)
);

BUFx8_ASAP7_75t_L g444 ( 
.A(n_265),
.Y(n_444)
);

INVx5_ASAP7_75t_L g445 ( 
.A(n_317),
.Y(n_445)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_317),
.Y(n_446)
);

BUFx12f_ASAP7_75t_L g447 ( 
.A(n_317),
.Y(n_447)
);

INVx6_ASAP7_75t_L g448 ( 
.A(n_257),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_281),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_257),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_281),
.B(n_12),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_337),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_337),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_257),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_282),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_290),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_338),
.B(n_13),
.Y(n_457)
);

INVx5_ASAP7_75t_L g458 ( 
.A(n_282),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_226),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_309),
.B(n_14),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_225),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_282),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_236),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_315),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_324),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_282),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_273),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_229),
.B(n_16),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_353),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_243),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_353),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_353),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_335),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_384),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_353),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_251),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_371),
.Y(n_477)
);

OA21x2_ASAP7_75t_L g478 ( 
.A1(n_371),
.A2(n_85),
.B(n_78),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_271),
.B(n_18),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_329),
.B(n_19),
.Y(n_480)
);

BUFx8_ASAP7_75t_SL g481 ( 
.A(n_400),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g482 ( 
.A1(n_377),
.A2(n_149),
.B(n_220),
.Y(n_482)
);

INVx5_ASAP7_75t_L g483 ( 
.A(n_376),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_275),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_377),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_237),
.Y(n_486)
);

OA21x2_ASAP7_75t_L g487 ( 
.A1(n_390),
.A2(n_148),
.B(n_219),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_278),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_269),
.B(n_19),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_390),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_239),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_400),
.Y(n_492)
);

OAI21x1_ASAP7_75t_L g493 ( 
.A1(n_228),
.A2(n_141),
.B(n_216),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_232),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_233),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_376),
.Y(n_496)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_376),
.Y(n_497)
);

INVx5_ASAP7_75t_L g498 ( 
.A(n_237),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_234),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_240),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_308),
.B(n_22),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_300),
.B(n_23),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_312),
.B(n_24),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_340),
.B(n_25),
.Y(n_504)
);

CKINVDCx6p67_ASAP7_75t_R g505 ( 
.A(n_235),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_242),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_237),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_426),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_407),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_426),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_439),
.Y(n_511)
);

AND3x2_ASAP7_75t_L g512 ( 
.A(n_422),
.B(n_378),
.C(n_326),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_451),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_410),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_413),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_408),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_451),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_461),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_411),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_467),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_403),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_404),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_411),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_461),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_474),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_403),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_474),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_481),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_481),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_434),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_434),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_492),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_447),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_418),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_468),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_414),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_409),
.Y(n_537)
);

INVxp33_ASAP7_75t_L g538 ( 
.A(n_463),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_491),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_468),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_453),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_463),
.Y(n_542)
);

BUFx10_ASAP7_75t_L g543 ( 
.A(n_419),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_416),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_416),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_453),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_412),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_446),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_479),
.Y(n_549)
);

AO22x2_ASAP7_75t_L g550 ( 
.A1(n_460),
.A2(n_375),
.B1(n_330),
.B2(n_345),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_446),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_480),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_R g553 ( 
.A(n_432),
.B(n_322),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_505),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_444),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_444),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_R g557 ( 
.A(n_432),
.B(n_322),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_420),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_445),
.B(n_224),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_445),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_445),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_445),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_R g563 ( 
.A(n_415),
.B(n_373),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_440),
.Y(n_564)
);

NOR2xp67_ASAP7_75t_L g565 ( 
.A(n_459),
.B(n_244),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_456),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_456),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_433),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_435),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_473),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_429),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_499),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_485),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_490),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_490),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_424),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_438),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_406),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_438),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_457),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_470),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_404),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_476),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_484),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_442),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_R g586 ( 
.A(n_488),
.B(n_373),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_494),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_R g588 ( 
.A(n_436),
.B(n_381),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_495),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_R g590 ( 
.A(n_425),
.B(n_280),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_464),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_489),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_465),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_R g594 ( 
.A(n_449),
.B(n_381),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_500),
.B(n_254),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_506),
.B(n_252),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_SL g597 ( 
.A(n_502),
.B(n_288),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_R g598 ( 
.A(n_452),
.B(n_397),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_477),
.B(n_255),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_443),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_504),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_417),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_501),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_503),
.B(n_276),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_428),
.Y(n_605)
);

NOR2xp67_ASAP7_75t_L g606 ( 
.A(n_486),
.B(n_262),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_425),
.Y(n_607)
);

OAI21x1_ASAP7_75t_L g608 ( 
.A1(n_482),
.A2(n_270),
.B(n_264),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_448),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_498),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_448),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_498),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_498),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_493),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_425),
.B(n_398),
.Y(n_615)
);

AOI21x1_ASAP7_75t_L g616 ( 
.A1(n_478),
.A2(n_277),
.B(n_274),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_458),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_458),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_404),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_458),
.B(n_295),
.Y(n_620)
);

BUFx10_ASAP7_75t_L g621 ( 
.A(n_507),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_483),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_483),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_483),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_478),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_478),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_497),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_507),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_R g629 ( 
.A(n_507),
.B(n_306),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_497),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_R g631 ( 
.A(n_507),
.B(n_311),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_497),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_404),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_487),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_405),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_405),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_405),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_405),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_421),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_421),
.B(n_320),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_423),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_423),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_423),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_496),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_487),
.A2(n_325),
.B1(n_334),
.B2(n_327),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_487),
.Y(n_646)
);

XOR2xp5_ASAP7_75t_L g647 ( 
.A(n_427),
.B(n_343),
.Y(n_647)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_496),
.B(n_350),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_427),
.Y(n_649)
);

BUFx10_ASAP7_75t_L g650 ( 
.A(n_427),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_579),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_591),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_587),
.B(n_589),
.Y(n_653)
);

NOR3xp33_ASAP7_75t_L g654 ( 
.A(n_602),
.B(n_539),
.C(n_511),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_591),
.Y(n_655)
);

BUFx5_ASAP7_75t_L g656 ( 
.A(n_614),
.Y(n_656)
);

INVx8_ASAP7_75t_L g657 ( 
.A(n_555),
.Y(n_657)
);

AND2x2_ASAP7_75t_SL g658 ( 
.A(n_597),
.B(n_357),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_548),
.B(n_238),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_547),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_551),
.B(n_313),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_538),
.B(n_359),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_541),
.Y(n_663)
);

OAI221xp5_ASAP7_75t_L g664 ( 
.A1(n_569),
.A2(n_358),
.B1(n_370),
.B2(n_369),
.C(n_363),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_516),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_572),
.B(n_227),
.Y(n_666)
);

NOR2x1p5_ASAP7_75t_L g667 ( 
.A(n_536),
.B(n_374),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_L g668 ( 
.A(n_607),
.B(n_230),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_546),
.Y(n_669)
);

NOR3xp33_ASAP7_75t_L g670 ( 
.A(n_518),
.B(n_389),
.C(n_380),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_609),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_578),
.B(n_231),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_574),
.B(n_241),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_581),
.B(n_246),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_611),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_575),
.B(n_248),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_604),
.B(n_583),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_570),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_519),
.A2(n_351),
.B1(n_247),
.B2(n_283),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_524),
.B(n_361),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_573),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_556),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_584),
.B(n_249),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_535),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_540),
.Y(n_685)
);

NOR2xp67_ASAP7_75t_L g686 ( 
.A(n_533),
.B(n_25),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_586),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_523),
.B(n_258),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_593),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_542),
.B(n_532),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_534),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_508),
.Y(n_692)
);

INVx8_ASAP7_75t_L g693 ( 
.A(n_554),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_576),
.B(n_261),
.Y(n_694)
);

NAND3xp33_ASAP7_75t_L g695 ( 
.A(n_645),
.B(n_259),
.C(n_297),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_577),
.B(n_263),
.Y(n_696)
);

INVx8_ASAP7_75t_L g697 ( 
.A(n_566),
.Y(n_697)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_647),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_510),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_513),
.Y(n_700)
);

A2O1A1Ixp33_ASAP7_75t_L g701 ( 
.A1(n_596),
.A2(n_599),
.B(n_517),
.C(n_549),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_595),
.B(n_299),
.Y(n_702)
);

INVx5_ASAP7_75t_L g703 ( 
.A(n_650),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_596),
.B(n_319),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_640),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_580),
.B(n_268),
.Y(n_706)
);

NAND3xp33_ASAP7_75t_L g707 ( 
.A(n_590),
.B(n_331),
.C(n_323),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_567),
.B(n_543),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_565),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_563),
.B(n_247),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_521),
.B(n_333),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_588),
.B(n_272),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_526),
.B(n_341),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_526),
.B(n_342),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_550),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_550),
.Y(n_716)
);

AO221x1_ASAP7_75t_L g717 ( 
.A1(n_563),
.A2(n_247),
.B1(n_351),
.B2(n_349),
.C(n_346),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_550),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_606),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_537),
.B(n_360),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_592),
.B(n_279),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_588),
.B(n_284),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_560),
.B(n_285),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_561),
.B(n_286),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_562),
.B(n_287),
.Y(n_725)
);

NOR2xp67_ASAP7_75t_L g726 ( 
.A(n_544),
.B(n_27),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_620),
.B(n_289),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_559),
.B(n_291),
.Y(n_728)
);

AOI221xp5_ASAP7_75t_L g729 ( 
.A1(n_594),
.A2(n_247),
.B1(n_351),
.B2(n_362),
.C(n_366),
.Y(n_729)
);

INVxp67_ASAP7_75t_SL g730 ( 
.A(n_615),
.Y(n_730)
);

INVx8_ASAP7_75t_L g731 ( 
.A(n_509),
.Y(n_731)
);

INVxp33_ASAP7_75t_L g732 ( 
.A(n_598),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_601),
.B(n_294),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_558),
.B(n_296),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_585),
.B(n_301),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_603),
.B(n_302),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_605),
.Y(n_737)
);

AOI221xp5_ASAP7_75t_L g738 ( 
.A1(n_553),
.A2(n_557),
.B1(n_598),
.B2(n_552),
.C(n_568),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_605),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_557),
.B(n_304),
.Y(n_740)
);

NAND2xp33_ASAP7_75t_L g741 ( 
.A(n_634),
.B(n_307),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_571),
.B(n_310),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_512),
.B(n_314),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_600),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_608),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_621),
.Y(n_746)
);

NOR3xp33_ASAP7_75t_L g747 ( 
.A(n_564),
.B(n_387),
.C(n_385),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_625),
.B(n_328),
.Y(n_748)
);

INVx5_ASAP7_75t_L g749 ( 
.A(n_522),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_625),
.B(n_332),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_633),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_635),
.Y(n_752)
);

INVxp67_ASAP7_75t_L g753 ( 
.A(n_648),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_626),
.B(n_336),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_636),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_646),
.Y(n_756)
);

NOR3xp33_ASAP7_75t_L g757 ( 
.A(n_515),
.B(n_393),
.C(n_388),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_646),
.B(n_339),
.Y(n_758)
);

NOR3xp33_ASAP7_75t_L g759 ( 
.A(n_520),
.B(n_399),
.C(n_394),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_514),
.B(n_545),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_629),
.B(n_347),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_616),
.B(n_348),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_629),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_530),
.B(n_352),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_637),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_631),
.B(n_354),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_638),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_610),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_617),
.B(n_356),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_531),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_618),
.B(n_364),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_612),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_613),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_622),
.B(n_365),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_623),
.B(n_368),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_624),
.B(n_372),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_641),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_627),
.B(n_379),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_630),
.B(n_382),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_663),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_669),
.Y(n_781)
);

INVx4_ASAP7_75t_L g782 ( 
.A(n_703),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_684),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_715),
.A2(n_383),
.B1(n_386),
.B2(n_402),
.Y(n_784)
);

NOR3xp33_ASAP7_75t_SL g785 ( 
.A(n_664),
.B(n_529),
.C(n_528),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_660),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_665),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_756),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_690),
.B(n_525),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_685),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_697),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_692),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_653),
.Y(n_793)
);

NAND3xp33_ASAP7_75t_SL g794 ( 
.A(n_738),
.B(n_677),
.C(n_732),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_699),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_662),
.B(n_527),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_665),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_718),
.A2(n_392),
.B1(n_643),
.B2(n_642),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_653),
.B(n_632),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_687),
.Y(n_800)
);

INVx4_ASAP7_75t_L g801 ( 
.A(n_703),
.Y(n_801)
);

BUFx4f_ASAP7_75t_L g802 ( 
.A(n_657),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_L g803 ( 
.A1(n_701),
.A2(n_471),
.B1(n_431),
.B2(n_437),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_700),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_691),
.B(n_28),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_768),
.B(n_28),
.Y(n_806)
);

NOR2xp67_ASAP7_75t_L g807 ( 
.A(n_707),
.B(n_87),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_721),
.B(n_29),
.Y(n_808)
);

BUFx8_ASAP7_75t_L g809 ( 
.A(n_770),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_697),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_703),
.Y(n_811)
);

NOR2x1p5_ASAP7_75t_L g812 ( 
.A(n_682),
.B(n_29),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_733),
.B(n_30),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_697),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_746),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_707),
.A2(n_471),
.B1(n_431),
.B2(n_437),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_731),
.B(n_31),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_731),
.B(n_36),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_736),
.B(n_742),
.Y(n_819)
);

OR2x6_ASAP7_75t_L g820 ( 
.A(n_731),
.B(n_430),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_777),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_672),
.B(n_37),
.Y(n_822)
);

OR2x4_ASAP7_75t_L g823 ( 
.A(n_760),
.B(n_37),
.Y(n_823)
);

INVx5_ASAP7_75t_L g824 ( 
.A(n_777),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_SL g825 ( 
.A1(n_658),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_R g826 ( 
.A(n_693),
.B(n_40),
.Y(n_826)
);

NAND2x1p5_ASAP7_75t_L g827 ( 
.A(n_708),
.B(n_667),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_678),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_681),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_689),
.Y(n_830)
);

NOR2xp67_ASAP7_75t_L g831 ( 
.A(n_695),
.B(n_88),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_705),
.A2(n_628),
.B(n_430),
.C(n_469),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_657),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_657),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_693),
.Y(n_835)
);

NOR3xp33_ASAP7_75t_SL g836 ( 
.A(n_743),
.B(n_44),
.C(n_45),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_777),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_693),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_695),
.A2(n_471),
.B1(n_437),
.B2(n_441),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_702),
.B(n_49),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_772),
.B(n_773),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_651),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_668),
.A2(n_471),
.B1(n_437),
.B2(n_441),
.Y(n_843)
);

AND2x6_ASAP7_75t_SL g844 ( 
.A(n_764),
.B(n_51),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_671),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_698),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_674),
.B(n_683),
.Y(n_847)
);

BUFx12f_ASAP7_75t_L g848 ( 
.A(n_680),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_652),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_675),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_655),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_711),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_753),
.B(n_52),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_706),
.B(n_55),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_717),
.A2(n_472),
.B1(n_450),
.B2(n_454),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_710),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_704),
.B(n_56),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_709),
.B(n_56),
.Y(n_858)
);

AO22x1_ASAP7_75t_L g859 ( 
.A1(n_730),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_704),
.B(n_61),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_757),
.A2(n_472),
.B1(n_450),
.B2(n_454),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_759),
.A2(n_472),
.B1(n_450),
.B2(n_454),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_737),
.B(n_63),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_739),
.B(n_63),
.Y(n_864)
);

CKINVDCx11_ASAP7_75t_R g865 ( 
.A(n_763),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_711),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_713),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_670),
.A2(n_496),
.B1(n_455),
.B2(n_462),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_719),
.B(n_66),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_713),
.A2(n_496),
.B1(n_455),
.B2(n_462),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_726),
.B(n_67),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_745),
.A2(n_644),
.B(n_619),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_751),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_694),
.B(n_68),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_714),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_729),
.A2(n_469),
.B1(n_455),
.B2(n_462),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_744),
.B(n_714),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_720),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_659),
.B(n_661),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_750),
.A2(n_649),
.B(n_639),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_720),
.Y(n_881)
);

INVx4_ASAP7_75t_L g882 ( 
.A(n_749),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_654),
.B(n_466),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_712),
.B(n_89),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_696),
.B(n_91),
.Y(n_885)
);

NOR2x2_ASAP7_75t_L g886 ( 
.A(n_752),
.B(n_93),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_688),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_755),
.Y(n_888)
);

XOR2x2_ASAP7_75t_L g889 ( 
.A(n_747),
.B(n_94),
.Y(n_889)
);

O2A1O1Ixp5_ASAP7_75t_L g890 ( 
.A1(n_762),
.A2(n_639),
.B(n_582),
.C(n_522),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_740),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_765),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_741),
.A2(n_475),
.B1(n_639),
.B2(n_522),
.Y(n_893)
);

AND2x6_ASAP7_75t_L g894 ( 
.A(n_758),
.B(n_475),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_767),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_722),
.Y(n_896)
);

INVx5_ASAP7_75t_L g897 ( 
.A(n_749),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_686),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_769),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_673),
.B(n_522),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_793),
.B(n_666),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_852),
.A2(n_867),
.B1(n_875),
.B2(n_866),
.Y(n_902)
);

AOI22x1_ASAP7_75t_L g903 ( 
.A1(n_880),
.A2(n_582),
.B1(n_639),
.B2(n_656),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_809),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_878),
.B(n_676),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_877),
.A2(n_872),
.B(n_881),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_877),
.A2(n_748),
.B(n_754),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_780),
.B(n_771),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_781),
.B(n_771),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_822),
.A2(n_679),
.B(n_734),
.C(n_735),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_789),
.B(n_778),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_SL g912 ( 
.A(n_802),
.B(n_775),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_824),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_819),
.B(n_774),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_792),
.B(n_774),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_795),
.B(n_727),
.Y(n_916)
);

INVx4_ASAP7_75t_L g917 ( 
.A(n_802),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_782),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_794),
.B(n_779),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_857),
.A2(n_766),
.B1(n_761),
.B2(n_724),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_796),
.B(n_728),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_824),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_887),
.B(n_723),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_786),
.B(n_725),
.Y(n_924)
);

INVx4_ASAP7_75t_L g925 ( 
.A(n_782),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_821),
.B(n_776),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_804),
.B(n_749),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_801),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_828),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_788),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_860),
.A2(n_108),
.B(n_110),
.C(n_112),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_829),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_860),
.A2(n_121),
.B(n_125),
.C(n_127),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_830),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_SL g935 ( 
.A(n_835),
.B(n_134),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_833),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_834),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_840),
.A2(n_164),
.B(n_166),
.C(n_169),
.Y(n_938)
);

NOR2x1_ASAP7_75t_L g939 ( 
.A(n_838),
.B(n_181),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_809),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_817),
.Y(n_941)
);

BUFx2_ASAP7_75t_SL g942 ( 
.A(n_897),
.Y(n_942)
);

NOR3xp33_ASAP7_75t_SL g943 ( 
.A(n_891),
.B(n_899),
.C(n_854),
.Y(n_943)
);

BUFx4f_ASAP7_75t_L g944 ( 
.A(n_820),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_826),
.Y(n_945)
);

INVx5_ASAP7_75t_L g946 ( 
.A(n_820),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_801),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_847),
.B(n_892),
.Y(n_948)
);

CKINVDCx10_ASAP7_75t_R g949 ( 
.A(n_820),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_811),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_837),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_900),
.A2(n_212),
.B(n_213),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_846),
.B(n_810),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_841),
.B(n_214),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_805),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_806),
.A2(n_223),
.B1(n_808),
.B2(n_813),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_806),
.B(n_785),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_874),
.A2(n_858),
.B1(n_869),
.B2(n_853),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_791),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_841),
.B(n_814),
.Y(n_960)
);

OAI21x1_ASAP7_75t_L g961 ( 
.A1(n_893),
.A2(n_864),
.B(n_863),
.Y(n_961)
);

OAI21x1_ASAP7_75t_L g962 ( 
.A1(n_893),
.A2(n_864),
.B(n_863),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_799),
.B(n_874),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_783),
.B(n_790),
.Y(n_964)
);

AND2x6_ASAP7_75t_L g965 ( 
.A(n_858),
.B(n_885),
.Y(n_965)
);

AOI221xp5_ASAP7_75t_L g966 ( 
.A1(n_800),
.A2(n_869),
.B1(n_895),
.B2(n_873),
.C(n_859),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_897),
.Y(n_967)
);

INVx5_ASAP7_75t_L g968 ( 
.A(n_815),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_SL g969 ( 
.A1(n_855),
.A2(n_884),
.B(n_839),
.C(n_862),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_888),
.B(n_885),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_831),
.A2(n_807),
.B(n_868),
.C(n_856),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_807),
.A2(n_832),
.B(n_842),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_818),
.B(n_871),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_812),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_845),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_850),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_883),
.B(n_882),
.Y(n_977)
);

BUFx8_ASAP7_75t_L g978 ( 
.A(n_848),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_896),
.B(n_827),
.Y(n_979)
);

BUFx8_ASAP7_75t_L g980 ( 
.A(n_871),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_849),
.Y(n_981)
);

NOR2xp67_ASAP7_75t_L g982 ( 
.A(n_898),
.B(n_798),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_851),
.Y(n_983)
);

AOI22xp33_ASAP7_75t_L g984 ( 
.A1(n_865),
.A2(n_825),
.B1(n_787),
.B2(n_797),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_797),
.A2(n_889),
.B1(n_784),
.B2(n_798),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_823),
.B(n_844),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_816),
.A2(n_861),
.B(n_870),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_894),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_870),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_836),
.B(n_868),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_894),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_894),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_894),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_844),
.B(n_843),
.Y(n_994)
);

AOI22xp33_ASAP7_75t_L g995 ( 
.A1(n_876),
.A2(n_715),
.B1(n_718),
.B2(n_716),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_886),
.B(n_660),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_793),
.B(n_715),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_793),
.B(n_586),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_793),
.B(n_586),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_793),
.B(n_715),
.Y(n_1000)
);

NAND2x1p5_ASAP7_75t_L g1001 ( 
.A(n_802),
.B(n_833),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_824),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_821),
.Y(n_1003)
);

AO32x1_ASAP7_75t_L g1004 ( 
.A1(n_803),
.A2(n_615),
.A3(n_856),
.B1(n_883),
.B2(n_745),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_880),
.A2(n_877),
.B(n_756),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_872),
.A2(n_890),
.B(n_745),
.Y(n_1006)
);

INVxp67_ASAP7_75t_L g1007 ( 
.A(n_809),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_802),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_793),
.B(n_586),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_809),
.Y(n_1010)
);

BUFx4f_ASAP7_75t_L g1011 ( 
.A(n_820),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_780),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_809),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_794),
.A2(n_664),
.B(n_701),
.C(n_677),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_793),
.B(n_715),
.Y(n_1015)
);

BUFx4f_ASAP7_75t_L g1016 ( 
.A(n_820),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_793),
.B(n_660),
.Y(n_1017)
);

AOI21xp33_ASAP7_75t_L g1018 ( 
.A1(n_879),
.A2(n_733),
.B(n_721),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_793),
.B(n_578),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_880),
.A2(n_877),
.B(n_756),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_793),
.B(n_715),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_852),
.A2(n_866),
.B1(n_875),
.B2(n_867),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_793),
.A2(n_603),
.B1(n_571),
.B2(n_547),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_780),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_1006),
.A2(n_903),
.B(n_1005),
.Y(n_1025)
);

CKINVDCx16_ASAP7_75t_R g1026 ( 
.A(n_945),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_978),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_1020),
.A2(n_962),
.B(n_961),
.Y(n_1028)
);

BUFx2_ASAP7_75t_SL g1029 ( 
.A(n_917),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_978),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_904),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_1010),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_906),
.A2(n_907),
.B(n_902),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_1013),
.Y(n_1034)
);

BUFx12f_ASAP7_75t_L g1035 ( 
.A(n_917),
.Y(n_1035)
);

INVx5_ASAP7_75t_L g1036 ( 
.A(n_967),
.Y(n_1036)
);

INVx1_ASAP7_75t_SL g1037 ( 
.A(n_942),
.Y(n_1037)
);

BUFx2_ASAP7_75t_SL g1038 ( 
.A(n_1008),
.Y(n_1038)
);

INVx3_ASAP7_75t_SL g1039 ( 
.A(n_1008),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1012),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_949),
.Y(n_1041)
);

NAND2x1p5_ASAP7_75t_L g1042 ( 
.A(n_944),
.B(n_1011),
.Y(n_1042)
);

INVxp67_ASAP7_75t_SL g1043 ( 
.A(n_1022),
.Y(n_1043)
);

CKINVDCx20_ASAP7_75t_R g1044 ( 
.A(n_980),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_1014),
.A2(n_916),
.B(n_910),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_SL g1046 ( 
.A1(n_965),
.A2(n_980),
.B1(n_954),
.B2(n_986),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_937),
.Y(n_1047)
);

AO21x2_ASAP7_75t_L g1048 ( 
.A1(n_987),
.A2(n_969),
.B(n_989),
.Y(n_1048)
);

OAI22xp33_ASAP7_75t_SL g1049 ( 
.A1(n_996),
.A2(n_963),
.B1(n_935),
.B2(n_944),
.Y(n_1049)
);

CKINVDCx11_ASAP7_75t_R g1050 ( 
.A(n_1002),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_SL g1051 ( 
.A1(n_970),
.A2(n_966),
.B(n_991),
.Y(n_1051)
);

NAND2x1p5_ASAP7_75t_L g1052 ( 
.A(n_1011),
.B(n_1016),
.Y(n_1052)
);

BUFx12f_ASAP7_75t_L g1053 ( 
.A(n_1001),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_929),
.B(n_932),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_SL g1055 ( 
.A(n_1016),
.B(n_965),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_954),
.B(n_923),
.Y(n_1056)
);

INVx6_ASAP7_75t_L g1057 ( 
.A(n_922),
.Y(n_1057)
);

AOI22x1_ASAP7_75t_L g1058 ( 
.A1(n_990),
.A2(n_952),
.B1(n_928),
.B2(n_925),
.Y(n_1058)
);

AOI22x1_ASAP7_75t_L g1059 ( 
.A1(n_925),
.A2(n_928),
.B1(n_993),
.B2(n_955),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_934),
.Y(n_1060)
);

INVx6_ASAP7_75t_L g1061 ( 
.A(n_922),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1019),
.B(n_914),
.Y(n_1062)
);

BUFx2_ASAP7_75t_R g1063 ( 
.A(n_901),
.Y(n_1063)
);

INVx1_ASAP7_75t_SL g1064 ( 
.A(n_953),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_946),
.Y(n_1065)
);

BUFx8_ASAP7_75t_L g1066 ( 
.A(n_957),
.Y(n_1066)
);

INVx4_ASAP7_75t_L g1067 ( 
.A(n_946),
.Y(n_1067)
);

OR2x2_ASAP7_75t_L g1068 ( 
.A(n_1023),
.B(n_1017),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_946),
.Y(n_1069)
);

BUFx12f_ASAP7_75t_L g1070 ( 
.A(n_960),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_968),
.Y(n_1071)
);

INVx6_ASAP7_75t_L g1072 ( 
.A(n_968),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_968),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1024),
.B(n_905),
.Y(n_1074)
);

INVx4_ASAP7_75t_L g1075 ( 
.A(n_940),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_SL g1076 ( 
.A1(n_939),
.A2(n_956),
.B(n_909),
.Y(n_1076)
);

AO21x2_ASAP7_75t_L g1077 ( 
.A1(n_931),
.A2(n_933),
.B(n_920),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_926),
.A2(n_938),
.B(n_950),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_921),
.B(n_1018),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_960),
.B(n_958),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_941),
.B(n_948),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_964),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_1003),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_1003),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_918),
.Y(n_1085)
);

BUFx12f_ASAP7_75t_L g1086 ( 
.A(n_959),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_SL g1087 ( 
.A(n_965),
.B(n_988),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_913),
.Y(n_1088)
);

NOR2x1_ASAP7_75t_L g1089 ( 
.A(n_918),
.B(n_947),
.Y(n_1089)
);

INVxp67_ASAP7_75t_SL g1090 ( 
.A(n_988),
.Y(n_1090)
);

AO21x2_ASAP7_75t_L g1091 ( 
.A1(n_982),
.A2(n_983),
.B(n_927),
.Y(n_1091)
);

OR2x6_ASAP7_75t_L g1092 ( 
.A(n_1007),
.B(n_974),
.Y(n_1092)
);

INVx6_ASAP7_75t_L g1093 ( 
.A(n_977),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_923),
.B(n_965),
.Y(n_1094)
);

INVx4_ASAP7_75t_L g1095 ( 
.A(n_951),
.Y(n_1095)
);

CKINVDCx11_ASAP7_75t_R g1096 ( 
.A(n_992),
.Y(n_1096)
);

NAND2x1p5_ASAP7_75t_L g1097 ( 
.A(n_992),
.B(n_977),
.Y(n_1097)
);

BUFx2_ASAP7_75t_R g1098 ( 
.A(n_973),
.Y(n_1098)
);

BUFx4_ASAP7_75t_SL g1099 ( 
.A(n_975),
.Y(n_1099)
);

AO21x2_ASAP7_75t_L g1100 ( 
.A1(n_908),
.A2(n_915),
.B(n_919),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_936),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_930),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_976),
.Y(n_1103)
);

BUFx2_ASAP7_75t_R g1104 ( 
.A(n_998),
.Y(n_1104)
);

CKINVDCx6p67_ASAP7_75t_R g1105 ( 
.A(n_999),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_995),
.A2(n_997),
.B(n_1015),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_981),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_979),
.Y(n_1108)
);

INVx1_ASAP7_75t_SL g1109 ( 
.A(n_1000),
.Y(n_1109)
);

BUFx2_ASAP7_75t_SL g1110 ( 
.A(n_1009),
.Y(n_1110)
);

INVx6_ASAP7_75t_L g1111 ( 
.A(n_912),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_1021),
.Y(n_1112)
);

AO21x2_ASAP7_75t_L g1113 ( 
.A1(n_1004),
.A2(n_994),
.B(n_924),
.Y(n_1113)
);

INVx6_ASAP7_75t_L g1114 ( 
.A(n_943),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_984),
.B(n_985),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_1004),
.Y(n_1116)
);

BUFx12f_ASAP7_75t_L g1117 ( 
.A(n_911),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1019),
.B(n_793),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_963),
.B(n_793),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1019),
.B(n_793),
.Y(n_1120)
);

OR2x6_ASAP7_75t_L g1121 ( 
.A(n_942),
.B(n_917),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_949),
.Y(n_1122)
);

BUFx12f_ASAP7_75t_L g1123 ( 
.A(n_904),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_967),
.Y(n_1124)
);

NAND2x1p5_ASAP7_75t_L g1125 ( 
.A(n_944),
.B(n_1011),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_902),
.B(n_852),
.Y(n_1126)
);

INVx1_ASAP7_75t_SL g1127 ( 
.A(n_942),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_978),
.Y(n_1128)
);

AO21x2_ASAP7_75t_L g1129 ( 
.A1(n_971),
.A2(n_972),
.B(n_962),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1062),
.B(n_1118),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_SL g1131 ( 
.A1(n_1115),
.A2(n_1056),
.B1(n_1055),
.B2(n_1043),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1036),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_1036),
.Y(n_1133)
);

CKINVDCx11_ASAP7_75t_R g1134 ( 
.A(n_1123),
.Y(n_1134)
);

CKINVDCx8_ASAP7_75t_R g1135 ( 
.A(n_1029),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1115),
.A2(n_1079),
.B1(n_1117),
.B2(n_1046),
.Y(n_1136)
);

NAND2x1p5_ASAP7_75t_L g1137 ( 
.A(n_1036),
.B(n_1037),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_1053),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1054),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1054),
.Y(n_1140)
);

OR2x2_ASAP7_75t_L g1141 ( 
.A(n_1064),
.B(n_1074),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_1036),
.Y(n_1142)
);

AO21x2_ASAP7_75t_L g1143 ( 
.A1(n_1033),
.A2(n_1028),
.B(n_1025),
.Y(n_1143)
);

INVxp33_ASAP7_75t_L g1144 ( 
.A(n_1050),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1068),
.B(n_1079),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1060),
.Y(n_1146)
);

BUFx2_ASAP7_75t_R g1147 ( 
.A(n_1027),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_SL g1148 ( 
.A1(n_1056),
.A2(n_1126),
.B(n_1049),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_1121),
.Y(n_1149)
);

INVx2_ASAP7_75t_SL g1150 ( 
.A(n_1099),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1046),
.A2(n_1100),
.B1(n_1080),
.B2(n_1043),
.Y(n_1151)
);

OAI22xp33_ASAP7_75t_SL g1152 ( 
.A1(n_1055),
.A2(n_1111),
.B1(n_1037),
.B2(n_1127),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_1094),
.B(n_1073),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_1044),
.Y(n_1154)
);

INVxp67_ASAP7_75t_SL g1155 ( 
.A(n_1102),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_1044),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1082),
.A2(n_1109),
.B1(n_1074),
.B2(n_1063),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1119),
.A2(n_1114),
.B1(n_1100),
.B2(n_1094),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1045),
.B(n_1106),
.Y(n_1159)
);

NAND2x1p5_ASAP7_75t_L g1160 ( 
.A(n_1127),
.B(n_1071),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1030),
.Y(n_1161)
);

OAI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1109),
.A2(n_1063),
.B1(n_1102),
.B2(n_1045),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1040),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_1099),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_1096),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1107),
.Y(n_1166)
);

NAND2xp33_ASAP7_75t_L g1167 ( 
.A(n_1042),
.B(n_1052),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_SL g1168 ( 
.A1(n_1051),
.A2(n_1076),
.B(n_1059),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_1128),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1120),
.B(n_1119),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_SL g1171 ( 
.A1(n_1049),
.A2(n_1087),
.B1(n_1125),
.B2(n_1052),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1103),
.Y(n_1172)
);

NAND2x1p5_ASAP7_75t_L g1173 ( 
.A(n_1071),
.B(n_1067),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1064),
.B(n_1101),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1106),
.B(n_1112),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_1121),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_1112),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1081),
.Y(n_1178)
);

OAI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1087),
.A2(n_1042),
.B1(n_1125),
.B2(n_1111),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_1035),
.Y(n_1180)
);

OAI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1111),
.A2(n_1041),
.B1(n_1105),
.B2(n_1112),
.Y(n_1181)
);

NAND2x1p5_ASAP7_75t_L g1182 ( 
.A(n_1067),
.B(n_1065),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1041),
.Y(n_1183)
);

NAND2x1p5_ASAP7_75t_L g1184 ( 
.A(n_1065),
.B(n_1047),
.Y(n_1184)
);

INVx5_ASAP7_75t_L g1185 ( 
.A(n_1072),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1114),
.Y(n_1186)
);

INVx4_ASAP7_75t_L g1187 ( 
.A(n_1039),
.Y(n_1187)
);

OAI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1088),
.A2(n_1122),
.B1(n_1075),
.B2(n_1069),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1114),
.Y(n_1189)
);

NAND2x1p5_ASAP7_75t_L g1190 ( 
.A(n_1073),
.B(n_1075),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1078),
.A2(n_1116),
.B(n_1058),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1101),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_SL g1193 ( 
.A1(n_1110),
.A2(n_1113),
.B1(n_1038),
.B2(n_1066),
.Y(n_1193)
);

NAND2xp33_ASAP7_75t_R g1194 ( 
.A(n_1031),
.B(n_1032),
.Y(n_1194)
);

BUFx4f_ASAP7_75t_L g1195 ( 
.A(n_1039),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1070),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_SL g1197 ( 
.A1(n_1113),
.A2(n_1066),
.B1(n_1093),
.B2(n_1116),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_1096),
.Y(n_1198)
);

OR2x6_ASAP7_75t_L g1199 ( 
.A(n_1148),
.B(n_1097),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1170),
.B(n_1108),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1159),
.B(n_1091),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1145),
.A2(n_1091),
.B1(n_1093),
.B2(n_1050),
.Y(n_1202)
);

CKINVDCx16_ASAP7_75t_R g1203 ( 
.A(n_1138),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_1177),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1159),
.B(n_1048),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_1195),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_1134),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_SL g1208 ( 
.A1(n_1157),
.A2(n_1097),
.B(n_1098),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1155),
.B(n_1124),
.Y(n_1209)
);

BUFx10_ASAP7_75t_L g1210 ( 
.A(n_1150),
.Y(n_1210)
);

NAND2xp33_ASAP7_75t_R g1211 ( 
.A(n_1149),
.B(n_1034),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_R g1212 ( 
.A(n_1135),
.B(n_1026),
.Y(n_1212)
);

OR2x6_ASAP7_75t_L g1213 ( 
.A(n_1162),
.B(n_1164),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1156),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1139),
.B(n_1048),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_1174),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_1195),
.Y(n_1217)
);

HB1xp67_ASAP7_75t_L g1218 ( 
.A(n_1155),
.Y(n_1218)
);

NAND2xp33_ASAP7_75t_R g1219 ( 
.A(n_1176),
.B(n_1092),
.Y(n_1219)
);

OAI222xp33_ASAP7_75t_L g1220 ( 
.A1(n_1157),
.A2(n_1089),
.B1(n_1085),
.B2(n_1092),
.C1(n_1095),
.C2(n_1098),
.Y(n_1220)
);

NOR2x1_ASAP7_75t_L g1221 ( 
.A(n_1187),
.B(n_1095),
.Y(n_1221)
);

OR2x6_ASAP7_75t_L g1222 ( 
.A(n_1162),
.B(n_1061),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1186),
.B(n_1086),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1130),
.B(n_1093),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1178),
.B(n_1057),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1146),
.Y(n_1226)
);

NOR3xp33_ASAP7_75t_SL g1227 ( 
.A(n_1194),
.B(n_1104),
.C(n_1090),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1141),
.Y(n_1228)
);

CKINVDCx11_ASAP7_75t_R g1229 ( 
.A(n_1154),
.Y(n_1229)
);

NAND3xp33_ASAP7_75t_SL g1230 ( 
.A(n_1171),
.B(n_1190),
.C(n_1136),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1161),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1187),
.Y(n_1232)
);

OR2x4_ASAP7_75t_L g1233 ( 
.A(n_1165),
.B(n_1124),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1131),
.A2(n_1057),
.B1(n_1061),
.B2(n_1077),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1171),
.A2(n_1167),
.B(n_1131),
.C(n_1151),
.Y(n_1235)
);

NAND3xp33_ASAP7_75t_SL g1236 ( 
.A(n_1190),
.B(n_1104),
.C(n_1084),
.Y(n_1236)
);

OR2x6_ASAP7_75t_L g1237 ( 
.A(n_1168),
.B(n_1072),
.Y(n_1237)
);

NAND2xp33_ASAP7_75t_R g1238 ( 
.A(n_1169),
.B(n_1092),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1175),
.A2(n_1084),
.B(n_1083),
.Y(n_1239)
);

BUFx10_ASAP7_75t_L g1240 ( 
.A(n_1180),
.Y(n_1240)
);

CKINVDCx16_ASAP7_75t_R g1241 ( 
.A(n_1165),
.Y(n_1241)
);

OR2x6_ASAP7_75t_L g1242 ( 
.A(n_1137),
.B(n_1072),
.Y(n_1242)
);

INVx4_ASAP7_75t_L g1243 ( 
.A(n_1237),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1205),
.B(n_1143),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1205),
.B(n_1143),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1215),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_SL g1247 ( 
.A(n_1232),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1233),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1218),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1230),
.A2(n_1189),
.B1(n_1158),
.B2(n_1140),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1201),
.Y(n_1251)
);

INVx2_ASAP7_75t_SL g1252 ( 
.A(n_1233),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1201),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1230),
.A2(n_1213),
.B1(n_1200),
.B2(n_1224),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_1222),
.B(n_1191),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1216),
.B(n_1129),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1213),
.A2(n_1228),
.B1(n_1222),
.B2(n_1225),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1204),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1226),
.B(n_1197),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1237),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1253),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1256),
.B(n_1197),
.Y(n_1262)
);

NOR2x1_ASAP7_75t_L g1263 ( 
.A(n_1248),
.B(n_1236),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1249),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1255),
.B(n_1199),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_1249),
.B(n_1251),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_1249),
.B(n_1251),
.Y(n_1267)
);

BUFx2_ASAP7_75t_SL g1268 ( 
.A(n_1247),
.Y(n_1268)
);

NOR2xp67_ASAP7_75t_L g1269 ( 
.A(n_1243),
.B(n_1208),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1255),
.B(n_1199),
.Y(n_1270)
);

AND2x2_ASAP7_75t_SL g1271 ( 
.A(n_1243),
.B(n_1209),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1248),
.B(n_1188),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1258),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1256),
.B(n_1239),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1256),
.B(n_1239),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1246),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1262),
.B(n_1244),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1273),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1266),
.Y(n_1279)
);

OR2x2_ASAP7_75t_L g1280 ( 
.A(n_1266),
.B(n_1253),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1267),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1261),
.B(n_1246),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1264),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1261),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1262),
.B(n_1244),
.Y(n_1285)
);

AND3x1_ASAP7_75t_L g1286 ( 
.A(n_1263),
.B(n_1208),
.C(n_1254),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1274),
.B(n_1244),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1274),
.B(n_1245),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_1268),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1275),
.B(n_1245),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1282),
.Y(n_1291)
);

INVx1_ASAP7_75t_SL g1292 ( 
.A(n_1289),
.Y(n_1292)
);

INVx1_ASAP7_75t_SL g1293 ( 
.A(n_1283),
.Y(n_1293)
);

OA222x2_ASAP7_75t_L g1294 ( 
.A1(n_1283),
.A2(n_1213),
.B1(n_1248),
.B2(n_1260),
.C1(n_1264),
.C2(n_1269),
.Y(n_1294)
);

NOR2xp67_ASAP7_75t_L g1295 ( 
.A(n_1278),
.B(n_1243),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1284),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1277),
.B(n_1275),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1279),
.B(n_1276),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1287),
.B(n_1245),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1287),
.B(n_1265),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1284),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1279),
.B(n_1144),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1288),
.B(n_1265),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1281),
.B(n_1265),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1277),
.B(n_1276),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1282),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1281),
.B(n_1265),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_1286),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1308),
.A2(n_1286),
.B(n_1272),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1300),
.B(n_1288),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1304),
.A2(n_1254),
.B1(n_1270),
.B2(n_1257),
.Y(n_1311)
);

OR2x6_ASAP7_75t_L g1312 ( 
.A(n_1295),
.B(n_1268),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1296),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_1302),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1299),
.B(n_1285),
.Y(n_1315)
);

NOR3xp33_ASAP7_75t_L g1316 ( 
.A(n_1292),
.B(n_1188),
.C(n_1220),
.Y(n_1316)
);

OAI21xp33_ASAP7_75t_L g1317 ( 
.A1(n_1293),
.A2(n_1285),
.B(n_1290),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1309),
.B(n_1299),
.Y(n_1318)
);

AOI21xp33_ASAP7_75t_L g1319 ( 
.A1(n_1314),
.A2(n_1211),
.B(n_1219),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1315),
.B(n_1305),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1311),
.A2(n_1295),
.B1(n_1304),
.B2(n_1307),
.Y(n_1321)
);

OAI221xp5_ASAP7_75t_L g1322 ( 
.A1(n_1316),
.A2(n_1250),
.B1(n_1257),
.B2(n_1235),
.C(n_1306),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1313),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1317),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1310),
.B(n_1291),
.Y(n_1325)
);

OAI221xp5_ASAP7_75t_L g1326 ( 
.A1(n_1312),
.A2(n_1250),
.B1(n_1306),
.B2(n_1291),
.C(n_1298),
.Y(n_1326)
);

OAI221xp5_ASAP7_75t_SL g1327 ( 
.A1(n_1312),
.A2(n_1202),
.B1(n_1294),
.B2(n_1181),
.C(n_1300),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_SL g1328 ( 
.A1(n_1319),
.A2(n_1217),
.B(n_1206),
.Y(n_1328)
);

XNOR2x2_ASAP7_75t_SL g1329 ( 
.A(n_1324),
.B(n_1147),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1318),
.B(n_1290),
.Y(n_1330)
);

O2A1O1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1327),
.A2(n_1231),
.B(n_1207),
.C(n_1196),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1326),
.B(n_1321),
.Y(n_1332)
);

AOI221xp5_ASAP7_75t_L g1333 ( 
.A1(n_1322),
.A2(n_1304),
.B1(n_1307),
.B2(n_1297),
.C(n_1212),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1320),
.B(n_1203),
.Y(n_1334)
);

NOR2x1_ASAP7_75t_L g1335 ( 
.A(n_1323),
.B(n_1221),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_SL g1336 ( 
.A1(n_1331),
.A2(n_1333),
.B(n_1329),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1330),
.B(n_1325),
.Y(n_1337)
);

NAND2x1_ASAP7_75t_L g1338 ( 
.A(n_1335),
.B(n_1243),
.Y(n_1338)
);

AOI211x1_ASAP7_75t_L g1339 ( 
.A1(n_1332),
.A2(n_1303),
.B(n_1181),
.C(n_1236),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1334),
.B(n_1307),
.Y(n_1340)
);

NOR3x1_ASAP7_75t_L g1341 ( 
.A(n_1328),
.B(n_1147),
.C(n_1229),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1334),
.Y(n_1342)
);

O2A1O1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1336),
.A2(n_1223),
.B(n_1184),
.C(n_1183),
.Y(n_1343)
);

NAND3xp33_ASAP7_75t_SL g1344 ( 
.A(n_1338),
.B(n_1214),
.C(n_1227),
.Y(n_1344)
);

OAI211xp5_ASAP7_75t_L g1345 ( 
.A1(n_1339),
.A2(n_1217),
.B(n_1165),
.C(n_1198),
.Y(n_1345)
);

O2A1O1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1342),
.A2(n_1184),
.B(n_1152),
.C(n_1160),
.Y(n_1346)
);

O2A1O1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1340),
.A2(n_1160),
.B(n_1179),
.C(n_1137),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1337),
.A2(n_1241),
.B(n_1217),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1341),
.A2(n_1298),
.B1(n_1303),
.B2(n_1271),
.Y(n_1349)
);

AOI221xp5_ASAP7_75t_L g1350 ( 
.A1(n_1339),
.A2(n_1192),
.B1(n_1296),
.B2(n_1301),
.C(n_1234),
.Y(n_1350)
);

AO22x2_ASAP7_75t_L g1351 ( 
.A1(n_1345),
.A2(n_1240),
.B1(n_1238),
.B2(n_1210),
.Y(n_1351)
);

OAI211xp5_ASAP7_75t_SL g1352 ( 
.A1(n_1343),
.A2(n_1240),
.B(n_1193),
.C(n_1210),
.Y(n_1352)
);

INVxp33_ASAP7_75t_L g1353 ( 
.A(n_1344),
.Y(n_1353)
);

NOR2xp67_ASAP7_75t_L g1354 ( 
.A(n_1353),
.B(n_1348),
.Y(n_1354)
);

OAI221xp5_ASAP7_75t_L g1355 ( 
.A1(n_1352),
.A2(n_1347),
.B1(n_1346),
.B2(n_1350),
.C(n_1349),
.Y(n_1355)
);

AOI31xp33_ASAP7_75t_SL g1356 ( 
.A1(n_1351),
.A2(n_1259),
.A3(n_1198),
.B(n_1280),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1354),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1356),
.Y(n_1358)
);

OA22x2_ASAP7_75t_L g1359 ( 
.A1(n_1358),
.A2(n_1355),
.B1(n_1242),
.B2(n_1243),
.Y(n_1359)
);

AO22x2_ASAP7_75t_L g1360 ( 
.A1(n_1357),
.A2(n_1172),
.B1(n_1142),
.B2(n_1133),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1357),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1361),
.Y(n_1362)
);

OAI31xp33_ASAP7_75t_L g1363 ( 
.A1(n_1360),
.A2(n_1179),
.A3(n_1173),
.B(n_1182),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1359),
.B(n_1301),
.Y(n_1364)
);

AOI221xp5_ASAP7_75t_L g1365 ( 
.A1(n_1362),
.A2(n_1198),
.B1(n_1247),
.B2(n_1166),
.C(n_1163),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1365),
.B(n_1363),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1366),
.B(n_1364),
.Y(n_1367)
);

AOI322xp5_ASAP7_75t_L g1368 ( 
.A1(n_1367),
.A2(n_1271),
.A3(n_1270),
.B1(n_1185),
.B2(n_1252),
.C1(n_1193),
.C2(n_1153),
.Y(n_1368)
);

OR2x6_ASAP7_75t_L g1369 ( 
.A(n_1368),
.B(n_1173),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1369),
.A2(n_1247),
.B1(n_1185),
.B2(n_1132),
.Y(n_1370)
);


endmodule