module fake_jpeg_28906_n_384 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_384);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_384;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_8),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_54),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_8),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_48),
.B(n_39),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g88 ( 
.A(n_52),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_53),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_18),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_76),
.Y(n_120)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_38),
.B(n_7),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_24),
.Y(n_80)
);

NAND2xp33_ASAP7_75t_SL g108 ( 
.A(n_80),
.B(n_84),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

AO22x1_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_29),
.B1(n_26),
.B2(n_24),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_91),
.B(n_29),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_82),
.B1(n_81),
.B2(n_77),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_110),
.B1(n_118),
.B2(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_76),
.B(n_39),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_102),
.B(n_112),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_55),
.A2(n_62),
.B1(n_80),
.B2(n_68),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_21),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_21),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_49),
.A2(n_32),
.B1(n_37),
.B2(n_28),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_57),
.A2(n_32),
.B1(n_37),
.B2(n_28),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_65),
.A2(n_32),
.B1(n_43),
.B2(n_35),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_128),
.A2(n_43),
.B1(n_35),
.B2(n_34),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_130),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_89),
.B(n_91),
.C(n_106),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_133),
.B(n_150),
.Y(n_163)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_140),
.B1(n_158),
.B2(n_160),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_108),
.A2(n_83),
.B1(n_66),
.B2(n_56),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_138),
.A2(n_152),
.B1(n_155),
.B2(n_157),
.Y(n_177)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_139),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_118),
.A2(n_60),
.B1(n_20),
.B2(n_34),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_142),
.Y(n_169)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_144),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_89),
.B(n_27),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_35),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_154),
.Y(n_179)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_147),
.Y(n_173)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_149),
.Y(n_178)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_107),
.Y(n_151)
);

BUFx24_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_103),
.A2(n_27),
.B1(n_34),
.B2(n_40),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_153),
.Y(n_164)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_97),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_159),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_27),
.B1(n_40),
.B2(n_75),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_111),
.A2(n_25),
.B1(n_42),
.B2(n_36),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_92),
.B1(n_119),
.B2(n_126),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_125),
.B(n_25),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_26),
.B(n_42),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_94),
.C(n_113),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_135),
.C(n_96),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_170),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_175),
.A2(n_161),
.B1(n_99),
.B2(n_146),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_132),
.A2(n_128),
.B1(n_119),
.B2(n_126),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_180),
.A2(n_160),
.B1(n_159),
.B2(n_156),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_145),
.A2(n_43),
.B(n_110),
.C(n_88),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_182),
.A2(n_98),
.B(n_142),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_184),
.A2(n_185),
.B1(n_187),
.B2(n_200),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_177),
.A2(n_130),
.B1(n_139),
.B2(n_143),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_160),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_186),
.B(n_190),
.Y(n_218)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_150),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_180),
.A2(n_151),
.B1(n_148),
.B2(n_134),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_175),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_98),
.B(n_149),
.Y(n_192)
);

O2A1O1Ixp33_ASAP7_75t_SL g205 ( 
.A1(n_192),
.A2(n_194),
.B(n_196),
.C(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_182),
.A2(n_154),
.B(n_153),
.Y(n_194)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_168),
.Y(n_209)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_172),
.A2(n_75),
.B1(n_73),
.B2(n_51),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_171),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_203),
.B(n_216),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_204),
.A2(n_205),
.B(n_192),
.Y(n_220)
);

AO21x2_ASAP7_75t_L g206 ( 
.A1(n_196),
.A2(n_163),
.B(n_172),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_SL g224 ( 
.A1(n_206),
.A2(n_214),
.B(n_191),
.C(n_197),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_187),
.A2(n_188),
.B1(n_193),
.B2(n_186),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_184),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_209),
.B(n_173),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_201),
.A2(n_163),
.B1(n_169),
.B2(n_171),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_210),
.A2(n_173),
.B1(n_184),
.B2(n_165),
.Y(n_226)
);

OAI22x1_ASAP7_75t_SL g214 ( 
.A1(n_194),
.A2(n_169),
.B1(n_170),
.B2(n_166),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_199),
.B(n_136),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_198),
.B(n_190),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_216),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_205),
.B(n_206),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_214),
.A2(n_194),
.B(n_197),
.Y(n_221)
);

AO21x1_ASAP7_75t_L g244 ( 
.A1(n_221),
.A2(n_224),
.B(n_206),
.Y(n_244)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

AO22x1_ASAP7_75t_L g223 ( 
.A1(n_206),
.A2(n_191),
.B1(n_200),
.B2(n_185),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_223),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_225),
.B(n_229),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_226),
.A2(n_204),
.B1(n_207),
.B2(n_195),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_215),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_227),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_231),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_209),
.B(n_88),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

FAx1_ASAP7_75t_SL g231 ( 
.A(n_208),
.B(n_164),
.CI(n_165),
.CON(n_231),
.SN(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_217),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_212),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.Y(n_240)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_164),
.C(n_166),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_207),
.Y(n_241)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_239),
.A2(n_220),
.B(n_221),
.Y(n_255)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_226),
.C(n_224),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_206),
.B1(n_205),
.B2(n_213),
.Y(n_242)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_250),
.Y(n_260)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_245),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_234),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_248),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_249),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_235),
.B(n_227),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_36),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_262),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_225),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_259),
.Y(n_293)
);

A2O1A1O1Ixp25_ASAP7_75t_L g259 ( 
.A1(n_239),
.A2(n_224),
.B(n_223),
.C(n_229),
.D(n_231),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_231),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_261),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_224),
.B(n_228),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_236),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_267),
.Y(n_278)
);

OA22x2_ASAP7_75t_L g268 ( 
.A1(n_247),
.A2(n_224),
.B1(n_204),
.B2(n_195),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_274),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_249),
.Y(n_269)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

HAxp5_ASAP7_75t_SL g270 ( 
.A(n_246),
.B(n_232),
.CON(n_270),
.SN(n_270)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_270),
.A2(n_174),
.B(n_1),
.Y(n_295)
);

A2O1A1O1Ixp25_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_174),
.B(n_202),
.C(n_181),
.D(n_52),
.Y(n_271)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_167),
.B1(n_176),
.B2(n_181),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_202),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_241),
.C(n_267),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_277),
.C(n_279),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_263),
.A2(n_254),
.B1(n_251),
.B2(n_243),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_276),
.A2(n_280),
.B1(n_287),
.B2(n_174),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_250),
.C(n_245),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_254),
.C(n_251),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_243),
.B1(n_247),
.B2(n_248),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_202),
.C(n_189),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_281),
.B(n_282),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_181),
.C(n_167),
.Y(n_282)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_283),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_174),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_268),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_264),
.A2(n_176),
.B1(n_147),
.B2(n_131),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_286),
.A2(n_271),
.B1(n_268),
.B2(n_121),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_261),
.A2(n_176),
.B1(n_17),
.B2(n_18),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_176),
.C(n_127),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_294),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_129),
.C(n_121),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_295),
.B(n_174),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_269),
.A2(n_272),
.B(n_256),
.Y(n_296)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_296),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_291),
.A2(n_268),
.B1(n_259),
.B2(n_270),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_298),
.B(n_302),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_257),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_306),
.Y(n_324)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_274),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_305),
.B(n_308),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_288),
.A2(n_292),
.B1(n_289),
.B2(n_291),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_281),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_307),
.B(n_311),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_309),
.A2(n_303),
.B1(n_302),
.B2(n_297),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_285),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_275),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_312),
.B(n_316),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_277),
.A2(n_67),
.B1(n_79),
.B2(n_72),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_313),
.B(n_314),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_284),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_282),
.A2(n_13),
.B(n_15),
.Y(n_315)
);

AO21x1_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_10),
.B(n_9),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_293),
.A2(n_10),
.B1(n_18),
.B2(n_17),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_290),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_317),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_305),
.Y(n_319)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_319),
.Y(n_335)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_320),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_304),
.A2(n_294),
.B1(n_293),
.B2(n_3),
.Y(n_323)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_323),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_84),
.C(n_9),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_328),
.B(n_332),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_310),
.B(n_52),
.C(n_85),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_29),
.C(n_2),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_330),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_299),
.C(n_313),
.Y(n_332)
);

MAJx2_ASAP7_75t_L g333 ( 
.A(n_298),
.B(n_6),
.C(n_16),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_333),
.B(n_320),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_326),
.B(n_316),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_334),
.B(n_341),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_336),
.B(n_343),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_308),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_337),
.B(n_342),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_321),
.A2(n_7),
.B(n_16),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_339),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_7),
.C(n_16),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_322),
.B(n_5),
.Y(n_342)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_325),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_346),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_335),
.Y(n_349)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_349),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_338),
.B(n_324),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_351),
.B(n_352),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_336),
.B(n_318),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_342),
.B(n_331),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_354),
.B(n_343),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_345),
.Y(n_355)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_355),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_340),
.B(n_329),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_356),
.B(n_357),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_344),
.B(n_327),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_353),
.B(n_333),
.Y(n_359)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_359),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_348),
.B(n_337),
.Y(n_361)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_361),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_363),
.B(n_365),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_358),
.B(n_339),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_349),
.A2(n_323),
.B(n_5),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_367),
.B(n_347),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_370),
.B(n_372),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_355),
.Y(n_372)
);

OAI21x1_ASAP7_75t_SL g373 ( 
.A1(n_362),
.A2(n_360),
.B(n_364),
.Y(n_373)
);

OAI21x1_ASAP7_75t_L g376 ( 
.A1(n_373),
.A2(n_5),
.B(n_10),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_371),
.B(n_366),
.C(n_350),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_375),
.B(n_369),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_376),
.A2(n_377),
.B(n_15),
.Y(n_379)
);

AOI21xp33_ASAP7_75t_L g377 ( 
.A1(n_368),
.A2(n_15),
.B(n_2),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_378),
.B(n_379),
.C(n_374),
.Y(n_380)
);

BUFx24_ASAP7_75t_SL g381 ( 
.A(n_380),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_381),
.A2(n_0),
.B(n_3),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_382),
.A2(n_0),
.B(n_4),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_383),
.B(n_0),
.Y(n_384)
);


endmodule