module real_aes_1173_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_746;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_0), .B(n_134), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_1), .A2(n_143), .B(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_2), .B(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_3), .B(n_134), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_4), .B(n_150), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_5), .B(n_150), .Y(n_514) );
INVx1_ASAP7_75t_L g141 ( .A(n_6), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_7), .B(n_150), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g791 ( .A(n_8), .Y(n_791) );
NAND2xp33_ASAP7_75t_L g495 ( .A(n_9), .B(n_152), .Y(n_495) );
AND2x2_ASAP7_75t_L g170 ( .A(n_10), .B(n_159), .Y(n_170) );
AND2x2_ASAP7_75t_L g179 ( .A(n_11), .B(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g156 ( .A(n_12), .Y(n_156) );
AOI221x1_ASAP7_75t_L g536 ( .A1(n_13), .A2(n_25), .B1(n_134), .B2(n_143), .C(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_14), .B(n_150), .Y(n_189) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_15), .Y(n_115) );
AND3x1_ASAP7_75t_L g788 ( .A(n_15), .B(n_38), .C(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_16), .B(n_134), .Y(n_491) );
AO21x2_ASAP7_75t_L g489 ( .A1(n_17), .A2(n_159), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_18), .B(n_154), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_19), .B(n_150), .Y(n_474) );
AO21x1_ASAP7_75t_L g509 ( .A1(n_20), .A2(n_134), .B(n_510), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_21), .Y(n_793) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_22), .B(n_134), .Y(n_204) );
INVx1_ASAP7_75t_L g119 ( .A(n_23), .Y(n_119) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_24), .A2(n_90), .B1(n_134), .B2(n_243), .Y(n_242) );
NAND2x1_ASAP7_75t_L g523 ( .A(n_26), .B(n_150), .Y(n_523) );
NAND2x1_ASAP7_75t_L g484 ( .A(n_27), .B(n_152), .Y(n_484) );
OR2x2_ASAP7_75t_L g157 ( .A(n_28), .B(n_87), .Y(n_157) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_28), .A2(n_87), .B(n_156), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_29), .B(n_152), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_30), .B(n_150), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_31), .Y(n_121) );
AO21x2_ASAP7_75t_L g184 ( .A1(n_32), .A2(n_180), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_33), .B(n_152), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_34), .A2(n_143), .B(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_35), .B(n_150), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_36), .A2(n_143), .B(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g140 ( .A(n_37), .B(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g144 ( .A(n_37), .B(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g251 ( .A(n_37), .Y(n_251) );
OR2x6_ASAP7_75t_L g117 ( .A(n_38), .B(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_39), .B(n_134), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_40), .B(n_134), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_41), .B(n_150), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_42), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_43), .B(n_152), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_44), .B(n_134), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_45), .A2(n_143), .B(n_175), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_46), .A2(n_143), .B(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_47), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_48), .B(n_152), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_49), .B(n_134), .Y(n_186) );
INVx1_ASAP7_75t_L g137 ( .A(n_50), .Y(n_137) );
INVx1_ASAP7_75t_L g147 ( .A(n_50), .Y(n_147) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_51), .A2(n_67), .B1(n_777), .B2(n_778), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_51), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_52), .B(n_150), .Y(n_177) );
AND2x2_ASAP7_75t_L g215 ( .A(n_53), .B(n_154), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_54), .B(n_152), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_55), .B(n_150), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_56), .B(n_152), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_57), .A2(n_143), .B(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_58), .B(n_134), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_59), .B(n_134), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_60), .A2(n_143), .B(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g210 ( .A(n_61), .B(n_155), .Y(n_210) );
AO21x1_ASAP7_75t_L g511 ( .A1(n_62), .A2(n_143), .B(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_63), .B(n_134), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_64), .A2(n_81), .B1(n_757), .B2(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_64), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_65), .B(n_152), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_66), .B(n_134), .Y(n_486) );
INVx1_ASAP7_75t_L g778 ( .A(n_67), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_68), .B(n_152), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_69), .A2(n_95), .B1(n_143), .B2(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_70), .B(n_150), .Y(n_207) );
AND2x2_ASAP7_75t_L g559 ( .A(n_71), .B(n_155), .Y(n_559) );
INVx1_ASAP7_75t_L g139 ( .A(n_72), .Y(n_139) );
INVx1_ASAP7_75t_L g145 ( .A(n_72), .Y(n_145) );
AND2x2_ASAP7_75t_L g487 ( .A(n_73), .B(n_180), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_74), .B(n_152), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_75), .A2(n_143), .B(n_219), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_76), .A2(n_143), .B(n_148), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_77), .A2(n_143), .B(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g201 ( .A(n_78), .B(n_155), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_79), .B(n_154), .Y(n_240) );
INVx1_ASAP7_75t_L g120 ( .A(n_80), .Y(n_120) );
INVx1_ASAP7_75t_L g758 ( .A(n_81), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_82), .B(n_134), .Y(n_476) );
AND2x2_ASAP7_75t_L g497 ( .A(n_83), .B(n_180), .Y(n_497) );
AOI22xp33_ASAP7_75t_SL g759 ( .A1(n_84), .A2(n_756), .B1(n_760), .B2(n_764), .Y(n_759) );
AND2x2_ASAP7_75t_L g158 ( .A(n_85), .B(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g510 ( .A(n_86), .B(n_191), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_88), .B(n_152), .Y(n_475) );
AND2x2_ASAP7_75t_L g526 ( .A(n_89), .B(n_180), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_91), .B(n_150), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_92), .A2(n_143), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_93), .B(n_152), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_94), .A2(n_143), .B(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_96), .B(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_97), .B(n_150), .Y(n_502) );
BUFx2_ASAP7_75t_L g209 ( .A(n_98), .Y(n_209) );
BUFx2_ASAP7_75t_L g107 ( .A(n_99), .Y(n_107) );
BUFx2_ASAP7_75t_SL g772 ( .A(n_99), .Y(n_772) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_100), .A2(n_143), .B(n_493), .Y(n_492) );
AOI21xp33_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_782), .B(n_792), .Y(n_101) );
OA21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_122), .B(n_768), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_108), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g773 ( .A1(n_109), .A2(n_774), .B(n_780), .Y(n_773) );
NOR2xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_121), .Y(n_109) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g781 ( .A(n_114), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AND2x6_ASAP7_75t_SL g461 ( .A(n_115), .B(n_117), .Y(n_461) );
OR2x6_ASAP7_75t_SL g755 ( .A(n_115), .B(n_116), .Y(n_755) );
OR2x2_ASAP7_75t_L g767 ( .A(n_115), .B(n_117), .Y(n_767) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g787 ( .A(n_118), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
OAI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_756), .B(n_759), .Y(n_122) );
INVxp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_460), .B1(n_462), .B2(n_753), .Y(n_124) );
INVx1_ASAP7_75t_L g761 ( .A(n_125), .Y(n_761) );
OAI22xp5_ASAP7_75t_SL g774 ( .A1(n_125), .A2(n_775), .B1(n_776), .B2(n_779), .Y(n_774) );
INVx5_ASAP7_75t_L g775 ( .A(n_125), .Y(n_775) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_364), .Y(n_125) );
NOR3xp33_ASAP7_75t_L g126 ( .A(n_127), .B(n_289), .C(n_325), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_263), .Y(n_127) );
AOI211xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_181), .B(n_211), .C(n_236), .Y(n_128) );
AND2x2_ASAP7_75t_L g354 ( .A(n_129), .B(n_213), .Y(n_354) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_161), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_130), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g387 ( .A(n_130), .B(n_269), .Y(n_387) );
AND2x2_ASAP7_75t_L g403 ( .A(n_130), .B(n_228), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_130), .B(n_413), .Y(n_412) );
NAND2x1p5_ASAP7_75t_L g436 ( .A(n_130), .B(n_437), .Y(n_436) );
INVx4_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x4_ASAP7_75t_SL g223 ( .A(n_131), .B(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g258 ( .A(n_131), .Y(n_258) );
AND2x2_ASAP7_75t_L g305 ( .A(n_131), .B(n_238), .Y(n_305) );
AND2x2_ASAP7_75t_L g324 ( .A(n_131), .B(n_161), .Y(n_324) );
BUFx2_ASAP7_75t_L g329 ( .A(n_131), .Y(n_329) );
AND2x2_ASAP7_75t_L g373 ( .A(n_131), .B(n_171), .Y(n_373) );
AND2x4_ASAP7_75t_L g445 ( .A(n_131), .B(n_446), .Y(n_445) );
NOR2x1_ASAP7_75t_L g457 ( .A(n_131), .B(n_227), .Y(n_457) );
OR2x6_ASAP7_75t_L g131 ( .A(n_132), .B(n_158), .Y(n_131) );
AOI21xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_142), .B(n_154), .Y(n_132) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_140), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
AND2x6_ASAP7_75t_L g152 ( .A(n_136), .B(n_145), .Y(n_152) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g150 ( .A(n_138), .B(n_147), .Y(n_150) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx5_ASAP7_75t_L g153 ( .A(n_140), .Y(n_153) );
AND2x2_ASAP7_75t_L g146 ( .A(n_141), .B(n_147), .Y(n_146) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_141), .Y(n_246) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
BUFx3_ASAP7_75t_L g247 ( .A(n_144), .Y(n_247) );
INVx2_ASAP7_75t_L g253 ( .A(n_145), .Y(n_253) );
AND2x4_ASAP7_75t_L g249 ( .A(n_146), .B(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g245 ( .A(n_147), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_151), .B(n_153), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_152), .B(n_209), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_153), .A2(n_167), .B(n_168), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_153), .A2(n_176), .B(n_177), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_153), .A2(n_189), .B(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_153), .A2(n_198), .B(n_199), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_153), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_153), .A2(n_220), .B(n_221), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_153), .A2(n_474), .B(n_475), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_153), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_153), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_153), .A2(n_502), .B(n_503), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_153), .A2(n_513), .B(n_514), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_153), .A2(n_523), .B(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_153), .A2(n_538), .B(n_539), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_153), .A2(n_556), .B(n_557), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_154), .Y(n_163) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_154), .A2(n_242), .B(n_248), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_154), .A2(n_499), .B(n_500), .Y(n_498) );
OA21x2_ASAP7_75t_L g535 ( .A1(n_154), .A2(n_536), .B(n_540), .Y(n_535) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_154), .A2(n_536), .B(n_540), .Y(n_547) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AND2x2_ASAP7_75t_SL g155 ( .A(n_156), .B(n_157), .Y(n_155) );
AND2x4_ASAP7_75t_L g191 ( .A(n_156), .B(n_157), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_159), .A2(n_204), .B(n_205), .Y(n_203) );
BUFx4f_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g172 ( .A(n_160), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_161), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g376 ( .A(n_161), .Y(n_376) );
BUFx2_ASAP7_75t_L g425 ( .A(n_161), .Y(n_425) );
INVx1_ASAP7_75t_L g447 ( .A(n_161), .Y(n_447) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_171), .Y(n_161) );
INVx3_ASAP7_75t_L g224 ( .A(n_162), .Y(n_224) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_162), .Y(n_413) );
AOI21x1_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_170), .Y(n_162) );
AO21x2_ASAP7_75t_L g480 ( .A1(n_163), .A2(n_481), .B(n_487), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_165), .B(n_169), .Y(n_164) );
INVx2_ASAP7_75t_L g227 ( .A(n_171), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_171), .B(n_224), .Y(n_228) );
INVx2_ASAP7_75t_L g313 ( .A(n_171), .Y(n_313) );
OR2x2_ASAP7_75t_L g320 ( .A(n_171), .B(n_269), .Y(n_320) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_179), .Y(n_171) );
INVx4_ASAP7_75t_L g180 ( .A(n_172), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_174), .B(n_178), .Y(n_173) );
INVx3_ASAP7_75t_L g194 ( .A(n_180), .Y(n_194) );
AND2x2_ASAP7_75t_L g275 ( .A(n_181), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g309 ( .A(n_181), .B(n_272), .Y(n_309) );
AND2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_192), .Y(n_181) );
AND2x2_ASAP7_75t_L g345 ( .A(n_182), .B(n_234), .Y(n_345) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g302 ( .A(n_183), .B(n_193), .Y(n_302) );
AND2x2_ASAP7_75t_L g421 ( .A(n_183), .B(n_202), .Y(n_421) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g233 ( .A(n_184), .Y(n_233) );
INVx1_ASAP7_75t_L g261 ( .A(n_184), .Y(n_261) );
AND2x2_ASAP7_75t_L g317 ( .A(n_184), .B(n_193), .Y(n_317) );
AND2x2_ASAP7_75t_L g322 ( .A(n_184), .B(n_214), .Y(n_322) );
OR2x2_ASAP7_75t_L g385 ( .A(n_184), .B(n_202), .Y(n_385) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_184), .Y(n_394) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_191), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_191), .A2(n_217), .B(n_218), .Y(n_216) );
INVx1_ASAP7_75t_SL g470 ( .A(n_191), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_191), .A2(n_491), .B(n_492), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_191), .B(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g213 ( .A(n_192), .B(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g262 ( .A(n_192), .Y(n_262) );
NOR2x1_ASAP7_75t_SL g192 ( .A(n_193), .B(n_202), .Y(n_192) );
AO21x1_ASAP7_75t_SL g193 ( .A1(n_194), .A2(n_195), .B(n_201), .Y(n_193) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_194), .A2(n_195), .B(n_201), .Y(n_235) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_194), .A2(n_520), .B(n_526), .Y(n_519) );
AO21x2_ASAP7_75t_L g552 ( .A1(n_194), .A2(n_553), .B(n_559), .Y(n_552) );
AO21x2_ASAP7_75t_L g588 ( .A1(n_194), .A2(n_553), .B(n_559), .Y(n_588) );
AO21x2_ASAP7_75t_L g591 ( .A1(n_194), .A2(n_520), .B(n_526), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_200), .Y(n_195) );
AND2x2_ASAP7_75t_L g230 ( .A(n_202), .B(n_231), .Y(n_230) );
INVx2_ASAP7_75t_SL g288 ( .A(n_202), .Y(n_288) );
NAND2x1_ASAP7_75t_L g298 ( .A(n_202), .B(n_214), .Y(n_298) );
OR2x2_ASAP7_75t_L g303 ( .A(n_202), .B(n_231), .Y(n_303) );
BUFx2_ASAP7_75t_L g359 ( .A(n_202), .Y(n_359) );
AND2x2_ASAP7_75t_L g395 ( .A(n_202), .B(n_274), .Y(n_395) );
AND2x2_ASAP7_75t_L g406 ( .A(n_202), .B(n_234), .Y(n_406) );
OR2x6_ASAP7_75t_L g202 ( .A(n_203), .B(n_210), .Y(n_202) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_222), .B1(n_228), .B2(n_229), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_213), .A2(n_403), .B1(n_453), .B2(n_458), .Y(n_452) );
INVx4_ASAP7_75t_L g231 ( .A(n_214), .Y(n_231) );
INVx2_ASAP7_75t_L g272 ( .A(n_214), .Y(n_272) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_214), .Y(n_343) );
OR2x2_ASAP7_75t_L g358 ( .A(n_214), .B(n_234), .Y(n_358) );
OR2x2_ASAP7_75t_SL g384 ( .A(n_214), .B(n_385), .Y(n_384) );
OR2x6_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
AND2x2_ASAP7_75t_SL g222 ( .A(n_223), .B(n_225), .Y(n_222) );
INVx2_ASAP7_75t_SL g265 ( .A(n_223), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_223), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g333 ( .A(n_223), .B(n_281), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_223), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g255 ( .A(n_224), .Y(n_255) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_224), .Y(n_280) );
AND2x2_ASAP7_75t_L g336 ( .A(n_224), .B(n_313), .Y(n_336) );
INVx1_ASAP7_75t_L g446 ( .A(n_224), .Y(n_446) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_226), .B(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_226), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g254 ( .A(n_227), .B(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_228), .B(n_387), .Y(n_386) );
AOI321xp33_ASAP7_75t_L g408 ( .A1(n_229), .A2(n_310), .A3(n_378), .B1(n_409), .B2(n_410), .C(n_414), .Y(n_408) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_232), .Y(n_229) );
INVxp67_ASAP7_75t_SL g307 ( .A(n_230), .Y(n_307) );
AND2x2_ASAP7_75t_L g332 ( .A(n_230), .B(n_261), .Y(n_332) );
AND2x2_ASAP7_75t_L g407 ( .A(n_230), .B(n_317), .Y(n_407) );
INVx1_ASAP7_75t_L g276 ( .A(n_231), .Y(n_276) );
BUFx2_ASAP7_75t_L g286 ( .A(n_231), .Y(n_286) );
NOR2xp67_ASAP7_75t_L g393 ( .A(n_231), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g331 ( .A(n_232), .Y(n_331) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
BUFx2_ASAP7_75t_L g338 ( .A(n_233), .Y(n_338) );
INVx2_ASAP7_75t_L g274 ( .A(n_234), .Y(n_274) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_234), .Y(n_297) );
INVx3_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AOI21xp33_ASAP7_75t_SL g236 ( .A1(n_237), .A2(n_256), .B(n_259), .Y(n_236) );
NOR2xp67_ASAP7_75t_L g390 ( .A(n_237), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_254), .Y(n_238) );
INVx3_ASAP7_75t_L g281 ( .A(n_239), .Y(n_281) );
AND2x2_ASAP7_75t_L g312 ( .A(n_239), .B(n_313), .Y(n_312) );
AND2x4_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
AND2x4_ASAP7_75t_L g269 ( .A(n_240), .B(n_241), .Y(n_269) );
AND2x4_ASAP7_75t_L g243 ( .A(n_244), .B(n_247), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
NOR2x1p5_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g352 ( .A(n_254), .Y(n_352) );
INVx1_ASAP7_75t_SL g437 ( .A(n_255), .Y(n_437) );
INVxp33_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_258), .B(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g363 ( .A(n_258), .B(n_320), .Y(n_363) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
AND2x2_ASAP7_75t_L g367 ( .A(n_260), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_260), .B(n_382), .Y(n_381) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_261), .B(n_298), .Y(n_353) );
NOR4xp25_ASAP7_75t_L g448 ( .A(n_261), .B(n_292), .C(n_449), .D(n_450), .Y(n_448) );
OR2x2_ASAP7_75t_L g416 ( .A(n_262), .B(n_417), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_270), .B1(n_275), .B2(n_277), .C(n_282), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
AND2x2_ASAP7_75t_L g291 ( .A(n_266), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g328 ( .A(n_267), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g348 ( .A(n_268), .Y(n_348) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx3_ASAP7_75t_L g371 ( .A(n_269), .Y(n_371) );
AND2x2_ASAP7_75t_L g378 ( .A(n_269), .B(n_379), .Y(n_378) );
INVxp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
OR2x2_ASAP7_75t_L g315 ( .A(n_272), .B(n_316), .Y(n_315) );
INVxp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_274), .B(n_288), .Y(n_287) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx2_ASAP7_75t_L g292 ( .A(n_279), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_279), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g284 ( .A(n_281), .Y(n_284) );
OAI321xp33_ASAP7_75t_L g396 ( .A1(n_281), .A2(n_389), .A3(n_397), .B1(n_402), .B2(n_404), .C(n_408), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
OR2x2_ASAP7_75t_L g351 ( .A(n_284), .B(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g451 ( .A(n_287), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_288), .B(n_331), .Y(n_330) );
NAND2xp33_ASAP7_75t_SL g431 ( .A(n_288), .B(n_302), .Y(n_431) );
OAI211xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_293), .B(n_304), .C(n_308), .Y(n_289) );
INVxp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2x1_ASAP7_75t_L g293 ( .A(n_294), .B(n_299), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g400 ( .A(n_297), .Y(n_400) );
INVx3_ASAP7_75t_L g339 ( .A(n_298), .Y(n_339) );
OR2x2_ASAP7_75t_L g442 ( .A(n_298), .B(n_316), .Y(n_442) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_300), .A2(n_384), .B1(n_386), .B2(n_388), .Y(n_383) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_SL g382 ( .A(n_303), .Y(n_382) );
OR2x2_ASAP7_75t_L g459 ( .A(n_303), .B(n_316), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AOI21xp5_ASAP7_75t_SL g308 ( .A1(n_309), .A2(n_310), .B(n_314), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_312), .B(n_329), .Y(n_428) );
AND2x2_ASAP7_75t_L g434 ( .A(n_312), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g379 ( .A(n_313), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_318), .B1(n_321), .B2(n_323), .Y(n_314) );
A2O1A1Ixp33_ASAP7_75t_L g360 ( .A1(n_316), .A2(n_359), .B(n_361), .C(n_363), .Y(n_360) );
INVx2_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_319), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_319), .B(n_411), .Y(n_433) );
INVx2_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g405 ( .A(n_322), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
A2O1A1Ixp33_ASAP7_75t_L g355 ( .A1(n_324), .A2(n_356), .B(n_359), .C(n_360), .Y(n_355) );
NAND3xp33_ASAP7_75t_SL g325 ( .A(n_326), .B(n_340), .C(n_355), .Y(n_325) );
AOI222xp33_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_330), .B1(n_332), .B2(n_333), .C1(n_334), .C2(n_337), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g389 ( .A(n_329), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_329), .B(n_362), .Y(n_415) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_SL g349 ( .A(n_336), .Y(n_349) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
OR2x2_ASAP7_75t_L g454 ( .A(n_338), .B(n_371), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_339), .A2(n_430), .B1(n_432), .B2(n_434), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_346), .B1(n_350), .B2(n_353), .C(n_354), .Y(n_340) );
INVx2_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI21xp5_ASAP7_75t_SL g414 ( .A1(n_347), .A2(n_415), .B(n_416), .Y(n_414) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx2_ASAP7_75t_L g362 ( .A(n_348), .Y(n_362) );
AND2x2_ASAP7_75t_L g456 ( .A(n_348), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g440 ( .A(n_352), .Y(n_440) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g369 ( .A(n_358), .B(n_359), .Y(n_369) );
INVx1_ASAP7_75t_L g422 ( .A(n_358), .Y(n_422) );
NOR3xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_396), .C(n_418), .Y(n_364) );
OAI211xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_370), .B(n_372), .C(n_377), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI21xp33_ASAP7_75t_L g372 ( .A1(n_367), .A2(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI211xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_380), .B(n_383), .C(n_390), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g401 ( .A(n_384), .Y(n_401) );
INVxp67_ASAP7_75t_SL g426 ( .A(n_385), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_387), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g449 ( .A(n_387), .Y(n_449) );
AND2x2_ASAP7_75t_L g439 ( .A(n_389), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g409 ( .A(n_391), .Y(n_409) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
INVx1_ASAP7_75t_L g417 ( .A(n_393), .Y(n_417) );
INVx2_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_399), .B(n_401), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g438 ( .A1(n_405), .A2(n_439), .B1(n_441), .B2(n_443), .C(n_448), .Y(n_438) );
OAI21xp33_ASAP7_75t_SL g453 ( .A1(n_410), .A2(n_454), .B(n_455), .Y(n_453) );
INVx2_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND4xp25_ASAP7_75t_L g418 ( .A(n_419), .B(n_429), .C(n_438), .D(n_452), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_423), .B1(n_426), .B2(n_427), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_447), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx3_ASAP7_75t_SL g763 ( .A(n_460), .Y(n_763) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_463), .A2(n_755), .B1(n_761), .B2(n_762), .Y(n_760) );
OR2x6_ASAP7_75t_L g463 ( .A(n_464), .B(n_651), .Y(n_463) );
NAND3xp33_ASAP7_75t_SL g464 ( .A(n_465), .B(n_563), .C(n_618), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_504), .B1(n_527), .B2(n_531), .C(n_541), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_488), .Y(n_466) );
AND2x2_ASAP7_75t_SL g529 ( .A(n_467), .B(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g562 ( .A(n_467), .Y(n_562) );
AND2x2_ASAP7_75t_L g607 ( .A(n_467), .B(n_544), .Y(n_607) );
AND2x4_ASAP7_75t_L g467 ( .A(n_468), .B(n_479), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g595 ( .A(n_469), .Y(n_595) );
INVx1_ASAP7_75t_L g605 ( .A(n_469), .Y(n_605) );
AO21x2_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B(n_477), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_470), .B(n_478), .Y(n_477) );
AO21x2_ASAP7_75t_L g569 ( .A1(n_470), .A2(n_471), .B(n_477), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_476), .Y(n_471) );
OR2x2_ASAP7_75t_L g584 ( .A(n_479), .B(n_489), .Y(n_584) );
NAND2x1p5_ASAP7_75t_L g615 ( .A(n_479), .B(n_530), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_479), .B(n_496), .Y(n_628) );
INVx2_ASAP7_75t_L g637 ( .A(n_479), .Y(n_637) );
AND2x2_ASAP7_75t_L g658 ( .A(n_479), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g742 ( .A(n_479), .B(n_561), .Y(n_742) );
INVx4_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g570 ( .A(n_480), .B(n_496), .Y(n_570) );
AND2x2_ASAP7_75t_L g703 ( .A(n_480), .B(n_530), .Y(n_703) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_480), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_486), .Y(n_481) );
AND2x4_ASAP7_75t_L g657 ( .A(n_488), .B(n_658), .Y(n_657) );
AOI321xp33_ASAP7_75t_L g671 ( .A1(n_488), .A2(n_600), .A3(n_601), .B1(n_633), .B2(n_672), .C(n_675), .Y(n_671) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_496), .Y(n_488) );
BUFx3_ASAP7_75t_L g528 ( .A(n_489), .Y(n_528) );
INVx2_ASAP7_75t_L g561 ( .A(n_489), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_489), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g594 ( .A(n_489), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g627 ( .A(n_489), .Y(n_627) );
INVx5_ASAP7_75t_L g530 ( .A(n_496), .Y(n_530) );
NOR2x1_ASAP7_75t_SL g579 ( .A(n_496), .B(n_569), .Y(n_579) );
BUFx2_ASAP7_75t_L g674 ( .A(n_496), .Y(n_674) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
INVxp67_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_517), .Y(n_505) );
NOR2xp33_ASAP7_75t_SL g572 ( .A(n_506), .B(n_573), .Y(n_572) );
NOR4xp25_ASAP7_75t_L g675 ( .A(n_506), .B(n_669), .C(n_673), .D(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g713 ( .A(n_506), .Y(n_713) );
AND2x2_ASAP7_75t_L g747 ( .A(n_506), .B(n_687), .Y(n_747) );
BUFx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g548 ( .A(n_507), .Y(n_548) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g602 ( .A(n_508), .Y(n_602) );
OAI21x1_ASAP7_75t_SL g508 ( .A1(n_509), .A2(n_511), .B(n_515), .Y(n_508) );
INVx1_ASAP7_75t_L g516 ( .A(n_510), .Y(n_516) );
AOI33xp33_ASAP7_75t_L g743 ( .A1(n_517), .A2(n_545), .A3(n_576), .B1(n_592), .B2(n_698), .B3(n_744), .Y(n_743) );
INVx1_ASAP7_75t_SL g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g533 ( .A(n_518), .B(n_534), .Y(n_533) );
AND2x4_ASAP7_75t_L g543 ( .A(n_518), .B(n_544), .Y(n_543) );
BUFx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g550 ( .A(n_519), .Y(n_550) );
INVxp67_ASAP7_75t_L g631 ( .A(n_519), .Y(n_631) );
AND2x2_ASAP7_75t_L g687 ( .A(n_519), .B(n_552), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_527), .A2(n_709), .B(n_710), .Y(n_708) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
AND2x2_ASAP7_75t_L g696 ( .A(n_528), .B(n_570), .Y(n_696) );
AND3x2_ASAP7_75t_L g698 ( .A(n_528), .B(n_582), .C(n_637), .Y(n_698) );
INVx3_ASAP7_75t_SL g650 ( .A(n_529), .Y(n_650) );
INVx4_ASAP7_75t_L g544 ( .A(n_530), .Y(n_544) );
AND2x2_ASAP7_75t_L g582 ( .A(n_530), .B(n_569), .Y(n_582) );
INVxp67_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx2_ASAP7_75t_L g576 ( .A(n_534), .Y(n_576) );
AND2x4_ASAP7_75t_L g601 ( .A(n_534), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g664 ( .A(n_534), .B(n_552), .Y(n_664) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g634 ( .A(n_535), .Y(n_634) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_535), .Y(n_656) );
O2A1O1Ixp33_ASAP7_75t_R g541 ( .A1(n_542), .A2(n_545), .B(n_549), .C(n_560), .Y(n_541) );
CKINVDCx16_ASAP7_75t_R g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g593 ( .A(n_544), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_544), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_544), .B(n_561), .Y(n_722) );
INVx1_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g704 ( .A(n_546), .B(n_694), .Y(n_704) );
AND2x2_ASAP7_75t_SL g546 ( .A(n_547), .B(n_548), .Y(n_546) );
AND2x2_ASAP7_75t_L g551 ( .A(n_547), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g573 ( .A(n_547), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g589 ( .A(n_547), .B(n_590), .Y(n_589) );
AND2x4_ASAP7_75t_L g622 ( .A(n_547), .B(n_602), .Y(n_622) );
AND2x4_ASAP7_75t_L g587 ( .A(n_548), .B(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g611 ( .A(n_548), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g649 ( .A(n_548), .B(n_574), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
AND2x2_ASAP7_75t_L g577 ( .A(n_550), .B(n_574), .Y(n_577) );
AND2x2_ASAP7_75t_L g592 ( .A(n_550), .B(n_552), .Y(n_592) );
BUFx2_ASAP7_75t_L g648 ( .A(n_550), .Y(n_648) );
AND2x2_ASAP7_75t_L g662 ( .A(n_550), .B(n_573), .Y(n_662) );
INVx2_ASAP7_75t_L g574 ( .A(n_552), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_554), .B(n_558), .Y(n_553) );
OAI22xp33_ASAP7_75t_L g610 ( .A1(n_560), .A2(n_611), .B1(n_613), .B2(n_617), .Y(n_610) );
INVx2_ASAP7_75t_SL g641 ( .A(n_560), .Y(n_641) );
OR2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
AND2x2_ASAP7_75t_L g616 ( .A(n_561), .B(n_569), .Y(n_616) );
INVx1_ASAP7_75t_L g723 ( .A(n_562), .Y(n_723) );
NOR3xp33_ASAP7_75t_L g563 ( .A(n_564), .B(n_596), .C(n_610), .Y(n_563) );
OAI221xp5_ASAP7_75t_SL g564 ( .A1(n_565), .A2(n_571), .B1(n_575), .B2(n_578), .C(n_580), .Y(n_564) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_570), .Y(n_566) );
INVxp67_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g624 ( .A(n_568), .Y(n_624) );
INVxp67_ASAP7_75t_SL g752 ( .A(n_568), .Y(n_752) );
INVx1_ASAP7_75t_L g715 ( .A(n_570), .Y(n_715) );
AND2x2_ASAP7_75t_SL g725 ( .A(n_570), .B(n_594), .Y(n_725) );
INVxp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_574), .B(n_602), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
OR2x2_ASAP7_75t_L g608 ( .A(n_576), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g686 ( .A(n_576), .Y(n_686) );
AND2x2_ASAP7_75t_L g621 ( .A(n_577), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g667 ( .A(n_579), .B(n_627), .Y(n_667) );
AND2x2_ASAP7_75t_L g744 ( .A(n_579), .B(n_742), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_585), .B1(n_592), .B2(n_593), .Y(n_580) );
AND2x4_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g603 ( .A(n_584), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
INVx2_ASAP7_75t_L g609 ( .A(n_587), .Y(n_609) );
AND2x4_ASAP7_75t_L g633 ( .A(n_587), .B(n_634), .Y(n_633) );
OAI21xp33_ASAP7_75t_SL g663 ( .A1(n_587), .A2(n_664), .B(n_665), .Y(n_663) );
AND2x2_ASAP7_75t_L g690 ( .A(n_587), .B(n_648), .Y(n_690) );
INVx2_ASAP7_75t_L g612 ( .A(n_588), .Y(n_612) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_588), .Y(n_645) );
INVx1_ASAP7_75t_SL g669 ( .A(n_589), .Y(n_669) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
BUFx2_ASAP7_75t_L g600 ( .A(n_591), .Y(n_600) );
AND2x4_ASAP7_75t_SL g694 ( .A(n_591), .B(n_612), .Y(n_694) );
AND2x2_ASAP7_75t_L g691 ( .A(n_594), .B(n_637), .Y(n_691) );
AND2x2_ASAP7_75t_L g717 ( .A(n_594), .B(n_703), .Y(n_717) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_595), .Y(n_639) );
INVx1_ASAP7_75t_L g659 ( .A(n_595), .Y(n_659) );
OAI22xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_603), .B1(n_606), .B2(n_608), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_601), .B(n_612), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_601), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g740 ( .A(n_601), .Y(n_740) );
INVx2_ASAP7_75t_SL g665 ( .A(n_603), .Y(n_665) );
AND2x2_ASAP7_75t_L g677 ( .A(n_605), .B(n_637), .Y(n_677) );
INVx2_ASAP7_75t_L g683 ( .A(n_605), .Y(n_683) );
INVxp33_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g642 ( .A(n_608), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_611), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g733 ( .A(n_611), .Y(n_733) );
INVx1_ASAP7_75t_L g661 ( .A(n_613), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_614), .B(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g672 ( .A(n_616), .B(n_673), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_616), .A2(n_746), .B1(n_747), .B2(n_748), .Y(n_745) );
NOR3xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_640), .C(n_643), .Y(n_618) );
OAI221xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_623), .B1(n_625), .B2(n_629), .C(n_632), .Y(n_619) );
INVx1_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g738 ( .A(n_623), .Y(n_738) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g707 ( .A(n_624), .B(n_673), .Y(n_707) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_628), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g638 ( .A(n_627), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g709 ( .A(n_629), .Y(n_709) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx1_ASAP7_75t_L g706 ( .A(n_630), .Y(n_706) );
INVx1_ASAP7_75t_L g712 ( .A(n_631), .Y(n_712) );
OR2x2_ASAP7_75t_L g735 ( .A(n_631), .B(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
INVx1_ASAP7_75t_SL g644 ( .A(n_634), .Y(n_644) );
AND2x2_ASAP7_75t_L g714 ( .A(n_634), .B(n_694), .Y(n_714) );
AND2x2_ASAP7_75t_SL g746 ( .A(n_634), .B(n_647), .Y(n_746) );
INVx1_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
INVx1_ASAP7_75t_L g751 ( .A(n_637), .Y(n_751) );
INVx1_ASAP7_75t_L g701 ( .A(n_639), .Y(n_701) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
O2A1O1Ixp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B(n_646), .C(n_650), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_644), .B(n_694), .Y(n_718) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_647), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
AND2x2_ASAP7_75t_L g655 ( .A(n_649), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g736 ( .A(n_649), .Y(n_736) );
NAND4xp75_ASAP7_75t_L g651 ( .A(n_652), .B(n_708), .C(n_724), .D(n_745), .Y(n_651) );
NOR3x1_ASAP7_75t_L g652 ( .A(n_653), .B(n_670), .C(n_692), .Y(n_652) );
NAND4xp75_ASAP7_75t_L g653 ( .A(n_654), .B(n_660), .C(n_663), .D(n_666), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_655), .B(n_657), .Y(n_654) );
AND2x2_ASAP7_75t_L g705 ( .A(n_656), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g730 ( .A(n_657), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g660 ( .A(n_661), .B(n_662), .Y(n_660) );
INVx1_ASAP7_75t_SL g719 ( .A(n_662), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_678), .Y(n_670) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_674), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_684), .B(n_688), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OAI322xp33_ASAP7_75t_L g710 ( .A1(n_682), .A2(n_711), .A3(n_715), .B1(n_716), .B2(n_718), .C1(n_719), .C2(n_720), .Y(n_710) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_683), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_686), .B(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_687), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
OAI211xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_695), .B(n_697), .C(n_699), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_704), .B1(n_705), .B2(n_707), .Y(n_699) );
NOR2xp33_ASAP7_75t_SL g700 ( .A(n_701), .B(n_702), .Y(n_700) );
INVx2_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_713), .B(n_714), .Y(n_711) );
INVxp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_717), .B(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_721), .B(n_723), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g727 ( .A(n_722), .B(n_728), .Y(n_727) );
O2A1O1Ixp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_726), .B(n_731), .C(n_734), .Y(n_724) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_727), .B(n_730), .Y(n_726) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OAI221xp5_ASAP7_75t_SL g734 ( .A1(n_735), .A2(n_737), .B1(n_739), .B2(n_741), .C(n_743), .Y(n_734) );
INVxp67_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
CKINVDCx11_ASAP7_75t_R g754 ( .A(n_755), .Y(n_754) );
CKINVDCx6p67_ASAP7_75t_R g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_773), .Y(n_768) );
CKINVDCx5p33_ASAP7_75t_R g769 ( .A(n_770), .Y(n_769) );
CKINVDCx11_ASAP7_75t_R g770 ( .A(n_771), .Y(n_770) );
CKINVDCx8_ASAP7_75t_R g771 ( .A(n_772), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_776), .Y(n_779) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_SL g794 ( .A(n_785), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g785 ( .A(n_786), .Y(n_785) );
AND2x2_ASAP7_75t_SL g786 ( .A(n_787), .B(n_788), .Y(n_786) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .Y(n_792) );
endmodule