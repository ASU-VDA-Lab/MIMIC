module fake_jpeg_23248_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx3_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_3),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_23),
.B(n_25),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_4),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_L g27 ( 
.A1(n_11),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_28),
.B1(n_18),
.B2(n_20),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_12),
.A2(n_15),
.B1(n_11),
.B2(n_20),
.Y(n_28)
);

OAI32xp33_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_13),
.A3(n_12),
.B1(n_19),
.B2(n_15),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_29),
.A2(n_30),
.B1(n_33),
.B2(n_40),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_18),
.B1(n_13),
.B2(n_19),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_26),
.B1(n_17),
.B2(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_22),
.B(n_5),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_17),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_39),
.B(n_17),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_6),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_38),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_31),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_44),
.C(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_56),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_32),
.B(n_29),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_54),
.A2(n_55),
.B1(n_51),
.B2(n_45),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_52),
.A2(n_43),
.B1(n_30),
.B2(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_60),
.Y(n_65)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_62),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_47),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_61),
.C(n_60),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_64),
.A2(n_58),
.B(n_42),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_65),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_63),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_64),
.B1(n_33),
.B2(n_40),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_SL g70 ( 
.A1(n_68),
.A2(n_69),
.B(n_39),
.C(n_53),
.Y(n_70)
);

MAJx2_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_39),
.C(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);


endmodule