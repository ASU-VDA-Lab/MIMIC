module real_jpeg_26733_n_17 (n_5, n_4, n_8, n_0, n_12, n_315, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_315;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_0),
.A2(n_34),
.B1(n_35),
.B2(n_54),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_0),
.A2(n_48),
.B1(n_51),
.B2(n_54),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_54),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_1),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_1),
.A2(n_28),
.B1(n_64),
.B2(n_65),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_1),
.A2(n_28),
.B1(n_48),
.B2(n_51),
.Y(n_239)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_2),
.Y(n_84)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_2),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_3),
.A2(n_64),
.B1(n_65),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_3),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_70),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_70),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_3),
.A2(n_48),
.B1(n_51),
.B2(n_70),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_4),
.B(n_35),
.Y(n_149)
);

A2O1A1O1Ixp25_ASAP7_75t_L g151 ( 
.A1(n_4),
.A2(n_35),
.B(n_43),
.C(n_149),
.D(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_4),
.B(n_32),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_4),
.Y(n_181)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_4),
.A2(n_83),
.B(n_166),
.Y(n_186)
);

A2O1A1O1Ixp25_ASAP7_75t_L g198 ( 
.A1(n_4),
.A2(n_30),
.B(n_31),
.C(n_199),
.D(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_4),
.B(n_30),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_4),
.A2(n_29),
.B(n_62),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_4),
.A2(n_64),
.B1(n_65),
.B2(n_181),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_5),
.A2(n_40),
.B1(n_48),
.B2(n_51),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_8),
.A2(n_64),
.B1(n_65),
.B2(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_8),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_8),
.A2(n_48),
.B1(n_51),
.B2(n_135),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_135),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_135),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_10),
.A2(n_64),
.B1(n_65),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_10),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_98),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_10),
.A2(n_48),
.B1(n_51),
.B2(n_98),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_98),
.Y(n_201)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_11),
.B(n_35),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_11),
.A2(n_45),
.B1(n_48),
.B2(n_51),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_11),
.B(n_48),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_12),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_12),
.A2(n_48),
.B1(n_51),
.B2(n_161),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_161),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_12),
.A2(n_64),
.B1(n_65),
.B2(n_161),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_13),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_13),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_67),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_13),
.A2(n_48),
.B1(n_51),
.B2(n_67),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_13),
.A2(n_34),
.B1(n_35),
.B2(n_67),
.Y(n_255)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_16),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_114),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_113),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_99),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_21),
.B(n_99),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_72),
.C(n_80),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_22),
.A2(n_23),
.B1(n_72),
.B2(n_73),
.Y(n_139)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_57),
.B2(n_71),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_41),
.B1(n_55),
.B2(n_56),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_26),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_26),
.B(n_56),
.C(n_57),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_27),
.A2(n_31),
.B1(n_32),
.B2(n_78),
.Y(n_77)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_29),
.A2(n_30),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_29),
.A2(n_30),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

AOI32xp33_ASAP7_75t_L g209 ( 
.A1(n_29),
.A2(n_35),
.A3(n_199),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_31),
.B(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_31),
.A2(n_32),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_34),
.Y(n_35)
);

AOI32xp33_ASAP7_75t_L g148 ( 
.A1(n_34),
.A2(n_45),
.A3(n_51),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

NAND2xp33_ASAP7_75t_SL g211 ( 
.A(n_34),
.B(n_37),
.Y(n_211)
);

O2A1O1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_44),
.B(n_46),
.C(n_47),
.Y(n_43)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_37),
.Y(n_210)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_39),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_41),
.A2(n_56),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_52),
.B(n_53),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_42),
.A2(n_52),
.B1(n_93),
.B2(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_42),
.A2(n_228),
.B(n_229),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_42),
.A2(n_52),
.B1(n_129),
.B2(n_255),
.Y(n_274)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_47),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_43),
.A2(n_47),
.B1(n_75),
.B2(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_43),
.B(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_43),
.A2(n_47),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_48),
.B(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_51),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_52),
.B(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_52),
.A2(n_160),
.B(n_162),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_52),
.B(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_52),
.A2(n_162),
.B(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_71),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_58),
.A2(n_68),
.B1(n_69),
.B2(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_58),
.A2(n_133),
.B(n_136),
.Y(n_132)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_59),
.B(n_97),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_59),
.A2(n_246),
.B(n_247),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_59),
.A2(n_60),
.B1(n_134),
.B2(n_269),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_60),
.B(n_97),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_61),
.A2(n_64),
.B(n_181),
.C(n_242),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_64),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_66),
.A2(n_68),
.B(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_68),
.B(n_181),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_68),
.A2(n_96),
.B(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_73),
.A2(n_74),
.B(n_77),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_79),
.A2(n_108),
.B1(n_110),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_80),
.A2(n_81),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_89),
.B(n_94),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_94),
.B1(n_95),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_82),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_82),
.A2(n_90),
.B1(n_91),
.B2(n_120),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_85),
.B(n_88),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_83),
.A2(n_85),
.B1(n_88),
.B2(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_83),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_83),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_83),
.B(n_168),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_83),
.A2(n_85),
.B1(n_208),
.B2(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_83),
.A2(n_87),
.B1(n_127),
.B2(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_85),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_85),
.A2(n_173),
.B(n_183),
.Y(n_182)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_86),
.B(n_167),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_86),
.A2(n_184),
.B(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_86),
.A2(n_174),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_119),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_112),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_108),
.A2(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_110),
.B(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_110),
.A2(n_218),
.B(n_219),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_110),
.A2(n_131),
.B(n_219),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_140),
.B(n_313),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_137),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_116),
.B(n_137),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_123),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_301)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_123),
.B(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_130),
.C(n_132),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_124),
.A2(n_125),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_126),
.B(n_128),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_130),
.B(n_132),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_136),
.Y(n_247)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI321xp33_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_293),
.A3(n_302),
.B1(n_307),
.B2(n_312),
.C(n_315),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_257),
.C(n_289),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_231),
.B(n_256),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_213),
.B(n_230),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_194),
.B(n_212),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_169),
.B(n_193),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_154),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_147),
.B(n_154),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_151),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_152),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_153),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_164),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_159),
.C(n_164),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_160),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_165),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_178),
.B(n_192),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_171),
.B(n_177),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_185),
.B(n_191),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_180),
.B(n_182),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_189),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_195),
.B(n_196),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_205),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_202),
.C(n_205),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_200),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_204),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_209),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_214),
.B(n_215),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_225),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_226),
.C(n_227),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_221),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_222),
.C(n_223),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_218),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_224),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_232),
.B(n_233),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_244),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_235),
.B(n_236),
.C(n_244),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_240),
.B1(n_241),
.B2(n_243),
.Y(n_236)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_239),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_243),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_248),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_250),
.C(n_253),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_253),
.B2(n_254),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_252),
.Y(n_265)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_258),
.A2(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_276),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_259),
.B(n_276),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_271),
.C(n_275),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_263),
.C(n_270),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_267),
.B2(n_270),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_267),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_275),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_274),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_276)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_277),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_285),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_278),
.B(n_285),
.C(n_288),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_282),
.C(n_283),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_286),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_291),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_300),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_300),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_298),
.C(n_299),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_298),
.Y(n_306)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_303),
.A2(n_308),
.B(n_311),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_304),
.B(n_305),
.Y(n_311)
);


endmodule