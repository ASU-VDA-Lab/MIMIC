module fake_jpeg_12546_n_622 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_622);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_622;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_14),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_29),
.B(n_16),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_66),
.B(n_68),
.Y(n_128)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_67),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_44),
.B(n_14),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_70),
.Y(n_163)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_19),
.B(n_11),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_72),
.B(n_80),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_73),
.Y(n_172)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_75),
.Y(n_179)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_77),
.Y(n_166)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_78),
.Y(n_155)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_79),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_24),
.B(n_13),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_81),
.Y(n_168)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_83),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_84),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_19),
.B(n_11),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_85),
.B(n_88),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx5_ASAP7_75t_SL g138 ( 
.A(n_87),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_28),
.B(n_13),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_90),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_17),
.Y(n_91)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_91),
.Y(n_186)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_17),
.Y(n_95)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_17),
.Y(n_96)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_17),
.Y(n_97)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_28),
.B(n_11),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_102),
.B(n_106),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_103),
.Y(n_177)
);

BUFx8_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_105),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_40),
.B(n_10),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_109),
.Y(n_203)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_41),
.B(n_10),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_111),
.B(n_112),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_41),
.B(n_9),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_26),
.Y(n_115)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_115),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_116),
.Y(n_189)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_117),
.Y(n_205)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_43),
.Y(n_118)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_26),
.Y(n_119)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g120 ( 
.A(n_20),
.Y(n_120)
);

INVx4_ASAP7_75t_SL g183 ( 
.A(n_120),
.Y(n_183)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_121),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_20),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_122),
.B(n_125),
.Y(n_187)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_20),
.Y(n_123)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_43),
.Y(n_124)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_124),
.Y(n_198)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_20),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_120),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_126),
.B(n_156),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_72),
.B(n_42),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_140),
.B(n_200),
.Y(n_220)
);

BUFx4f_ASAP7_75t_SL g143 ( 
.A(n_120),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g227 ( 
.A(n_143),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_80),
.A2(n_36),
.B1(n_56),
.B2(n_48),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_144),
.A2(n_184),
.B1(n_197),
.B2(n_199),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_115),
.A2(n_37),
.B1(n_26),
.B2(n_34),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_150),
.A2(n_34),
.B1(n_83),
.B2(n_90),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_66),
.B(n_43),
.Y(n_152)
);

NAND2x1_ASAP7_75t_L g261 ( 
.A(n_152),
.B(n_59),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_53),
.Y(n_156)
);

INVx6_ASAP7_75t_SL g169 ( 
.A(n_87),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_169),
.Y(n_250)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_85),
.Y(n_171)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_98),
.A2(n_36),
.B1(n_56),
.B2(n_48),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_175),
.A2(n_185),
.B1(n_107),
.B2(n_34),
.Y(n_217)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_102),
.Y(n_176)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_96),
.A2(n_36),
.B1(n_48),
.B2(n_56),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_86),
.A2(n_34),
.B1(n_37),
.B2(n_47),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_112),
.B(n_42),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_194),
.B(n_46),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_60),
.A2(n_37),
.B1(n_38),
.B2(n_55),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_64),
.A2(n_38),
.B1(n_39),
.B2(n_55),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_104),
.B(n_57),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_70),
.Y(n_201)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_122),
.B(n_53),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_202),
.B(n_173),
.Y(n_252)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_73),
.Y(n_204)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_75),
.Y(n_207)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_138),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_208),
.B(n_260),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g283 ( 
.A(n_213),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_152),
.B(n_128),
.C(n_147),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_215),
.B(n_261),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_217),
.A2(n_240),
.B1(n_243),
.B2(n_254),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_218),
.Y(n_299)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_219),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_142),
.A2(n_109),
.B1(n_91),
.B2(n_105),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_222),
.A2(n_232),
.B1(n_258),
.B2(n_264),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_223),
.A2(n_268),
.B1(n_275),
.B2(n_174),
.Y(n_303)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_138),
.Y(n_224)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_224),
.Y(n_310)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_183),
.Y(n_225)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_225),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_142),
.B(n_57),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_226),
.B(n_241),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_135),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_228),
.Y(n_302)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_133),
.Y(n_229)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_229),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_230),
.Y(n_295)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_231),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_156),
.A2(n_84),
.B1(n_103),
.B2(n_100),
.Y(n_232)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_149),
.Y(n_233)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_233),
.Y(n_297)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_159),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_234),
.Y(n_290)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_235),
.Y(n_313)
);

AO22x2_ASAP7_75t_L g236 ( 
.A1(n_150),
.A2(n_59),
.B1(n_97),
.B2(n_95),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_236),
.B(n_243),
.Y(n_292)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_129),
.Y(n_238)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_238),
.Y(n_287)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_146),
.Y(n_239)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_239),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_189),
.A2(n_107),
.B1(n_34),
.B2(n_47),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_161),
.B(n_40),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_167),
.Y(n_242)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_242),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_134),
.A2(n_34),
.B1(n_47),
.B2(n_23),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g244 ( 
.A(n_135),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_244),
.Y(n_329)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_154),
.Y(n_245)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_245),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_161),
.B(n_54),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_246),
.B(n_262),
.Y(n_335)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_160),
.Y(n_247)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_247),
.Y(n_307)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_195),
.Y(n_248)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_248),
.Y(n_333)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_170),
.Y(n_249)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_249),
.Y(n_336)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_165),
.Y(n_251)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_251),
.Y(n_315)
);

NAND3xp33_ASAP7_75t_L g331 ( 
.A(n_252),
.B(n_270),
.C(n_3),
.Y(n_331)
);

BUFx2_ASAP7_75t_SL g253 ( 
.A(n_168),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_253),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_132),
.A2(n_23),
.B1(n_27),
.B2(n_35),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_182),
.Y(n_255)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_255),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_148),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_256),
.Y(n_314)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_180),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_257),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_141),
.A2(n_54),
.B1(n_25),
.B2(n_51),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_136),
.A2(n_27),
.B1(n_35),
.B2(n_50),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_259),
.A2(n_266),
.B1(n_269),
.B2(n_277),
.Y(n_330)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_148),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_194),
.B(n_51),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_202),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_265),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_175),
.A2(n_185),
.B1(n_199),
.B2(n_197),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_158),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_137),
.A2(n_166),
.B1(n_155),
.B2(n_127),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_141),
.B(n_128),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_267),
.B(n_273),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_144),
.A2(n_39),
.B1(n_25),
.B2(n_50),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_157),
.A2(n_46),
.B1(n_9),
.B2(n_2),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_151),
.Y(n_271)
);

INVx8_ASAP7_75t_L g311 ( 
.A(n_271),
.Y(n_311)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_198),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_278),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_130),
.B(n_8),
.C(n_1),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_173),
.B(n_0),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_274),
.B(n_187),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_203),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_275)
);

BUFx6f_ASAP7_75t_SL g276 ( 
.A(n_143),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_276),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_191),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_277)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_131),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_162),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_280),
.Y(n_293)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_186),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_230),
.B(n_139),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_284),
.B(n_312),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_292),
.A2(n_277),
.B1(n_269),
.B2(n_225),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_296),
.B(n_300),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_221),
.B(n_205),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_303),
.A2(n_237),
.B1(n_236),
.B2(n_223),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_276),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_305),
.B(n_323),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_209),
.B(n_205),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_308),
.B(n_309),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_220),
.B(n_153),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_212),
.B(n_164),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_273),
.B(n_145),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_316),
.B(n_318),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_215),
.B(n_190),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_250),
.B(n_196),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_320),
.B(n_322),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_208),
.B(n_181),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_261),
.B(n_151),
.Y(n_323)
);

INVxp33_ASAP7_75t_SL g326 ( 
.A(n_224),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_326),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_216),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_327),
.B(n_3),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_214),
.B(n_206),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_328),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_331),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_217),
.A2(n_206),
.B1(n_192),
.B2(n_179),
.Y(n_334)
);

OR2x6_ASAP7_75t_L g344 ( 
.A(n_334),
.B(n_236),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_240),
.C(n_211),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_338),
.B(n_349),
.C(n_355),
.Y(n_397)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_310),
.Y(n_339)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_339),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_342),
.A2(n_344),
.B1(n_351),
.B2(n_358),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_310),
.Y(n_343)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_343),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_303),
.A2(n_256),
.B1(n_233),
.B2(n_260),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_346),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_295),
.A2(n_254),
.B(n_259),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_347),
.A2(n_376),
.B(n_381),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_288),
.B(n_210),
.C(n_266),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_287),
.Y(n_350)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_306),
.A2(n_236),
.B1(n_280),
.B2(n_278),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_302),
.Y(n_352)
);

INVx8_ASAP7_75t_L g413 ( 
.A(n_352),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_354),
.A2(n_362),
.B1(n_364),
.B2(n_290),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_288),
.B(n_235),
.C(n_228),
.Y(n_355)
);

OAI32xp33_ASAP7_75t_L g357 ( 
.A1(n_309),
.A2(n_282),
.A3(n_284),
.B1(n_316),
.B2(n_296),
.Y(n_357)
);

AOI32xp33_ASAP7_75t_L g390 ( 
.A1(n_357),
.A2(n_294),
.A3(n_335),
.B1(n_301),
.B2(n_315),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_306),
.A2(n_192),
.B1(n_163),
.B2(n_179),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_287),
.Y(n_359)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_359),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_282),
.B(n_271),
.C(n_229),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_360),
.B(n_370),
.C(n_374),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_292),
.A2(n_172),
.B1(n_163),
.B2(n_234),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_361),
.A2(n_371),
.B1(n_281),
.B2(n_319),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_291),
.A2(n_172),
.B1(n_248),
.B2(n_255),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_330),
.A2(n_244),
.B1(n_219),
.B2(n_231),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_366),
.B(n_380),
.Y(n_385)
);

INVx8_ASAP7_75t_L g367 ( 
.A(n_329),
.Y(n_367)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_367),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_285),
.A2(n_218),
.B1(n_213),
.B2(n_244),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_368),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_312),
.B(n_227),
.C(n_4),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_323),
.A2(n_227),
.B1(n_4),
.B2(n_5),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_313),
.Y(n_372)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_372),
.Y(n_418)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_298),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_373),
.B(n_375),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_317),
.A2(n_227),
.B(n_4),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_374),
.A2(n_337),
.B(n_290),
.Y(n_396)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_298),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_317),
.A2(n_3),
.B(n_5),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_290),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_377),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_311),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_378),
.B(n_379),
.Y(n_398)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_301),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_327),
.B(n_6),
.Y(n_380)
);

O2A1O1Ixp33_ASAP7_75t_L g381 ( 
.A1(n_317),
.A2(n_8),
.B(n_314),
.C(n_286),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_386),
.B(n_371),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_356),
.B(n_293),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_388),
.B(n_392),
.Y(n_428)
);

AO21x1_ASAP7_75t_L g440 ( 
.A1(n_390),
.A2(n_353),
.B(n_370),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_365),
.Y(n_392)
);

MAJx2_ASAP7_75t_L g393 ( 
.A(n_365),
.B(n_307),
.C(n_315),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_393),
.B(n_400),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_369),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_395),
.B(n_369),
.Y(n_429)
);

AND2x2_ASAP7_75t_SL g449 ( 
.A(n_396),
.B(n_289),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_338),
.A2(n_307),
.B1(n_333),
.B2(n_325),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_399),
.A2(n_403),
.B1(n_408),
.B2(n_411),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_355),
.B(n_360),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_341),
.B(n_340),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_401),
.B(n_414),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_357),
.B(n_325),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_402),
.B(n_412),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_349),
.A2(n_333),
.B1(n_313),
.B2(n_324),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_366),
.B(n_297),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_405),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_380),
.B(n_297),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_344),
.A2(n_324),
.B1(n_311),
.B2(n_302),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_410),
.A2(n_379),
.B1(n_359),
.B2(n_375),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_344),
.A2(n_302),
.B1(n_319),
.B2(n_281),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_363),
.B(n_336),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_341),
.B(n_336),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_348),
.B(n_321),
.Y(n_415)
);

XNOR2x1_ASAP7_75t_L g425 ( 
.A(n_415),
.B(n_416),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_406),
.A2(n_347),
.B(n_381),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_419),
.A2(n_424),
.B(n_426),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_386),
.A2(n_344),
.B1(n_351),
.B2(n_342),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_421),
.A2(n_430),
.B1(n_450),
.B2(n_384),
.Y(n_463)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_383),
.Y(n_423)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_423),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_411),
.A2(n_361),
.B(n_344),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_382),
.A2(n_344),
.B(n_345),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_392),
.B(n_340),
.Y(n_427)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_427),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_429),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_398),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_431),
.B(n_438),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_388),
.B(n_348),
.Y(n_433)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_433),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_382),
.A2(n_358),
.B(n_364),
.Y(n_434)
);

XOR2x1_ASAP7_75t_SL g484 ( 
.A(n_434),
.B(n_442),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_435),
.A2(n_440),
.B1(n_403),
.B2(n_390),
.Y(n_454)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_387),
.Y(n_436)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_436),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_409),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_437),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_396),
.B(n_376),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_406),
.A2(n_373),
.B(n_350),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_439),
.B(n_412),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_404),
.B(n_339),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_441),
.B(n_443),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_402),
.A2(n_409),
.B(n_408),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_387),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_389),
.A2(n_378),
.B1(n_353),
.B2(n_352),
.Y(n_446)
);

XOR2x1_ASAP7_75t_L g475 ( 
.A(n_446),
.B(n_449),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_384),
.B(n_372),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_447),
.B(n_418),
.Y(n_469)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_407),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_451),
.Y(n_476)
);

OAI22xp33_ASAP7_75t_SL g450 ( 
.A1(n_399),
.A2(n_378),
.B1(n_289),
.B2(n_299),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_405),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_407),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_452),
.B(n_453),
.Y(n_482)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_418),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_454),
.A2(n_420),
.B1(n_449),
.B2(n_437),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_425),
.B(n_400),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_457),
.B(n_468),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_425),
.B(n_397),
.C(n_416),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_458),
.B(n_481),
.C(n_438),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_429),
.A2(n_423),
.B1(n_446),
.B2(n_444),
.Y(n_459)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_459),
.Y(n_506)
);

OA21x2_ASAP7_75t_L g461 ( 
.A1(n_430),
.A2(n_410),
.B(n_391),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_461),
.A2(n_426),
.B(n_434),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_463),
.A2(n_466),
.B1(n_471),
.B2(n_435),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_450),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_464),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_421),
.A2(n_415),
.B1(n_397),
.B2(n_385),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_425),
.B(n_393),
.Y(n_468)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_469),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_470),
.A2(n_481),
.B(n_455),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_430),
.A2(n_385),
.B1(n_417),
.B2(n_413),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_444),
.B(n_332),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_472),
.B(n_480),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_422),
.B(n_417),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_473),
.B(n_445),
.Y(n_496)
);

AOI22x1_ASAP7_75t_L g478 ( 
.A1(n_430),
.A2(n_394),
.B1(n_413),
.B2(n_367),
.Y(n_478)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_478),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_427),
.B(n_332),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_422),
.B(n_394),
.C(n_321),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_431),
.Y(n_483)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_483),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_451),
.B(n_299),
.Y(n_485)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_485),
.Y(n_501)
);

INVx13_ASAP7_75t_L g486 ( 
.A(n_485),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_486),
.Y(n_521)
);

AO22x1_ASAP7_75t_L g488 ( 
.A1(n_479),
.A2(n_437),
.B1(n_439),
.B2(n_419),
.Y(n_488)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_488),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_473),
.B(n_445),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_489),
.B(n_496),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_490),
.A2(n_492),
.B1(n_463),
.B2(n_471),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_461),
.A2(n_420),
.B1(n_449),
.B2(n_432),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_493),
.A2(n_508),
.B(n_484),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_483),
.B(n_428),
.Y(n_495)
);

CKINVDCx14_ASAP7_75t_R g515 ( 
.A(n_495),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_468),
.B(n_428),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_499),
.B(n_511),
.C(n_512),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_457),
.B(n_433),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_SL g522 ( 
.A(n_500),
.B(n_455),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_482),
.B(n_432),
.Y(n_502)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_502),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_462),
.B(n_452),
.Y(n_503)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_503),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_504),
.A2(n_461),
.B1(n_478),
.B2(n_424),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_474),
.B(n_447),
.Y(n_505)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_505),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_507),
.B(n_510),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_479),
.A2(n_442),
.B(n_449),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_482),
.Y(n_509)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_509),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_465),
.B(n_448),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_458),
.B(n_440),
.C(n_438),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_466),
.B(n_440),
.C(n_438),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_514),
.B(n_484),
.C(n_475),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_502),
.B(n_456),
.Y(n_518)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_518),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_522),
.B(n_489),
.Y(n_550)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_523),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_SL g547 ( 
.A1(n_525),
.A2(n_488),
.B(n_529),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_526),
.B(n_514),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_509),
.B(n_460),
.Y(n_527)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_527),
.Y(n_548)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_513),
.Y(n_528)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_528),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_506),
.A2(n_467),
.B1(n_476),
.B2(n_475),
.Y(n_530)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_530),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_511),
.B(n_476),
.C(n_467),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_532),
.B(n_533),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_486),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_500),
.B(n_478),
.C(n_460),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_535),
.B(n_537),
.C(n_507),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_536),
.A2(n_490),
.B1(n_492),
.B2(n_498),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_512),
.B(n_441),
.C(n_477),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_501),
.B(n_477),
.Y(n_538)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_538),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_501),
.B(n_436),
.Y(n_539)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_539),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_540),
.B(n_544),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_521),
.B(n_494),
.Y(n_541)
);

AOI21x1_ASAP7_75t_SL g562 ( 
.A1(n_541),
.A2(n_545),
.B(n_547),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_521),
.B(n_494),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_549),
.A2(n_523),
.B1(n_543),
.B2(n_553),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_550),
.B(n_508),
.Y(n_576)
);

CKINVDCx16_ASAP7_75t_R g552 ( 
.A(n_518),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_552),
.B(n_557),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_524),
.B(n_491),
.C(n_496),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_554),
.B(n_556),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_524),
.B(n_491),
.C(n_499),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_515),
.B(n_532),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_519),
.B(n_527),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_559),
.B(n_539),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_560),
.A2(n_565),
.B1(n_558),
.B2(n_542),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_546),
.B(n_520),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_563),
.B(n_566),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_543),
.A2(n_487),
.B1(n_516),
.B2(n_531),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_553),
.A2(n_487),
.B1(n_498),
.B2(n_536),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_SL g567 ( 
.A1(n_544),
.A2(n_529),
.B(n_525),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_567),
.A2(n_573),
.B(n_574),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_568),
.B(n_548),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_556),
.B(n_537),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_569),
.B(n_570),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_554),
.B(n_540),
.C(n_534),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_550),
.B(n_534),
.C(n_535),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_571),
.B(n_572),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_547),
.B(n_522),
.C(n_526),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_549),
.B(n_530),
.C(n_555),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_555),
.B(n_538),
.C(n_517),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_SL g590 ( 
.A(n_576),
.B(n_453),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g577 ( 
.A1(n_562),
.A2(n_541),
.B(n_545),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_577),
.B(n_581),
.Y(n_599)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_579),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_564),
.B(n_559),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_564),
.B(n_558),
.C(n_548),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_582),
.B(n_528),
.C(n_513),
.Y(n_600)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_584),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_569),
.B(n_542),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_586),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_574),
.B(n_488),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_587),
.B(n_589),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_L g588 ( 
.A1(n_562),
.A2(n_493),
.B(n_551),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_588),
.B(n_572),
.C(n_576),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_573),
.B(n_551),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_590),
.B(n_568),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_SL g591 ( 
.A1(n_585),
.A2(n_570),
.B(n_561),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_591),
.A2(n_582),
.B(n_586),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_595),
.B(n_596),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_578),
.B(n_575),
.C(n_571),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_597),
.B(n_600),
.Y(n_604)
);

BUFx24_ASAP7_75t_SL g602 ( 
.A(n_599),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_602),
.B(n_603),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_600),
.B(n_583),
.C(n_580),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_605),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_598),
.B(n_589),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_SL g612 ( 
.A1(n_606),
.A2(n_607),
.B1(n_497),
.B2(n_590),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_598),
.B(n_584),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_SL g608 ( 
.A1(n_601),
.A2(n_592),
.B1(n_594),
.B2(n_604),
.Y(n_608)
);

XOR2xp5_ASAP7_75t_L g615 ( 
.A(n_608),
.B(n_283),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_604),
.B(n_593),
.C(n_587),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_610),
.B(n_612),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_611),
.B(n_443),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_614),
.B(n_615),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_613),
.B(n_609),
.C(n_329),
.Y(n_617)
);

BUFx24_ASAP7_75t_SL g618 ( 
.A(n_617),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_618),
.A2(n_609),
.B(n_616),
.Y(n_619)
);

A2O1A1Ixp33_ASAP7_75t_L g620 ( 
.A1(n_619),
.A2(n_283),
.B(n_304),
.C(n_305),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_620),
.B(n_283),
.Y(n_621)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_621),
.B(n_283),
.Y(n_622)
);


endmodule