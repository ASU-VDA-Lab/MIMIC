module fake_netlist_1_738_n_668 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_668);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_668;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_476;
wire n_227;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_535;
wire n_225;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_494;
wire n_223;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_59), .Y(n_78) );
BUFx5_ASAP7_75t_L g79 ( .A(n_39), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_28), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_62), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_19), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_13), .Y(n_83) );
INVxp67_ASAP7_75t_L g84 ( .A(n_3), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_29), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_42), .Y(n_86) );
HB1xp67_ASAP7_75t_L g87 ( .A(n_21), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_74), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_26), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_72), .Y(n_90) );
HB1xp67_ASAP7_75t_L g91 ( .A(n_75), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_60), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_32), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_54), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_20), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_16), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_13), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_19), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_17), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_16), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_67), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_69), .Y(n_102) );
BUFx2_ASAP7_75t_L g103 ( .A(n_27), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_24), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_49), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_31), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_47), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_51), .Y(n_108) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_20), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_70), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_22), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_7), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_35), .Y(n_113) );
BUFx5_ASAP7_75t_L g114 ( .A(n_34), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_38), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_73), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_37), .Y(n_117) );
INVxp33_ASAP7_75t_L g118 ( .A(n_7), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_18), .Y(n_119) );
INVxp33_ASAP7_75t_SL g120 ( .A(n_17), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_56), .Y(n_121) );
INVxp67_ASAP7_75t_SL g122 ( .A(n_45), .Y(n_122) );
CKINVDCx16_ASAP7_75t_R g123 ( .A(n_36), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_18), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_26), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_88), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_123), .Y(n_127) );
BUFx3_ASAP7_75t_L g128 ( .A(n_103), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_88), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_90), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_117), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_90), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_82), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_79), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_102), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_79), .Y(n_136) );
BUFx3_ASAP7_75t_L g137 ( .A(n_103), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_117), .Y(n_138) );
NAND2xp33_ASAP7_75t_R g139 ( .A(n_93), .B(n_0), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_93), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_118), .B(n_0), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_102), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_116), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_78), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_116), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_120), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_95), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_120), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_80), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_91), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_95), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_81), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_89), .B(n_1), .Y(n_153) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_118), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_79), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_79), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_87), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_84), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_79), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_85), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_121), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_86), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_94), .B(n_1), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_121), .Y(n_164) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_89), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_83), .B(n_2), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_121), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_128), .B(n_101), .Y(n_168) );
BUFx2_ASAP7_75t_L g169 ( .A(n_154), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_153), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_154), .B(n_96), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_128), .B(n_108), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_128), .B(n_125), .Y(n_173) );
INVxp67_ASAP7_75t_SL g174 ( .A(n_137), .Y(n_174) );
OAI22xp5_ASAP7_75t_L g175 ( .A1(n_146), .A2(n_124), .B1(n_97), .B2(n_98), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_161), .Y(n_176) );
NOR3xp33_ASAP7_75t_L g177 ( .A(n_148), .B(n_100), .C(n_119), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_137), .B(n_105), .Y(n_179) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_161), .Y(n_180) );
NAND2x1p5_ASAP7_75t_L g181 ( .A(n_153), .B(n_110), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_137), .B(n_99), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_141), .A2(n_111), .B1(n_104), .B2(n_112), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_144), .B(n_106), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_161), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_153), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_161), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_153), .B(n_109), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_161), .Y(n_189) );
BUFx2_ASAP7_75t_L g190 ( .A(n_140), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_144), .B(n_113), .Y(n_191) );
INVx4_ASAP7_75t_L g192 ( .A(n_166), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_134), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_165), .B(n_109), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_149), .B(n_107), .Y(n_195) );
CKINVDCx11_ASAP7_75t_R g196 ( .A(n_147), .Y(n_196) );
INVx2_ASAP7_75t_SL g197 ( .A(n_165), .Y(n_197) );
OR2x2_ASAP7_75t_L g198 ( .A(n_141), .B(n_109), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_161), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_134), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_164), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_136), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_136), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_131), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_149), .B(n_115), .Y(n_205) );
INVx5_ASAP7_75t_L g206 ( .A(n_164), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_136), .Y(n_207) );
INVxp67_ASAP7_75t_L g208 ( .A(n_143), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_166), .B(n_109), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_155), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_166), .B(n_109), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_139), .A2(n_92), .B1(n_122), .B2(n_114), .Y(n_212) );
AND2x4_ASAP7_75t_SL g213 ( .A(n_166), .B(n_121), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_155), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_150), .B(n_121), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_164), .Y(n_216) );
BUFx3_ASAP7_75t_L g217 ( .A(n_155), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_156), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_126), .A2(n_114), .B(n_79), .C(n_4), .Y(n_219) );
NAND3xp33_ASAP7_75t_L g220 ( .A(n_160), .B(n_114), .C(n_79), .Y(n_220) );
OR2x6_ASAP7_75t_L g221 ( .A(n_163), .B(n_2), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_126), .B(n_3), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_156), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_164), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_164), .Y(n_225) );
BUFx2_ASAP7_75t_L g226 ( .A(n_145), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_156), .Y(n_227) );
NAND2x1p5_ASAP7_75t_L g228 ( .A(n_129), .B(n_114), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_228), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_197), .B(n_162), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_196), .Y(n_231) );
CKINVDCx8_ASAP7_75t_R g232 ( .A(n_204), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_217), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_197), .B(n_152), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_174), .B(n_142), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_172), .B(n_142), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_188), .Y(n_237) );
NOR2xp33_ASAP7_75t_R g238 ( .A(n_190), .B(n_133), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_169), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_222), .Y(n_240) );
INVx2_ASAP7_75t_SL g241 ( .A(n_170), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_169), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_179), .B(n_130), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_171), .B(n_127), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_222), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_190), .Y(n_246) );
BUFx2_ASAP7_75t_L g247 ( .A(n_221), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_177), .A2(n_158), .B1(n_139), .B2(n_163), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_168), .B(n_129), .Y(n_249) );
AO22x1_ASAP7_75t_L g250 ( .A1(n_226), .A2(n_138), .B1(n_151), .B2(n_157), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_228), .Y(n_251) );
OR2x2_ASAP7_75t_L g252 ( .A(n_226), .B(n_152), .Y(n_252) );
BUFx3_ASAP7_75t_L g253 ( .A(n_217), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_181), .A2(n_135), .B1(n_132), .B2(n_130), .Y(n_254) );
BUFx2_ASAP7_75t_L g255 ( .A(n_208), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_222), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_194), .B(n_135), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_222), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_221), .Y(n_259) );
NOR2x1_ASAP7_75t_L g260 ( .A(n_198), .B(n_132), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_217), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_194), .Y(n_262) );
OR2x2_ASAP7_75t_L g263 ( .A(n_171), .B(n_4), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_198), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_186), .B(n_159), .Y(n_265) );
AOI21xp33_ASAP7_75t_L g266 ( .A1(n_212), .A2(n_159), .B(n_6), .Y(n_266) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_221), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_173), .B(n_159), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_173), .B(n_114), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_221), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_181), .A2(n_167), .B1(n_164), .B2(n_8), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_228), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_209), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_209), .Y(n_274) );
INVxp67_ASAP7_75t_SL g275 ( .A(n_170), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_182), .B(n_114), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_218), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_221), .Y(n_278) );
OR2x6_ASAP7_75t_L g279 ( .A(n_181), .B(n_167), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_182), .B(n_114), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_170), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_209), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_188), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_218), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_212), .A2(n_167), .B1(n_6), .B2(n_8), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_175), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_192), .B(n_5), .Y(n_287) );
OR2x2_ASAP7_75t_L g288 ( .A(n_183), .B(n_5), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_186), .A2(n_167), .B1(n_10), .B2(n_11), .Y(n_289) );
INVx5_ASAP7_75t_L g290 ( .A(n_188), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_192), .B(n_167), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_183), .B(n_9), .Y(n_292) );
BUFx4f_ASAP7_75t_L g293 ( .A(n_209), .Y(n_293) );
INVx4_ASAP7_75t_L g294 ( .A(n_279), .Y(n_294) );
NOR2xp67_ASAP7_75t_SL g295 ( .A(n_229), .B(n_186), .Y(n_295) );
BUFx4f_ASAP7_75t_L g296 ( .A(n_287), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_237), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_237), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_237), .Y(n_299) );
A2O1A1Ixp33_ASAP7_75t_L g300 ( .A1(n_240), .A2(n_219), .B(n_211), .C(n_188), .Y(n_300) );
AOI21xp33_ASAP7_75t_SL g301 ( .A1(n_231), .A2(n_215), .B(n_191), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_265), .A2(n_186), .B(n_192), .Y(n_302) );
NOR2xp33_ASAP7_75t_SL g303 ( .A(n_232), .B(n_239), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_265), .A2(n_192), .B(n_213), .Y(n_304) );
AND2x4_ASAP7_75t_L g305 ( .A(n_234), .B(n_211), .Y(n_305) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_229), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_234), .B(n_211), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_283), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_229), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_283), .Y(n_310) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_229), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_283), .Y(n_312) );
INVx5_ASAP7_75t_L g313 ( .A(n_279), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_273), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_281), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_247), .A2(n_213), .B1(n_211), .B2(n_184), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_281), .Y(n_317) );
INVx2_ASAP7_75t_SL g318 ( .A(n_287), .Y(n_318) );
INVxp67_ASAP7_75t_L g319 ( .A(n_242), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g320 ( .A1(n_247), .A2(n_213), .B1(n_205), .B2(n_195), .Y(n_320) );
OAI21xp5_ASAP7_75t_L g321 ( .A1(n_233), .A2(n_261), .B(n_260), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g322 ( .A1(n_239), .A2(n_220), .B1(n_218), .B2(n_193), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_238), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_242), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_291), .A2(n_202), .B(n_178), .Y(n_325) );
INVx2_ASAP7_75t_SL g326 ( .A(n_287), .Y(n_326) );
INVxp67_ASAP7_75t_L g327 ( .A(n_246), .Y(n_327) );
INVx3_ASAP7_75t_SL g328 ( .A(n_231), .Y(n_328) );
INVx1_ASAP7_75t_SL g329 ( .A(n_252), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_234), .B(n_207), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_233), .Y(n_331) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_229), .B(n_202), .Y(n_332) );
BUFx3_ASAP7_75t_L g333 ( .A(n_253), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_274), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_282), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_245), .Y(n_336) );
O2A1O1Ixp5_ASAP7_75t_SL g337 ( .A1(n_266), .A2(n_218), .B(n_203), .C(n_210), .Y(n_337) );
INVx2_ASAP7_75t_SL g338 ( .A(n_279), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_281), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_244), .B(n_207), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_261), .Y(n_341) );
BUFx2_ASAP7_75t_L g342 ( .A(n_279), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_277), .Y(n_343) );
OA21x2_ASAP7_75t_L g344 ( .A1(n_300), .A2(n_269), .B(n_276), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_336), .Y(n_345) );
OR2x6_ASAP7_75t_L g346 ( .A(n_318), .B(n_259), .Y(n_346) );
A2O1A1Ixp33_ASAP7_75t_L g347 ( .A1(n_340), .A2(n_296), .B(n_258), .C(n_256), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_336), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_328), .Y(n_349) );
BUFx3_ASAP7_75t_L g350 ( .A(n_306), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_324), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_329), .B(n_286), .Y(n_352) );
INVxp33_ASAP7_75t_L g353 ( .A(n_303), .Y(n_353) );
OAI22xp33_ASAP7_75t_L g354 ( .A1(n_296), .A2(n_288), .B1(n_252), .B2(n_286), .Y(n_354) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_296), .A2(n_254), .B(n_249), .Y(n_355) );
OAI221xp5_ASAP7_75t_L g356 ( .A1(n_319), .A2(n_288), .B1(n_248), .B2(n_263), .C(n_230), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_330), .Y(n_357) );
INVx2_ASAP7_75t_SL g358 ( .A(n_313), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_305), .A2(n_292), .B1(n_270), .B2(n_267), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_314), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_318), .A2(n_280), .B(n_236), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_313), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_314), .Y(n_363) );
OAI21xp5_ASAP7_75t_L g364 ( .A1(n_337), .A2(n_293), .B(n_285), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_327), .B(n_255), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_313), .B(n_251), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_305), .A2(n_292), .B1(n_278), .B2(n_293), .Y(n_367) );
BUFx12f_ASAP7_75t_L g368 ( .A(n_323), .Y(n_368) );
INVx2_ASAP7_75t_SL g369 ( .A(n_313), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_313), .B(n_251), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_305), .B(n_263), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_307), .A2(n_293), .B1(n_264), .B2(n_262), .Y(n_372) );
AOI21x1_ASAP7_75t_L g373 ( .A1(n_295), .A2(n_176), .B(n_185), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_306), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_294), .B(n_251), .Y(n_375) );
INVxp33_ASAP7_75t_L g376 ( .A(n_365), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_345), .B(n_334), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_349), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_366), .Y(n_379) );
INVx3_ASAP7_75t_L g380 ( .A(n_366), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_361), .A2(n_326), .B(n_320), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_357), .B(n_326), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_357), .B(n_307), .Y(n_383) );
BUFx2_ASAP7_75t_L g384 ( .A(n_366), .Y(n_384) );
AOI22xp33_ASAP7_75t_SL g385 ( .A1(n_356), .A2(n_323), .B1(n_342), .B2(n_294), .Y(n_385) );
OAI221xp5_ASAP7_75t_L g386 ( .A1(n_356), .A2(n_301), .B1(n_243), .B2(n_289), .C(n_316), .Y(n_386) );
AOI222xp33_ASAP7_75t_L g387 ( .A1(n_354), .A2(n_250), .B1(n_335), .B2(n_328), .C1(n_334), .C2(n_257), .Y(n_387) );
NAND3xp33_ASAP7_75t_L g388 ( .A(n_364), .B(n_337), .C(n_321), .Y(n_388) );
NAND3xp33_ASAP7_75t_SL g389 ( .A(n_355), .B(n_342), .C(n_232), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_345), .Y(n_390) );
AO21x2_ASAP7_75t_L g391 ( .A1(n_364), .A2(n_271), .B(n_332), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_368), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_368), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_371), .A2(n_307), .B1(n_294), .B2(n_338), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_352), .B(n_298), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_371), .A2(n_268), .B1(n_338), .B2(n_297), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_348), .A2(n_268), .B1(n_308), .B2(n_297), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_348), .B(n_268), .Y(n_398) );
BUFx3_ASAP7_75t_L g399 ( .A(n_366), .Y(n_399) );
AOI222xp33_ASAP7_75t_L g400 ( .A1(n_360), .A2(n_235), .B1(n_308), .B2(n_299), .C1(n_310), .C2(n_312), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_359), .A2(n_309), .B1(n_306), .B2(n_311), .Y(n_401) );
OAI21xp5_ASAP7_75t_SL g402 ( .A1(n_353), .A2(n_322), .B(n_251), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_360), .A2(n_333), .B1(n_343), .B2(n_341), .Y(n_403) );
AO21x2_ASAP7_75t_L g404 ( .A1(n_388), .A2(n_347), .B(n_361), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_390), .Y(n_405) );
INVxp67_ASAP7_75t_SL g406 ( .A(n_398), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_390), .B(n_363), .Y(n_407) );
OAI211xp5_ASAP7_75t_L g408 ( .A1(n_387), .A2(n_351), .B(n_372), .C(n_367), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_390), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_387), .A2(n_355), .B1(n_362), .B2(n_363), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_398), .B(n_362), .Y(n_411) );
BUFx2_ASAP7_75t_L g412 ( .A(n_384), .Y(n_412) );
OAI22xp33_ASAP7_75t_L g413 ( .A1(n_376), .A2(n_346), .B1(n_358), .B2(n_369), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_376), .A2(n_395), .B1(n_386), .B2(n_385), .C(n_383), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_398), .B(n_375), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_377), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_378), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_385), .A2(n_368), .B1(n_346), .B2(n_375), .Y(n_418) );
NAND4xp75_ASAP7_75t_L g419 ( .A(n_395), .B(n_369), .C(n_358), .D(n_370), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_383), .B(n_375), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_383), .B(n_375), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_384), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_396), .A2(n_346), .B1(n_309), .B2(n_311), .Y(n_423) );
AOI222xp33_ASAP7_75t_L g424 ( .A1(n_386), .A2(n_290), .B1(n_295), .B2(n_343), .C1(n_275), .C2(n_341), .Y(n_424) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_396), .A2(n_344), .B1(n_346), .B2(n_304), .C(n_290), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g426 ( .A1(n_394), .A2(n_346), .B1(n_272), .B2(n_251), .Y(n_426) );
NAND4xp25_ASAP7_75t_L g427 ( .A(n_400), .B(n_302), .C(n_325), .D(n_11), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_382), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g429 ( .A(n_400), .B(n_306), .Y(n_429) );
OAI21x1_ASAP7_75t_SL g430 ( .A1(n_401), .A2(n_344), .B(n_373), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_380), .B(n_350), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_384), .B(n_344), .Y(n_432) );
NAND2xp33_ASAP7_75t_SL g433 ( .A(n_401), .B(n_306), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_389), .A2(n_344), .B1(n_333), .B2(n_281), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_379), .B(n_350), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_382), .B(n_290), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_379), .B(n_350), .Y(n_437) );
INVx3_ASAP7_75t_L g438 ( .A(n_405), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_409), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_432), .Y(n_440) );
INVx6_ASAP7_75t_L g441 ( .A(n_431), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_414), .A2(n_389), .B1(n_394), .B2(n_388), .C(n_402), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_433), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_432), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_412), .B(n_379), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_433), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_407), .Y(n_447) );
BUFx2_ASAP7_75t_L g448 ( .A(n_412), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_407), .Y(n_449) );
AOI22xp33_ASAP7_75t_SL g450 ( .A1(n_408), .A2(n_399), .B1(n_380), .B2(n_378), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_430), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_416), .B(n_380), .Y(n_452) );
OAI33xp33_ASAP7_75t_L g453 ( .A1(n_427), .A2(n_392), .A3(n_393), .B1(n_12), .B2(n_14), .B3(n_15), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_428), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_430), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_415), .B(n_380), .Y(n_456) );
NAND2xp33_ASAP7_75t_R g457 ( .A(n_417), .B(n_9), .Y(n_457) );
AOI33xp33_ASAP7_75t_L g458 ( .A1(n_410), .A2(n_397), .A3(n_382), .B1(n_403), .B2(n_15), .B3(n_21), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_415), .B(n_399), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_428), .B(n_402), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_406), .B(n_399), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_422), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_404), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_404), .Y(n_464) );
OR2x2_ASAP7_75t_SL g465 ( .A(n_435), .B(n_309), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_411), .B(n_397), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_404), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_429), .Y(n_468) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_420), .A2(n_381), .B1(n_403), .B2(n_290), .C(n_391), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_421), .B(n_381), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_431), .B(n_391), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_431), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_435), .B(n_391), .Y(n_473) );
INVx4_ASAP7_75t_L g474 ( .A(n_437), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_418), .B(n_436), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_426), .A2(n_391), .B1(n_331), .B2(n_272), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_423), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_437), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_434), .B(n_391), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_417), .B(n_374), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_419), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_419), .Y(n_482) );
NAND2x1p5_ASAP7_75t_L g483 ( .A(n_413), .B(n_374), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_424), .B(n_374), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_425), .B(n_374), .Y(n_485) );
NAND2x1p5_ASAP7_75t_L g486 ( .A(n_438), .B(n_309), .Y(n_486) );
AOI221xp5_ASAP7_75t_L g487 ( .A1(n_453), .A2(n_167), .B1(n_290), .B2(n_178), .C(n_214), .Y(n_487) );
INVxp33_ASAP7_75t_L g488 ( .A(n_478), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_438), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_449), .B(n_10), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_472), .B(n_50), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_438), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_443), .A2(n_309), .B(n_311), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_473), .B(n_12), .Y(n_494) );
OAI33xp33_ASAP7_75t_L g495 ( .A1(n_480), .A2(n_14), .A3(n_22), .B1(n_23), .B2(n_24), .B3(n_25), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_438), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_449), .B(n_23), .Y(n_497) );
NOR3xp33_ASAP7_75t_L g498 ( .A(n_450), .B(n_339), .C(n_317), .Y(n_498) );
INVx2_ASAP7_75t_SL g499 ( .A(n_441), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_462), .B(n_25), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_473), .B(n_311), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_447), .B(n_311), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_471), .B(n_30), .Y(n_503) );
NOR4xp25_ASAP7_75t_SL g504 ( .A(n_457), .B(n_33), .C(n_40), .D(n_41), .Y(n_504) );
INVxp67_ASAP7_75t_L g505 ( .A(n_448), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_439), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_471), .B(n_43), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_443), .A2(n_272), .B(n_339), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_454), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_440), .B(n_44), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_454), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_452), .Y(n_512) );
NAND2xp33_ASAP7_75t_SL g513 ( .A(n_474), .B(n_272), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_448), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_465), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_465), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_460), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_440), .B(n_46), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_466), .B(n_315), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_459), .B(n_315), .Y(n_520) );
NOR2x1_ASAP7_75t_L g521 ( .A(n_474), .B(n_317), .Y(n_521) );
BUFx3_ASAP7_75t_L g522 ( .A(n_441), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_459), .B(n_315), .Y(n_523) );
OAI222xp33_ASAP7_75t_L g524 ( .A1(n_474), .A2(n_373), .B1(n_331), .B2(n_241), .C1(n_277), .C2(n_284), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_440), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_445), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_445), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_444), .B(n_48), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_456), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_444), .B(n_52), .Y(n_530) );
NAND2xp33_ASAP7_75t_SL g531 ( .A(n_474), .B(n_272), .Y(n_531) );
INVx3_ASAP7_75t_L g532 ( .A(n_451), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_444), .B(n_53), .Y(n_533) );
INVx2_ASAP7_75t_SL g534 ( .A(n_441), .Y(n_534) );
INVx4_ASAP7_75t_L g535 ( .A(n_483), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_470), .B(n_55), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_456), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_479), .B(n_57), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_461), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_529), .B(n_472), .Y(n_540) );
O2A1O1Ixp33_ASAP7_75t_L g541 ( .A1(n_500), .A2(n_481), .B(n_475), .C(n_482), .Y(n_541) );
AOI221xp5_ASAP7_75t_L g542 ( .A1(n_495), .A2(n_442), .B1(n_463), .B2(n_464), .C(n_467), .Y(n_542) );
NOR2xp67_ASAP7_75t_SL g543 ( .A(n_497), .B(n_482), .Y(n_543) );
OAI322xp33_ASAP7_75t_L g544 ( .A1(n_517), .A2(n_468), .A3(n_481), .B1(n_464), .B2(n_463), .C1(n_467), .C2(n_477), .Y(n_544) );
OAI21xp33_ASAP7_75t_SL g545 ( .A1(n_535), .A2(n_468), .B(n_458), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_506), .Y(n_546) );
INVx2_ASAP7_75t_SL g547 ( .A(n_521), .Y(n_547) );
OAI22xp33_ASAP7_75t_L g548 ( .A1(n_535), .A2(n_482), .B1(n_446), .B2(n_483), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_509), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_511), .Y(n_550) );
OAI32xp33_ASAP7_75t_L g551 ( .A1(n_488), .A2(n_483), .A3(n_455), .B1(n_451), .B2(n_477), .Y(n_551) );
OAI332xp33_ASAP7_75t_L g552 ( .A1(n_497), .A2(n_485), .A3(n_455), .B1(n_451), .B2(n_469), .B3(n_446), .C1(n_479), .C2(n_476), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_537), .B(n_461), .Y(n_553) );
INVx1_ASAP7_75t_SL g554 ( .A(n_513), .Y(n_554) );
OAI22xp33_ASAP7_75t_SL g555 ( .A1(n_535), .A2(n_441), .B1(n_476), .B2(n_455), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_526), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_527), .B(n_484), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_513), .A2(n_441), .B1(n_484), .B2(n_281), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_539), .B(n_58), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_514), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_488), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_525), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_494), .B(n_61), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_512), .B(n_63), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_494), .B(n_64), .Y(n_565) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_505), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_515), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_501), .B(n_65), .Y(n_568) );
INVxp67_ASAP7_75t_L g569 ( .A(n_516), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_531), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_525), .B(n_66), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_528), .A2(n_241), .B1(n_284), .B2(n_253), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_490), .Y(n_573) );
INVx2_ASAP7_75t_SL g574 ( .A(n_522), .Y(n_574) );
NAND2x1_ASAP7_75t_SL g575 ( .A(n_538), .B(n_185), .Y(n_575) );
OAI21xp33_ASAP7_75t_L g576 ( .A1(n_538), .A2(n_189), .B(n_225), .Y(n_576) );
OAI321xp33_ASAP7_75t_L g577 ( .A1(n_487), .A2(n_68), .A3(n_71), .B1(n_76), .B2(n_77), .C(n_180), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_501), .B(n_176), .Y(n_578) );
NAND4xp75_ASAP7_75t_L g579 ( .A(n_499), .B(n_201), .C(n_185), .D(n_187), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_489), .B(n_224), .Y(n_580) );
OAI332xp33_ASAP7_75t_L g581 ( .A1(n_519), .A2(n_224), .A3(n_187), .B1(n_189), .B2(n_216), .B3(n_199), .C1(n_225), .C2(n_201), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_531), .A2(n_203), .B(n_223), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_498), .A2(n_201), .B1(n_187), .B2(n_189), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_534), .B(n_214), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_503), .A2(n_225), .B1(n_216), .B2(n_199), .Y(n_585) );
NAND2xp33_ASAP7_75t_L g586 ( .A(n_534), .B(n_210), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_524), .A2(n_193), .B(n_200), .Y(n_587) );
NAND2xp33_ASAP7_75t_L g588 ( .A(n_554), .B(n_503), .Y(n_588) );
XNOR2xp5_ASAP7_75t_L g589 ( .A(n_553), .B(n_507), .Y(n_589) );
OAI21xp33_ASAP7_75t_SL g590 ( .A1(n_554), .A2(n_507), .B(n_533), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_566), .B(n_522), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g592 ( .A(n_574), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_567), .B(n_532), .Y(n_593) );
NOR2xp33_ASAP7_75t_R g594 ( .A(n_586), .B(n_533), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_573), .B(n_536), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_561), .B(n_496), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_546), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_549), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_540), .B(n_496), .Y(n_599) );
INVxp67_ASAP7_75t_L g600 ( .A(n_543), .Y(n_600) );
XOR2x2_ASAP7_75t_L g601 ( .A(n_575), .B(n_520), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_550), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_560), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_541), .B(n_536), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_556), .Y(n_605) );
XOR2xp5_ASAP7_75t_L g606 ( .A(n_557), .B(n_523), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_570), .A2(n_528), .B1(n_492), .B2(n_489), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_542), .B(n_532), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_569), .B(n_532), .Y(n_609) );
OAI22xp5_ASAP7_75t_SL g610 ( .A1(n_570), .A2(n_486), .B1(n_491), .B2(n_502), .Y(n_610) );
INVxp67_ASAP7_75t_L g611 ( .A(n_547), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_562), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_584), .B(n_486), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_578), .B(n_486), .Y(n_614) );
XOR2x2_ASAP7_75t_L g615 ( .A(n_563), .B(n_491), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_580), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_580), .Y(n_617) );
AOI22xp33_ASAP7_75t_SL g618 ( .A1(n_555), .A2(n_491), .B1(n_530), .B2(n_518), .Y(n_618) );
NOR4xp25_ASAP7_75t_SL g619 ( .A(n_576), .B(n_504), .C(n_518), .D(n_510), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_544), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_552), .B(n_530), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_620), .B(n_552), .Y(n_622) );
OAI22xp33_ASAP7_75t_L g623 ( .A1(n_621), .A2(n_600), .B1(n_592), .B2(n_558), .Y(n_623) );
NOR2xp67_ASAP7_75t_SL g624 ( .A(n_613), .B(n_564), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_591), .Y(n_625) );
INVx1_ASAP7_75t_SL g626 ( .A(n_615), .Y(n_626) );
OAI21x1_ASAP7_75t_L g627 ( .A1(n_608), .A2(n_493), .B(n_508), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_590), .B(n_548), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_596), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_621), .A2(n_545), .B1(n_565), .B2(n_568), .Y(n_630) );
INVx1_ASAP7_75t_SL g631 ( .A(n_614), .Y(n_631) );
AOI321xp33_ASAP7_75t_L g632 ( .A1(n_604), .A2(n_551), .A3(n_581), .B1(n_572), .B2(n_559), .C(n_577), .Y(n_632) );
NOR2x1_ASAP7_75t_L g633 ( .A(n_588), .B(n_572), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_618), .A2(n_585), .B1(n_583), .B2(n_571), .Y(n_634) );
XOR2xp5_ASAP7_75t_L g635 ( .A(n_589), .B(n_579), .Y(n_635) );
OAI211xp5_ASAP7_75t_L g636 ( .A1(n_618), .A2(n_582), .B(n_587), .C(n_199), .Y(n_636) );
AOI322xp5_ASAP7_75t_L g637 ( .A1(n_595), .A2(n_611), .A3(n_600), .B1(n_605), .B2(n_603), .C1(n_602), .C2(n_598), .Y(n_637) );
AOI321xp33_ASAP7_75t_L g638 ( .A1(n_607), .A2(n_224), .A3(n_200), .B1(n_223), .B2(n_227), .C(n_180), .Y(n_638) );
A2O1A1Ixp33_ASAP7_75t_L g639 ( .A1(n_611), .A2(n_206), .B(n_227), .C(n_180), .Y(n_639) );
NOR2xp67_ASAP7_75t_L g640 ( .A(n_628), .B(n_607), .Y(n_640) );
AOI21xp33_ASAP7_75t_L g641 ( .A1(n_622), .A2(n_617), .B(n_616), .Y(n_641) );
INVx1_ASAP7_75t_SL g642 ( .A(n_625), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_630), .A2(n_610), .B1(n_606), .B2(n_593), .Y(n_643) );
INVx3_ASAP7_75t_SL g644 ( .A(n_631), .Y(n_644) );
NOR2xp33_ASAP7_75t_R g645 ( .A(n_630), .B(n_597), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_623), .A2(n_594), .B1(n_601), .B2(n_593), .Y(n_646) );
OAI211xp5_ASAP7_75t_L g647 ( .A1(n_628), .A2(n_619), .B(n_609), .C(n_612), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_637), .B(n_599), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_629), .B(n_180), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_633), .A2(n_180), .B1(n_206), .B2(n_626), .Y(n_650) );
NAND2x1p5_ASAP7_75t_L g651 ( .A(n_624), .B(n_206), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_636), .A2(n_180), .B1(n_206), .B2(n_635), .Y(n_652) );
A2O1A1Ixp33_ASAP7_75t_L g653 ( .A1(n_632), .A2(n_206), .B(n_638), .C(n_639), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_639), .A2(n_622), .B(n_623), .C(n_628), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_634), .A2(n_630), .B1(n_628), .B2(n_592), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_627), .Y(n_656) );
CKINVDCx5p33_ASAP7_75t_R g657 ( .A(n_644), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_642), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_642), .Y(n_659) );
NOR3xp33_ASAP7_75t_L g660 ( .A(n_647), .B(n_655), .C(n_654), .Y(n_660) );
A2O1A1Ixp33_ASAP7_75t_L g661 ( .A1(n_660), .A2(n_640), .B(n_643), .C(n_650), .Y(n_661) );
OAI221xp5_ASAP7_75t_L g662 ( .A1(n_659), .A2(n_646), .B1(n_648), .B2(n_653), .C(n_641), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_657), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_663), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_661), .Y(n_665) );
OA22x2_ASAP7_75t_L g666 ( .A1(n_665), .A2(n_658), .B1(n_662), .B2(n_656), .Y(n_666) );
AOI22xp33_ASAP7_75t_SL g667 ( .A1(n_666), .A2(n_664), .B1(n_645), .B2(n_651), .Y(n_667) );
AOI21xp5_ASAP7_75t_L g668 ( .A1(n_667), .A2(n_649), .B(n_652), .Y(n_668) );
endmodule