module fake_jpeg_23397_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_33),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_34),
.B(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_31),
.Y(n_49)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_40),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_43),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx5_ASAP7_75t_SL g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_32),
.B1(n_21),
.B2(n_20),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_47),
.A2(n_32),
.B1(n_16),
.B2(n_30),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_66),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_21),
.B1(n_20),
.B2(n_29),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_56),
.B1(n_25),
.B2(n_30),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_32),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_28),
.Y(n_70)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_59),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_21),
.B1(n_20),
.B2(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_64),
.Y(n_94)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_44),
.C(n_41),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_70),
.Y(n_103)
);

NAND3xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_22),
.C(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_73),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_69),
.A2(n_86),
.B(n_88),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_43),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_78),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_42),
.B1(n_24),
.B2(n_19),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_72),
.A2(n_76),
.B1(n_1),
.B2(n_2),
.Y(n_106)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

OR2x4_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_18),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_91),
.B(n_17),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_42),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_62),
.A2(n_24),
.B1(n_16),
.B2(n_22),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_81),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_29),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_84),
.Y(n_115)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_27),
.C(n_18),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_28),
.B1(n_19),
.B2(n_3),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_50),
.B(n_17),
.Y(n_89)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_60),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_28),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_65),
.B(n_17),
.Y(n_93)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_101),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_70),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_100),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_110),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_106),
.B(n_116),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_107),
.Y(n_129)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_112),
.Y(n_137)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_76),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_119),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_67),
.B1(n_77),
.B2(n_85),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_78),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_71),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_124),
.Y(n_152)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_122),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_82),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_109),
.B(n_75),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_136),
.B(n_114),
.Y(n_138)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_126),
.Y(n_142)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_128),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_91),
.Y(n_130)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_131),
.A2(n_134),
.B(n_135),
.Y(n_139)
);

AOI22x1_ASAP7_75t_SL g134 ( 
.A1(n_97),
.A2(n_72),
.B1(n_86),
.B2(n_1),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_4),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_138),
.B(n_131),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_99),
.C(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_153),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_98),
.B(n_104),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_148),
.B(n_151),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_123),
.A2(n_100),
.B1(n_113),
.B2(n_96),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_137),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_136),
.C(n_152),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_7),
.B(n_8),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_9),
.C(n_12),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_13),
.C(n_124),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_133),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_166),
.Y(n_173)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_162),
.Y(n_170)
);

BUFx12f_ASAP7_75t_SL g176 ( 
.A(n_157),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_158),
.B(n_161),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_146),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_126),
.Y(n_164)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_144),
.B(n_120),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_167),
.C(n_154),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_160),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_168),
.A2(n_169),
.B(n_135),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_159),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_167),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_175),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_157),
.B(n_145),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_171),
.Y(n_184)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_165),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_183),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_176),
.A2(n_143),
.B1(n_150),
.B2(n_139),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_181),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_143),
.B1(n_150),
.B2(n_153),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_170),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_184),
.A2(n_168),
.B(n_173),
.Y(n_189)
);

NOR2xp67_ASAP7_75t_SL g188 ( 
.A(n_185),
.B(n_150),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_172),
.B(n_169),
.Y(n_186)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_189),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_178),
.C(n_179),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_191),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_127),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_194),
.B(n_193),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_SL g198 ( 
.A1(n_192),
.A2(n_180),
.B(n_129),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_199),
.A2(n_196),
.B(n_127),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_200),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_128),
.Y(n_203)
);


endmodule