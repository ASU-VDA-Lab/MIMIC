module fake_netlist_1_813_n_701 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_701, n_699);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_701;
output n_699;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_25), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_5), .Y(n_79) );
INVxp33_ASAP7_75t_L g80 ( .A(n_41), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_48), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_43), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_28), .Y(n_83) );
BUFx2_ASAP7_75t_L g84 ( .A(n_37), .Y(n_84) );
CKINVDCx14_ASAP7_75t_R g85 ( .A(n_16), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_58), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_3), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_47), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_22), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_31), .Y(n_90) );
INVxp33_ASAP7_75t_SL g91 ( .A(n_44), .Y(n_91) );
CKINVDCx16_ASAP7_75t_R g92 ( .A(n_40), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_69), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_14), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_24), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_8), .Y(n_96) );
INVxp67_ASAP7_75t_L g97 ( .A(n_26), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_63), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_29), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_71), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_3), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_59), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_70), .Y(n_103) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_30), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_74), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_19), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_53), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_2), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_76), .Y(n_109) );
INVx3_ASAP7_75t_L g110 ( .A(n_38), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_49), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_56), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_13), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_42), .Y(n_114) );
OR2x2_ASAP7_75t_L g115 ( .A(n_75), .B(n_36), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_77), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_12), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_6), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_17), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_65), .Y(n_120) );
NOR2xp67_ASAP7_75t_L g121 ( .A(n_34), .B(n_27), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_73), .Y(n_122) );
INVxp67_ASAP7_75t_SL g123 ( .A(n_9), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_7), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_72), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_78), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_83), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_92), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_86), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_110), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_94), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_88), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_110), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_84), .B(n_0), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_80), .B(n_0), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_119), .B(n_1), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_89), .Y(n_137) );
NAND2xp33_ASAP7_75t_L g138 ( .A(n_109), .B(n_68), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_93), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_85), .Y(n_140) );
AND2x4_ASAP7_75t_SL g141 ( .A(n_82), .B(n_32), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_87), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_104), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_110), .Y(n_144) );
BUFx2_ASAP7_75t_L g145 ( .A(n_108), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_96), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_98), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_100), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_104), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_102), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_101), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_113), .B(n_1), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_105), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_106), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_118), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_124), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_104), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_112), .Y(n_158) );
NOR2xp33_ASAP7_75t_SL g159 ( .A(n_81), .B(n_33), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_108), .B(n_2), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_82), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_120), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_91), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_163) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_125), .A2(n_39), .B(n_66), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_104), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_115), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_111), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_97), .Y(n_168) );
NAND2x1p5_ASAP7_75t_L g169 ( .A(n_145), .B(n_121), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_130), .Y(n_170) );
INVx8_ASAP7_75t_L g171 ( .A(n_166), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_152), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g173 ( .A1(n_152), .A2(n_135), .B1(n_166), .B2(n_132), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_145), .B(n_114), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_128), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_166), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_152), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g178 ( .A1(n_135), .A2(n_91), .B1(n_123), .B2(n_117), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_143), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_168), .B(n_122), .Y(n_180) );
AND2x2_ASAP7_75t_SL g181 ( .A(n_141), .B(n_111), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_143), .Y(n_182) );
INVx4_ASAP7_75t_L g183 ( .A(n_166), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_130), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_143), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_168), .B(n_122), .Y(n_186) );
INVx6_ASAP7_75t_L g187 ( .A(n_166), .Y(n_187) );
INVx4_ASAP7_75t_SL g188 ( .A(n_143), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_161), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_133), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_158), .B(n_114), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_126), .B(n_127), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_143), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_126), .B(n_107), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_133), .Y(n_195) );
INVx5_ASAP7_75t_L g196 ( .A(n_151), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_128), .B(n_107), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_127), .B(n_99), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_149), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_129), .B(n_99), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_149), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_149), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_129), .B(n_90), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_132), .B(n_90), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_149), .Y(n_205) );
AND2x2_ASAP7_75t_SL g206 ( .A(n_141), .B(n_116), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_144), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_149), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_144), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_157), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_157), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_151), .B(n_81), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_151), .B(n_79), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_137), .B(n_103), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_157), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_137), .B(n_116), .Y(n_216) );
INVx4_ASAP7_75t_SL g217 ( .A(n_157), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_139), .B(n_147), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_139), .B(n_94), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_142), .Y(n_220) );
BUFx3_ASAP7_75t_L g221 ( .A(n_157), .Y(n_221) );
INVx4_ASAP7_75t_SL g222 ( .A(n_165), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_165), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_165), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_140), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_165), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_165), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_150), .Y(n_228) );
OR2x6_ASAP7_75t_L g229 ( .A(n_136), .B(n_4), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_147), .B(n_95), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_136), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_176), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_198), .B(n_148), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_180), .B(n_140), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_183), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_183), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_183), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_228), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_228), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_174), .B(n_155), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_178), .A2(n_160), .B1(n_134), .B2(n_138), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_176), .Y(n_242) );
INVx4_ASAP7_75t_L g243 ( .A(n_171), .Y(n_243) );
OR2x6_ASAP7_75t_L g244 ( .A(n_229), .B(n_156), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_187), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_198), .B(n_148), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_187), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_203), .B(n_154), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_218), .A2(n_146), .B(n_154), .C(n_150), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_187), .Y(n_250) );
INVx2_ASAP7_75t_SL g251 ( .A(n_212), .Y(n_251) );
NAND2x1p5_ASAP7_75t_L g252 ( .A(n_212), .B(n_163), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_203), .B(n_162), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_212), .B(n_159), .Y(n_254) );
INVx4_ASAP7_75t_L g255 ( .A(n_171), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_213), .B(n_162), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_171), .Y(n_257) );
AND3x2_ASAP7_75t_SL g258 ( .A(n_181), .B(n_167), .C(n_161), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_171), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_190), .Y(n_260) );
INVxp67_ASAP7_75t_L g261 ( .A(n_216), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_204), .B(n_153), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_213), .B(n_153), .Y(n_263) );
INVx2_ASAP7_75t_SL g264 ( .A(n_213), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_204), .B(n_172), .Y(n_265) );
BUFx12f_ASAP7_75t_L g266 ( .A(n_229), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_190), .Y(n_267) );
INVx5_ASAP7_75t_L g268 ( .A(n_170), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_229), .Y(n_269) );
INVx4_ASAP7_75t_L g270 ( .A(n_196), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_186), .B(n_197), .Y(n_271) );
AO22x1_ASAP7_75t_L g272 ( .A1(n_175), .A2(n_167), .B1(n_131), .B2(n_164), .Y(n_272) );
INVxp33_ASAP7_75t_L g273 ( .A(n_216), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_177), .B(n_164), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_200), .B(n_10), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_220), .B(n_164), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_195), .Y(n_277) );
INVxp67_ASAP7_75t_SL g278 ( .A(n_216), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_186), .B(n_164), .Y(n_279) );
INVx2_ASAP7_75t_SL g280 ( .A(n_196), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_196), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_173), .B(n_46), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_207), .Y(n_283) );
OAI22x1_ASAP7_75t_L g284 ( .A1(n_219), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_192), .A2(n_11), .B1(n_13), .B2(n_14), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_194), .B(n_15), .Y(n_286) );
BUFx8_ASAP7_75t_L g287 ( .A(n_219), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_191), .B(n_52), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_200), .B(n_51), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_189), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_230), .B(n_54), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_192), .B(n_50), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_196), .Y(n_293) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_169), .B(n_55), .Y(n_294) );
BUFx3_ASAP7_75t_L g295 ( .A(n_170), .Y(n_295) );
INVx2_ASAP7_75t_SL g296 ( .A(n_169), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_214), .B(n_15), .Y(n_297) );
NOR2x1_ASAP7_75t_L g298 ( .A(n_214), .B(n_18), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_244), .A2(n_219), .B1(n_181), .B2(n_206), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_244), .B(n_206), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_244), .A2(n_175), .B1(n_231), .B2(n_225), .Y(n_301) );
BUFx2_ASAP7_75t_L g302 ( .A(n_287), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_287), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_274), .A2(n_209), .B(n_184), .Y(n_304) );
OAI21xp33_ASAP7_75t_L g305 ( .A1(n_273), .A2(n_225), .B(n_170), .Y(n_305) );
INVxp67_ASAP7_75t_L g306 ( .A(n_269), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_243), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_275), .A2(n_184), .B1(n_221), .B2(n_224), .Y(n_308) );
O2A1O1Ixp33_ASAP7_75t_L g309 ( .A1(n_261), .A2(n_184), .B(n_221), .C(n_224), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_243), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_255), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_255), .B(n_188), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_266), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_271), .B(n_188), .Y(n_314) );
AO21x2_ASAP7_75t_L g315 ( .A1(n_279), .A2(n_208), .B(n_226), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_278), .A2(n_205), .B1(n_226), .B2(n_223), .Y(n_316) );
BUFx3_ASAP7_75t_L g317 ( .A(n_257), .Y(n_317) );
INVx5_ASAP7_75t_L g318 ( .A(n_281), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_275), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_296), .B(n_20), .Y(n_320) );
AO21x2_ASAP7_75t_L g321 ( .A1(n_279), .A2(n_205), .B(n_223), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_240), .B(n_21), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_290), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_274), .A2(n_182), .B(n_215), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_259), .Y(n_325) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_251), .B(n_188), .Y(n_326) );
INVxp67_ASAP7_75t_L g327 ( .A(n_297), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_238), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_276), .A2(n_215), .B(n_208), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_277), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_233), .B(n_23), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_283), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_281), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_281), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_233), .B(n_217), .Y(n_335) );
INVx3_ASAP7_75t_SL g336 ( .A(n_297), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_270), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_264), .A2(n_202), .B1(n_199), .B2(n_193), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_246), .B(n_35), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_276), .A2(n_202), .B(n_199), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_256), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_270), .Y(n_342) );
INVx2_ASAP7_75t_SL g343 ( .A(n_268), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_260), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_252), .A2(n_263), .B1(n_265), .B2(n_284), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_252), .A2(n_182), .B1(n_193), .B2(n_179), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_239), .Y(n_347) );
OR2x6_ASAP7_75t_L g348 ( .A(n_254), .B(n_227), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_267), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_328), .Y(n_350) );
OAI21x1_ASAP7_75t_L g351 ( .A1(n_329), .A2(n_298), .B(n_291), .Y(n_351) );
OAI21xp5_ASAP7_75t_L g352 ( .A1(n_304), .A2(n_265), .B(n_246), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_315), .Y(n_353) );
NAND3xp33_ASAP7_75t_L g354 ( .A(n_345), .B(n_272), .C(n_249), .Y(n_354) );
OR2x6_ASAP7_75t_L g355 ( .A(n_319), .B(n_294), .Y(n_355) );
OA21x2_ASAP7_75t_L g356 ( .A1(n_340), .A2(n_292), .B(n_288), .Y(n_356) );
INVx4_ASAP7_75t_L g357 ( .A(n_318), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_299), .A2(n_319), .B1(n_300), .B2(n_327), .Y(n_358) );
INVx2_ASAP7_75t_SL g359 ( .A(n_310), .Y(n_359) );
NOR2xp67_ASAP7_75t_SL g360 ( .A(n_334), .B(n_248), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_330), .B(n_248), .Y(n_361) );
OA21x2_ASAP7_75t_L g362 ( .A1(n_324), .A2(n_292), .B(n_286), .Y(n_362) );
AO21x2_ASAP7_75t_L g363 ( .A1(n_315), .A2(n_282), .B(n_262), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_328), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_347), .Y(n_365) );
OA21x2_ASAP7_75t_L g366 ( .A1(n_331), .A2(n_339), .B(n_322), .Y(n_366) );
O2A1O1Ixp33_ASAP7_75t_SL g367 ( .A1(n_314), .A2(n_289), .B(n_253), .C(n_262), .Y(n_367) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_334), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_323), .Y(n_369) );
OAI21x1_ASAP7_75t_L g370 ( .A1(n_346), .A2(n_253), .B(n_242), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_331), .A2(n_232), .B(n_285), .Y(n_371) );
OAI21x1_ASAP7_75t_L g372 ( .A1(n_339), .A2(n_293), .B(n_245), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_334), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_335), .A2(n_247), .B(n_250), .Y(n_374) );
OAI21xp5_ASAP7_75t_L g375 ( .A1(n_347), .A2(n_241), .B(n_235), .Y(n_375) );
A2O1A1Ixp33_ASAP7_75t_L g376 ( .A1(n_322), .A2(n_234), .B(n_237), .C(n_236), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_323), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_332), .Y(n_378) );
CKINVDCx11_ASAP7_75t_R g379 ( .A(n_313), .Y(n_379) );
OR2x6_ASAP7_75t_L g380 ( .A(n_310), .B(n_280), .Y(n_380) );
OAI21x1_ASAP7_75t_L g381 ( .A1(n_309), .A2(n_179), .B(n_268), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_361), .A2(n_301), .B1(n_300), .B2(n_303), .C(n_302), .Y(n_382) );
OAI221xp5_ASAP7_75t_L g383 ( .A1(n_358), .A2(n_336), .B1(n_305), .B2(n_302), .C(n_306), .Y(n_383) );
O2A1O1Ixp33_ASAP7_75t_L g384 ( .A1(n_376), .A2(n_336), .B(n_341), .C(n_348), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_361), .A2(n_308), .B1(n_258), .B2(n_316), .C(n_313), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_350), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_378), .B(n_317), .Y(n_387) );
OAI211xp5_ASAP7_75t_SL g388 ( .A1(n_378), .A2(n_258), .B(n_344), .C(n_338), .Y(n_388) );
AOI22xp33_ASAP7_75t_SL g389 ( .A1(n_366), .A2(n_311), .B1(n_307), .B2(n_320), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_377), .B(n_343), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_366), .A2(n_348), .B1(n_349), .B2(n_343), .Y(n_391) );
NAND2x1p5_ASAP7_75t_L g392 ( .A(n_357), .B(n_318), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_350), .B(n_268), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_364), .B(n_325), .Y(n_394) );
AOI22xp33_ASAP7_75t_SL g395 ( .A1(n_366), .A2(n_307), .B1(n_311), .B2(n_325), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_364), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_365), .Y(n_397) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_366), .A2(n_315), .B(n_321), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_365), .B(n_268), .Y(n_399) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_380), .A2(n_348), .B1(n_317), .B2(n_318), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_352), .A2(n_348), .B1(n_321), .B2(n_349), .Y(n_401) );
CKINVDCx11_ASAP7_75t_R g402 ( .A(n_379), .Y(n_402) );
OR2x6_ASAP7_75t_L g403 ( .A(n_380), .B(n_311), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_354), .A2(n_295), .B1(n_344), .B2(n_307), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_359), .B(n_318), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_380), .A2(n_318), .B1(n_344), .B2(n_337), .Y(n_406) );
INVx4_ASAP7_75t_L g407 ( .A(n_357), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_359), .A2(n_342), .B1(n_337), .B2(n_333), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_375), .A2(n_342), .B1(n_337), .B2(n_321), .C(n_326), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_386), .Y(n_410) );
INVx2_ASAP7_75t_SL g411 ( .A(n_392), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_396), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_397), .B(n_353), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_382), .B(n_354), .Y(n_414) );
OR2x6_ASAP7_75t_L g415 ( .A(n_403), .B(n_380), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_391), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_394), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_387), .B(n_353), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_398), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_403), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_395), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_403), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_407), .Y(n_423) );
INVx3_ASAP7_75t_L g424 ( .A(n_392), .Y(n_424) );
INVx3_ASAP7_75t_L g425 ( .A(n_407), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_393), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_400), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_399), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_405), .B(n_357), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_395), .Y(n_430) );
OAI33xp33_ASAP7_75t_L g431 ( .A1(n_388), .A2(n_353), .A3(n_312), .B1(n_355), .B2(n_369), .B3(n_367), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_401), .B(n_357), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_408), .Y(n_433) );
INVx3_ASAP7_75t_SL g434 ( .A(n_390), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_401), .B(n_380), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_385), .B(n_355), .Y(n_436) );
BUFx2_ASAP7_75t_L g437 ( .A(n_400), .Y(n_437) );
BUFx2_ASAP7_75t_L g438 ( .A(n_409), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_406), .B(n_355), .Y(n_439) );
AO21x2_ASAP7_75t_L g440 ( .A1(n_384), .A2(n_370), .B(n_372), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_383), .Y(n_441) );
AOI211xp5_ASAP7_75t_L g442 ( .A1(n_388), .A2(n_360), .B(n_342), .C(n_337), .Y(n_442) );
INVx3_ASAP7_75t_L g443 ( .A(n_389), .Y(n_443) );
AND2x4_ASAP7_75t_L g444 ( .A(n_404), .B(n_373), .Y(n_444) );
INVx5_ASAP7_75t_L g445 ( .A(n_415), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_413), .B(n_389), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_413), .B(n_363), .Y(n_447) );
NOR2x1_ASAP7_75t_SL g448 ( .A(n_415), .B(n_355), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_410), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_432), .B(n_372), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_410), .Y(n_451) );
AO21x2_ASAP7_75t_L g452 ( .A1(n_419), .A2(n_370), .B(n_374), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_410), .B(n_363), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_412), .Y(n_454) );
AO21x2_ASAP7_75t_L g455 ( .A1(n_419), .A2(n_374), .B(n_363), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_412), .B(n_373), .Y(n_456) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_414), .A2(n_371), .B(n_355), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_412), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_427), .A2(n_360), .B1(n_362), .B2(n_402), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_418), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_418), .Y(n_461) );
AOI21xp5_ASAP7_75t_SL g462 ( .A1(n_415), .A2(n_368), .B(n_362), .Y(n_462) );
AOI22xp33_ASAP7_75t_SL g463 ( .A1(n_427), .A2(n_373), .B1(n_368), .B2(n_337), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_434), .B(n_373), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_417), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_434), .B(n_342), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_417), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_435), .B(n_368), .Y(n_468) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_431), .A2(n_342), .B1(n_333), .B2(n_227), .C(n_201), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_435), .B(n_368), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_417), .Y(n_471) );
NOR2xp67_ASAP7_75t_L g472 ( .A(n_425), .B(n_368), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_426), .B(n_362), .Y(n_473) );
AOI221xp5_ASAP7_75t_L g474 ( .A1(n_421), .A2(n_333), .B1(n_227), .B2(n_211), .C(n_210), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_426), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_432), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_420), .B(n_351), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_442), .A2(n_362), .B(n_356), .Y(n_478) );
INVxp67_ASAP7_75t_L g479 ( .A(n_423), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_426), .B(n_371), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_428), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_425), .Y(n_482) );
NAND3xp33_ASAP7_75t_L g483 ( .A(n_441), .B(n_210), .C(n_185), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_416), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_437), .B(n_356), .Y(n_485) );
AND2x4_ASAP7_75t_L g486 ( .A(n_420), .B(n_351), .Y(n_486) );
OAI33xp33_ASAP7_75t_L g487 ( .A1(n_436), .A2(n_45), .A3(n_57), .B1(n_60), .B2(n_61), .B3(n_62), .Y(n_487) );
BUFx2_ASAP7_75t_L g488 ( .A(n_415), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_416), .Y(n_489) );
NOR2xp33_ASAP7_75t_SL g490 ( .A(n_434), .B(n_334), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_416), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_421), .Y(n_492) );
OAI221xp5_ASAP7_75t_L g493 ( .A1(n_441), .A2(n_356), .B1(n_334), .B2(n_185), .C(n_201), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_430), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_461), .B(n_460), .Y(n_495) );
AND4x1_ASAP7_75t_L g496 ( .A(n_490), .B(n_439), .C(n_430), .D(n_415), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_460), .B(n_428), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_492), .B(n_428), .Y(n_498) );
INVx1_ASAP7_75t_SL g499 ( .A(n_466), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_449), .Y(n_500) );
INVx1_ASAP7_75t_SL g501 ( .A(n_464), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_492), .B(n_441), .Y(n_502) );
INVx3_ASAP7_75t_L g503 ( .A(n_482), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_467), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_467), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_476), .B(n_443), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_479), .A2(n_423), .B(n_425), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_449), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_476), .B(n_443), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_446), .B(n_468), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_465), .Y(n_511) );
NAND2x1p5_ASAP7_75t_L g512 ( .A(n_445), .B(n_425), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_471), .B(n_437), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_472), .B(n_423), .Y(n_514) );
AND2x4_ASAP7_75t_L g515 ( .A(n_445), .B(n_443), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_475), .B(n_481), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_494), .B(n_420), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_494), .B(n_422), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_482), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_475), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_468), .B(n_429), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_488), .A2(n_443), .B1(n_438), .B2(n_439), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_481), .B(n_458), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_458), .B(n_422), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_470), .B(n_446), .Y(n_525) );
NAND4xp25_ASAP7_75t_L g526 ( .A(n_459), .B(n_438), .C(n_422), .D(n_429), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_470), .B(n_429), .Y(n_527) );
INVx2_ASAP7_75t_SL g528 ( .A(n_482), .Y(n_528) );
NOR2x1p5_ASAP7_75t_L g529 ( .A(n_485), .B(n_424), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_447), .B(n_473), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_447), .B(n_440), .Y(n_531) );
OR2x6_ASAP7_75t_L g532 ( .A(n_462), .B(n_411), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_472), .B(n_411), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_473), .B(n_440), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_451), .B(n_429), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_480), .B(n_440), .Y(n_536) );
NOR3xp33_ASAP7_75t_L g537 ( .A(n_487), .B(n_424), .C(n_433), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_451), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_456), .B(n_424), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_454), .B(n_424), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_454), .B(n_444), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_456), .B(n_444), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_480), .B(n_444), .Y(n_543) );
NAND2x1p5_ASAP7_75t_L g544 ( .A(n_445), .B(n_444), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_453), .B(n_433), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_488), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_453), .B(n_433), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_445), .B(n_440), .Y(n_548) );
OAI21xp33_ASAP7_75t_L g549 ( .A1(n_462), .A2(n_211), .B(n_227), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_485), .B(n_381), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_445), .B(n_356), .Y(n_551) );
BUFx3_ASAP7_75t_L g552 ( .A(n_445), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_450), .B(n_381), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_510), .B(n_450), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_495), .Y(n_555) );
INVxp67_ASAP7_75t_L g556 ( .A(n_532), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_510), .B(n_450), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_530), .B(n_450), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_530), .B(n_491), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_525), .B(n_491), .Y(n_560) );
AND2x4_ASAP7_75t_L g561 ( .A(n_515), .B(n_486), .Y(n_561) );
INVx2_ASAP7_75t_SL g562 ( .A(n_512), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_501), .B(n_489), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_504), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_497), .B(n_489), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_505), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_506), .B(n_486), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_511), .B(n_484), .Y(n_568) );
AOI22x1_ASAP7_75t_L g569 ( .A1(n_512), .A2(n_478), .B1(n_457), .B2(n_448), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_521), .B(n_448), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_513), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_499), .B(n_484), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_517), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_506), .B(n_486), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_498), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_527), .B(n_486), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_509), .B(n_477), .Y(n_577) );
INVxp67_ASAP7_75t_SL g578 ( .A(n_514), .Y(n_578) );
NOR3xp33_ASAP7_75t_L g579 ( .A(n_526), .B(n_469), .C(n_483), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_500), .Y(n_580) );
NAND2x1p5_ASAP7_75t_L g581 ( .A(n_533), .B(n_477), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_537), .A2(n_463), .B(n_493), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_500), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_508), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_509), .B(n_477), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_523), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_518), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_531), .B(n_477), .Y(n_588) );
NAND2x1_ASAP7_75t_L g589 ( .A(n_532), .B(n_452), .Y(n_589) );
NAND2x1_ASAP7_75t_SL g590 ( .A(n_515), .B(n_474), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_531), .B(n_455), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_542), .B(n_539), .Y(n_592) );
NAND3xp33_ASAP7_75t_L g593 ( .A(n_537), .B(n_211), .C(n_210), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_518), .B(n_455), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_532), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_524), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_516), .Y(n_597) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_508), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_520), .Y(n_599) );
NOR2xp67_ASAP7_75t_SL g600 ( .A(n_552), .B(n_64), .Y(n_600) );
OAI31xp33_ASAP7_75t_L g601 ( .A1(n_529), .A2(n_455), .A3(n_452), .B(n_67), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_535), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_538), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_546), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_522), .A2(n_452), .B1(n_201), .B2(n_210), .Y(n_605) );
NAND3xp33_ASAP7_75t_SL g606 ( .A(n_601), .B(n_496), .C(n_549), .Y(n_606) );
OAI322xp33_ASAP7_75t_L g607 ( .A1(n_587), .A2(n_543), .A3(n_502), .B1(n_550), .B2(n_541), .C1(n_545), .C2(n_547), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_580), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_579), .A2(n_522), .B1(n_515), .B2(n_553), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_588), .B(n_534), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_598), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_598), .Y(n_612) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_559), .Y(n_613) );
OAI21xp5_ASAP7_75t_L g614 ( .A1(n_593), .A2(n_507), .B(n_514), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_555), .B(n_533), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_564), .Y(n_616) );
AOI221x1_ASAP7_75t_L g617 ( .A1(n_579), .A2(n_503), .B1(n_548), .B2(n_540), .C(n_551), .Y(n_617) );
INVxp67_ASAP7_75t_L g618 ( .A(n_571), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_582), .A2(n_528), .B(n_548), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_566), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_568), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_562), .A2(n_544), .B1(n_552), .B2(n_528), .Y(n_622) );
OAI21xp33_ASAP7_75t_L g623 ( .A1(n_594), .A2(n_534), .B(n_536), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_580), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_588), .B(n_536), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_583), .Y(n_626) );
INVx3_ASAP7_75t_SL g627 ( .A(n_562), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_583), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_586), .Y(n_629) );
INVxp67_ASAP7_75t_SL g630 ( .A(n_578), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_558), .B(n_553), .Y(n_631) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_597), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_584), .Y(n_633) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_596), .Y(n_634) );
INVxp67_ASAP7_75t_SL g635 ( .A(n_578), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_602), .B(n_519), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_573), .B(n_548), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g638 ( .A1(n_556), .A2(n_544), .B1(n_503), .B2(n_211), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_584), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_575), .B(n_503), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_591), .B(n_560), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_599), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_613), .B(n_591), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_634), .Y(n_644) );
OR2x2_ASAP7_75t_L g645 ( .A(n_641), .B(n_554), .Y(n_645) );
AND2x2_ASAP7_75t_SL g646 ( .A(n_609), .B(n_570), .Y(n_646) );
A2O1A1Ixp33_ASAP7_75t_L g647 ( .A1(n_619), .A2(n_556), .B(n_590), .C(n_595), .Y(n_647) );
INVx1_ASAP7_75t_SL g648 ( .A(n_627), .Y(n_648) );
NAND2xp33_ASAP7_75t_L g649 ( .A(n_627), .B(n_595), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_606), .A2(n_589), .B(n_569), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_615), .A2(n_558), .B1(n_557), .B2(n_576), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_632), .B(n_604), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_616), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_616), .Y(n_654) );
XNOR2xp5_ASAP7_75t_L g655 ( .A(n_629), .B(n_592), .Y(n_655) );
INVxp67_ASAP7_75t_L g656 ( .A(n_630), .Y(n_656) );
BUFx2_ASAP7_75t_L g657 ( .A(n_635), .Y(n_657) );
O2A1O1Ixp33_ASAP7_75t_L g658 ( .A1(n_614), .A2(n_581), .B(n_563), .C(n_603), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_610), .B(n_567), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_642), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_621), .B(n_567), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g662 ( .A1(n_617), .A2(n_605), .B(n_600), .Y(n_662) );
NOR2xp33_ASAP7_75t_SL g663 ( .A(n_622), .B(n_581), .Y(n_663) );
A2O1A1Ixp33_ASAP7_75t_L g664 ( .A1(n_623), .A2(n_561), .B(n_577), .C(n_574), .Y(n_664) );
INVxp67_ASAP7_75t_L g665 ( .A(n_611), .Y(n_665) );
OAI211xp5_ASAP7_75t_L g666 ( .A1(n_650), .A2(n_617), .B(n_618), .C(n_637), .Y(n_666) );
OAI211xp5_ASAP7_75t_L g667 ( .A1(n_647), .A2(n_636), .B(n_640), .C(n_621), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_663), .B(n_638), .Y(n_668) );
INVx1_ASAP7_75t_SL g669 ( .A(n_648), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_657), .Y(n_670) );
NAND4xp25_ASAP7_75t_L g671 ( .A(n_662), .B(n_561), .C(n_620), .D(n_585), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_660), .Y(n_672) );
OAI21xp5_ASAP7_75t_L g673 ( .A1(n_656), .A2(n_611), .B(n_612), .Y(n_673) );
NAND2xp33_ASAP7_75t_R g674 ( .A(n_649), .B(n_612), .Y(n_674) );
INVx1_ASAP7_75t_SL g675 ( .A(n_644), .Y(n_675) );
OAI22xp33_ASAP7_75t_L g676 ( .A1(n_656), .A2(n_642), .B1(n_631), .B2(n_610), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_653), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_646), .B(n_658), .Y(n_678) );
INVx2_ASAP7_75t_SL g679 ( .A(n_655), .Y(n_679) );
O2A1O1Ixp33_ASAP7_75t_L g680 ( .A1(n_678), .A2(n_658), .B(n_664), .C(n_665), .Y(n_680) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_670), .Y(n_681) );
OAI221xp5_ASAP7_75t_SL g682 ( .A1(n_666), .A2(n_651), .B1(n_643), .B2(n_652), .C(n_661), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_671), .A2(n_665), .B1(n_654), .B2(n_659), .Y(n_683) );
NOR3xp33_ASAP7_75t_L g684 ( .A(n_668), .B(n_607), .C(n_639), .Y(n_684) );
OAI221xp5_ASAP7_75t_L g685 ( .A1(n_667), .A2(n_645), .B1(n_639), .B2(n_633), .C(n_628), .Y(n_685) );
NOR3xp33_ASAP7_75t_L g686 ( .A(n_667), .B(n_633), .C(n_628), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_679), .A2(n_625), .B1(n_631), .B2(n_626), .C(n_624), .Y(n_687) );
INVx5_ASAP7_75t_L g688 ( .A(n_681), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_684), .B(n_675), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_683), .Y(n_690) );
NOR4xp25_ASAP7_75t_L g691 ( .A(n_682), .B(n_669), .C(n_673), .D(n_676), .Y(n_691) );
NOR3xp33_ASAP7_75t_L g692 ( .A(n_689), .B(n_680), .C(n_685), .Y(n_692) );
NAND5xp2_ASAP7_75t_L g693 ( .A(n_690), .B(n_687), .C(n_686), .D(n_674), .E(n_673), .Y(n_693) );
OA22x2_ASAP7_75t_L g694 ( .A1(n_691), .A2(n_677), .B1(n_672), .B2(n_625), .Y(n_694) );
NAND4xp25_ASAP7_75t_L g695 ( .A(n_692), .B(n_688), .C(n_561), .D(n_572), .Y(n_695) );
OAI222xp33_ASAP7_75t_L g696 ( .A1(n_694), .A2(n_688), .B1(n_626), .B2(n_624), .C1(n_608), .C2(n_565), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_695), .A2(n_693), .B1(n_608), .B2(n_201), .Y(n_697) );
OAI21xp5_ASAP7_75t_L g698 ( .A1(n_697), .A2(n_696), .B(n_217), .Y(n_698) );
UNKNOWN g699 ( );
OAI22xp33_ASAP7_75t_L g700 ( .A1(n_699), .A2(n_185), .B1(n_217), .B2(n_222), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_700), .A2(n_185), .B1(n_222), .B2(n_692), .Y(n_701) );
endmodule