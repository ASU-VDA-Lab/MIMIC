module fake_jpeg_2748_n_121 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_32),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_11),
.B(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_6),
.B(n_24),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_52),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_0),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_34),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_42),
.Y(n_63)
);

NAND3xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_73),
.C(n_75),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_62),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_36),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_74),
.Y(n_79)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_37),
.Y(n_73)
);

AOI32xp33_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_45),
.A3(n_44),
.B1(n_40),
.B2(n_38),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_49),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_64),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_78),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_57),
.B(n_1),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_50),
.B1(n_48),
.B2(n_39),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_83),
.B1(n_7),
.B2(n_8),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_88),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_3),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_4),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_7),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_70),
.A2(n_5),
.B(n_6),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_5),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_10),
.C(n_12),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_97),
.B(n_98),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_99),
.A2(n_100),
.B1(n_25),
.B2(n_27),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_90),
.B(n_15),
.Y(n_106)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_29),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_20),
.C(n_22),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_110),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_108),
.Y(n_113)
);

OAI321xp33_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_93),
.A3(n_101),
.B1(n_100),
.B2(n_92),
.C(n_28),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_107),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_114),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

NAND2x1p5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_109),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_105),
.C(n_101),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_113),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_116),
.Y(n_121)
);


endmodule