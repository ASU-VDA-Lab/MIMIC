module real_jpeg_7218_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

BUFx10_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_1),
.B(n_5),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

AO22x1_ASAP7_75t_SL g14 ( 
.A1(n_3),
.A2(n_4),
.B1(n_15),
.B2(n_16),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

OA21x2_ASAP7_75t_L g20 ( 
.A1(n_4),
.A2(n_21),
.B(n_22),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_4),
.B(n_21),
.Y(n_22)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_SL g6 ( 
.A(n_7),
.B(n_29),
.Y(n_6)
);

OAI21xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_12),
.B(n_23),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_9),
.Y(n_8)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_9),
.B(n_24),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_11),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_13),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_17),
.B(n_19),
.Y(n_13)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_20),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);


endmodule