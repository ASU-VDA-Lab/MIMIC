module fake_jpeg_27594_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx5_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

AOI21xp33_ASAP7_75t_L g7 ( 
.A1(n_1),
.A2(n_2),
.B(n_0),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx2_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_L g14 ( 
.A1(n_7),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_14),
.A2(n_17),
.B1(n_18),
.B2(n_8),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_8),
.B(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_15),
.B(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_9),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_15),
.B(n_10),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_14),
.A2(n_12),
.B(n_6),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_23),
.B(n_16),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_25),
.B(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_22),
.Y(n_26)
);

OAI21x1_ASAP7_75t_R g27 ( 
.A1(n_21),
.A2(n_13),
.B(n_17),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_19),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_29),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_11),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_28),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_34),
.B1(n_32),
.B2(n_28),
.Y(n_35)
);

FAx1_ASAP7_75t_SL g34 ( 
.A(n_32),
.B(n_28),
.CI(n_31),
.CON(n_34),
.SN(n_34)
);

HAxp5_ASAP7_75t_SL g36 ( 
.A(n_35),
.B(n_34),
.CON(n_36),
.SN(n_36)
);


endmodule