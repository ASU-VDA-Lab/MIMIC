module fake_jpeg_10491_n_236 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_236);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx6_ASAP7_75t_SL g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_30),
.B(n_26),
.Y(n_49)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_29),
.A2(n_26),
.B1(n_14),
.B2(n_18),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_18),
.B1(n_14),
.B2(n_26),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_38),
.Y(n_56)
);

HB1xp67_ASAP7_75t_SL g81 ( 
.A(n_56),
.Y(n_81)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_18),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_43),
.Y(n_78)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_60),
.B(n_64),
.Y(n_84)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_33),
.B(n_30),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_42),
.B(n_62),
.Y(n_82)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_70),
.B1(n_24),
.B2(n_13),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_50),
.A2(n_23),
.B1(n_17),
.B2(n_21),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_68),
.A2(n_21),
.B1(n_17),
.B2(n_23),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_69),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_39),
.A2(n_14),
.B1(n_13),
.B2(n_24),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_63),
.C(n_55),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_76),
.B(n_88),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_27),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

NOR2x1p5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_69),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_43),
.C(n_46),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_94),
.B1(n_75),
.B2(n_64),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_91),
.B(n_93),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_83),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_98),
.B(n_99),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_42),
.B1(n_58),
.B2(n_54),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_53),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_87),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_76),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_71),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_102),
.Y(n_115)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_108),
.B(n_116),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_72),
.B(n_85),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_90),
.B1(n_100),
.B2(n_102),
.Y(n_133)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_113),
.Y(n_140)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_120),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_74),
.B(n_79),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_124),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_97),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_96),
.B(n_103),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_93),
.B(n_74),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_86),
.B(n_65),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_125),
.B(n_95),
.Y(n_135)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_86),
.B(n_88),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_106),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_99),
.C(n_96),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_132),
.C(n_136),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_128),
.B(n_137),
.Y(n_153)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_129),
.B(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_131),
.B(n_143),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_95),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_133),
.A2(n_135),
.B1(n_115),
.B2(n_117),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_90),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_13),
.B(n_24),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_47),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_111),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_114),
.A2(n_53),
.B1(n_60),
.B2(n_58),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_144),
.B1(n_112),
.B2(n_110),
.Y(n_152)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_107),
.A2(n_56),
.B1(n_41),
.B2(n_50),
.Y(n_144)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_142),
.Y(n_146)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_127),
.A2(n_115),
.B1(n_124),
.B2(n_111),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_151),
.B1(n_144),
.B2(n_138),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_159),
.C(n_160),
.Y(n_169)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_112),
.B1(n_17),
.B2(n_25),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_154),
.A2(n_25),
.B1(n_21),
.B2(n_22),
.Y(n_180)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_158),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_140),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_128),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_28),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_145),
.Y(n_162)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_162),
.Y(n_167)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_164),
.Y(n_165)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_157),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_168),
.A2(n_175),
.B(n_176),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_132),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_178),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_153),
.B(n_137),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_173),
.B(n_160),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_161),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_147),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_153),
.A2(n_22),
.B1(n_25),
.B2(n_23),
.Y(n_177)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_44),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_22),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_165),
.A2(n_152),
.B(n_154),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_181),
.A2(n_194),
.B(n_180),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_173),
.B(n_159),
.Y(n_182)
);

XNOR2x1_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_186),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_191),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_148),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_36),
.C(n_34),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_146),
.C(n_155),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_190),
.C(n_193),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_155),
.C(n_69),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_67),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_67),
.C(n_41),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_165),
.A2(n_9),
.B(n_12),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_166),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_202),
.C(n_203),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_167),
.Y(n_196)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_183),
.A2(n_179),
.B1(n_171),
.B2(n_177),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_197),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_198),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_170),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_201),
.B(n_193),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_190),
.A2(n_8),
.B(n_9),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_20),
.C(n_19),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_186),
.C(n_189),
.Y(n_208)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_208),
.B(n_210),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_182),
.C(n_20),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_6),
.B1(n_11),
.B2(n_10),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_211),
.A2(n_204),
.B1(n_200),
.B2(n_7),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_205),
.A2(n_6),
.B(n_11),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_213),
.A2(n_214),
.B(n_9),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_199),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_217),
.Y(n_223)
);

OAI211xp5_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_12),
.B(n_6),
.C(n_7),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_4),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_207),
.A2(n_7),
.B(n_11),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_219),
.A2(n_218),
.B(n_213),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_4),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_224),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_221),
.B(n_212),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_226),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_223),
.A2(n_216),
.B(n_10),
.Y(n_227)
);

XOR2x2_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_12),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_231),
.C(n_229),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_228),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_232),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_233),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_1),
.C(n_3),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_3),
.Y(n_236)
);


endmodule