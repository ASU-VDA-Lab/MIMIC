module fake_jpeg_16556_n_335 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_16),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_45),
.Y(n_66)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_46),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_26),
.B1(n_28),
.B2(n_33),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_48),
.B1(n_54),
.B2(n_70),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_28),
.B1(n_26),
.B2(n_33),
.Y(n_48)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_54)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_25),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_21),
.Y(n_95)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_20),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_18),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_38),
.A2(n_28),
.B1(n_26),
.B2(n_30),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_66),
.B(n_27),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_SL g111 ( 
.A(n_74),
.B(n_95),
.C(n_100),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_76),
.A2(n_34),
.B(n_22),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_67),
.B(n_18),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_77),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_30),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_51),
.Y(n_84)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_63),
.B(n_18),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_89),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_30),
.B1(n_43),
.B2(n_40),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_61),
.B1(n_27),
.B2(n_21),
.Y(n_127)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_20),
.Y(n_94)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_46),
.C(n_31),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_43),
.Y(n_120)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_20),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_98),
.A2(n_56),
.B1(n_60),
.B2(n_71),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_101),
.A2(n_117),
.B1(n_127),
.B2(n_130),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_29),
.B1(n_65),
.B2(n_64),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_73),
.B1(n_81),
.B2(n_90),
.Y(n_131)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_103),
.Y(n_143)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_74),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_113),
.B(n_23),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_74),
.A2(n_86),
.B(n_97),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_115),
.B(n_21),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_27),
.B(n_34),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_91),
.A2(n_69),
.B1(n_54),
.B2(n_29),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_32),
.Y(n_153)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_72),
.B(n_55),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_51),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_91),
.A2(n_29),
.B1(n_43),
.B2(n_40),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_133),
.B1(n_134),
.B2(n_138),
.Y(n_174)
);

O2A1O1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_120),
.A2(n_91),
.B(n_75),
.C(n_29),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_132),
.A2(n_153),
.B(n_129),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_73),
.B1(n_96),
.B2(n_97),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_99),
.B1(n_83),
.B2(n_87),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_31),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_142),
.C(n_124),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_110),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_152),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_79),
.B1(n_55),
.B2(n_84),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_17),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_135),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_147),
.B(n_115),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_22),
.B(n_34),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_127),
.A2(n_82),
.B1(n_22),
.B2(n_24),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_150),
.B1(n_108),
.B2(n_105),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_32),
.B1(n_24),
.B2(n_19),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_151),
.A2(n_123),
.B1(n_108),
.B2(n_125),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_106),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_164),
.B1(n_168),
.B2(n_175),
.Y(n_188)
);

OAI22x1_ASAP7_75t_SL g157 ( 
.A1(n_132),
.A2(n_139),
.B1(n_153),
.B2(n_146),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_166),
.B1(n_174),
.B2(n_161),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_126),
.Y(n_158)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_158),
.Y(n_208)
);

NOR2xp67_ASAP7_75t_R g186 ( 
.A(n_159),
.B(n_151),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_160),
.B(n_169),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_153),
.Y(n_161)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_142),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_101),
.B1(n_117),
.B2(n_112),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_112),
.C(n_130),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_167),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_121),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_166),
.A2(n_178),
.B1(n_165),
.B2(n_174),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_132),
.A2(n_109),
.B(n_121),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_140),
.A2(n_153),
.B1(n_134),
.B2(n_131),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_140),
.B(n_109),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_173),
.C(n_24),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_124),
.B(n_118),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_103),
.B1(n_118),
.B2(n_110),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_176),
.A2(n_181),
.B1(n_32),
.B2(n_19),
.Y(n_206)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_179),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_128),
.B(n_107),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_180),
.B(n_143),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_107),
.B1(n_11),
.B2(n_12),
.Y(n_181)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_137),
.Y(n_184)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_186),
.B(n_189),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_157),
.A2(n_138),
.A3(n_155),
.B1(n_143),
.B2(n_24),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_187),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_207),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_157),
.A2(n_149),
.B1(n_106),
.B2(n_141),
.Y(n_192)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_167),
.Y(n_194)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_141),
.Y(n_195)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_149),
.Y(n_196)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_181),
.C(n_162),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_162),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_199),
.B(n_179),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_17),
.Y(n_200)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_164),
.A2(n_180),
.B1(n_165),
.B2(n_156),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_201),
.A2(n_206),
.B1(n_166),
.B2(n_168),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_175),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_32),
.Y(n_229)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_17),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_209),
.A2(n_221),
.B1(n_229),
.B2(n_233),
.Y(n_255)
);

INVxp33_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_220),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_171),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_198),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_173),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_227),
.C(n_183),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_160),
.B1(n_176),
.B2(n_159),
.Y(n_221)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_195),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_226),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_197),
.Y(n_225)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_197),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_182),
.B(n_16),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_190),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_188),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_214),
.A2(n_206),
.B1(n_194),
.B2(n_190),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_234),
.Y(n_267)
);

NOR3xp33_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_186),
.C(n_202),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_250),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_239),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_201),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_207),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_244),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_189),
.B(n_184),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_242),
.A2(n_233),
.B(n_251),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_253),
.C(n_254),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_210),
.B(n_192),
.Y(n_244)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_187),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_248),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_210),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_252),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_208),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_212),
.B(n_208),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_214),
.A2(n_185),
.B1(n_199),
.B2(n_203),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_185),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_203),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_L g257 ( 
.A1(n_244),
.A2(n_231),
.B(n_212),
.C(n_217),
.Y(n_257)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_216),
.C(n_231),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_268),
.C(n_273),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_236),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_262),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_253),
.A2(n_211),
.B1(n_224),
.B2(n_213),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_264),
.A2(n_248),
.B1(n_246),
.B2(n_239),
.Y(n_276)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_269),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_211),
.C(n_193),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_238),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_270),
.B(n_273),
.Y(n_289)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_271),
.B(n_14),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_204),
.C(n_19),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_276),
.B(n_286),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_255),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_289),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_251),
.C(n_19),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_281),
.C(n_288),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_280),
.A2(n_257),
.B(n_2),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_256),
.C(n_263),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_3),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_285),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_258),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_10),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_270),
.C(n_274),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_17),
.C(n_2),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_272),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_298),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_275),
.A2(n_262),
.B1(n_267),
.B2(n_259),
.Y(n_292)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_274),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_297),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_272),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_266),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_302),
.C(n_277),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_6),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_283),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_303),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_17),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_17),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_293),
.A2(n_284),
.B(n_288),
.Y(n_306)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_306),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_279),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_307),
.B(n_311),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_302),
.A2(n_4),
.B(n_5),
.Y(n_310)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_310),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_294),
.A2(n_4),
.B(n_5),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_6),
.Y(n_317)
);

A2O1A1O1Ixp25_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_299),
.B(n_298),
.C(n_290),
.D(n_291),
.Y(n_315)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_315),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_317),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_309),
.B(n_290),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_313),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_7),
.C(n_8),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_SL g322 ( 
.A(n_308),
.B(n_307),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_305),
.B(n_308),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_323),
.A2(n_324),
.B(n_327),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_316),
.A2(n_313),
.B(n_8),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_328),
.A2(n_316),
.B(n_319),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_325),
.C(n_329),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_326),
.C(n_320),
.Y(n_332)
);

A2O1A1Ixp33_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_333)
);

O2A1O1Ixp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_9),
.Y(n_335)
);


endmodule