module fake_jpeg_3130_n_348 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_348);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_348;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_1),
.B(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_13),
.B(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_49),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_56),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_52),
.Y(n_140)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_54),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_28),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_61),
.B(n_64),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_21),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_81),
.Y(n_110)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_28),
.Y(n_64)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_68),
.Y(n_144)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_28),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_70),
.B(n_71),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g139 ( 
.A(n_74),
.Y(n_139)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_76),
.Y(n_155)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_83),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_79),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_21),
.B(n_0),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_22),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_87),
.B(n_88),
.Y(n_146)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_48),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_91),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_90),
.B(n_96),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_44),
.B(n_1),
.Y(n_91)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

HAxp5_ASAP7_75t_SL g117 ( 
.A(n_92),
.B(n_102),
.CON(n_117),
.SN(n_117)
);

INVx6_ASAP7_75t_SL g93 ( 
.A(n_25),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_94),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_48),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_22),
.B(n_1),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_99),
.Y(n_136)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_97),
.B(n_98),
.Y(n_107)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_27),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_101),
.Y(n_137)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_47),
.B(n_40),
.Y(n_106)
);

INVx2_ASAP7_75t_R g184 ( 
.A(n_106),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_36),
.B1(n_46),
.B2(n_43),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_108),
.A2(n_112),
.B1(n_118),
.B2(n_121),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_74),
.B1(n_82),
.B2(n_77),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_93),
.A2(n_36),
.B1(n_46),
.B2(n_43),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g174 ( 
.A1(n_113),
.A2(n_123),
.B1(n_133),
.B2(n_151),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_76),
.A2(n_35),
.B1(n_27),
.B2(n_38),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_55),
.A2(n_35),
.B1(n_40),
.B2(n_38),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_47),
.B1(n_37),
.B2(n_7),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_67),
.A2(n_37),
.B1(n_4),
.B2(n_8),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_124),
.A2(n_139),
.B1(n_149),
.B2(n_144),
.Y(n_181)
);

AND2x2_ASAP7_75t_SL g127 ( 
.A(n_58),
.B(n_2),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_127),
.B(n_91),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_2),
.B1(n_8),
.B2(n_11),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_128),
.A2(n_123),
.B1(n_116),
.B2(n_131),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_84),
.A2(n_8),
.B1(n_12),
.B2(n_14),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_98),
.B(n_14),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_141),
.B(n_150),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_15),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_65),
.A2(n_80),
.B1(n_60),
.B2(n_53),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_100),
.B(n_69),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_152),
.B(n_66),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_85),
.A2(n_90),
.B1(n_87),
.B2(n_68),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_109),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_110),
.B(n_72),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_159),
.B(n_160),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_73),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_137),
.A2(n_79),
.B1(n_92),
.B2(n_57),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_162),
.Y(n_203)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_163),
.Y(n_231)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_167),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_166),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_105),
.B(n_129),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_107),
.A2(n_146),
.B1(n_156),
.B2(n_147),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_168),
.Y(n_220)
);

BUFx12_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_106),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_197),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_127),
.A2(n_133),
.B1(n_113),
.B2(n_157),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_172),
.A2(n_177),
.B1(n_181),
.B2(n_189),
.Y(n_206)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_173),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_153),
.B1(n_134),
.B2(n_111),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_175),
.A2(n_180),
.B1(n_185),
.B2(n_191),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_122),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_178),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_145),
.A2(n_116),
.B1(n_139),
.B2(n_130),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_140),
.A2(n_138),
.B1(n_109),
.B2(n_143),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_120),
.C(n_114),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_182),
.Y(n_205)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_124),
.A2(n_149),
.B1(n_144),
.B2(n_115),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_140),
.B(n_142),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_186),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g187 ( 
.A(n_103),
.B(n_104),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_199),
.Y(n_226)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_126),
.Y(n_188)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_190),
.Y(n_221)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_126),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_192),
.Y(n_222)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_131),
.Y(n_193)
);

INVx13_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_194),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_117),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_195),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_138),
.A2(n_117),
.B1(n_154),
.B2(n_125),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_196),
.A2(n_194),
.B(n_191),
.Y(n_201)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_125),
.Y(n_197)
);

INVx6_ASAP7_75t_SL g198 ( 
.A(n_104),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_200),
.Y(n_216)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_111),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_172),
.A2(n_171),
.B(n_198),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_208),
.Y(n_237)
);

AND2x6_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_168),
.Y(n_215)
);

A2O1A1O1Ixp25_ASAP7_75t_L g244 ( 
.A1(n_215),
.A2(n_218),
.B(n_174),
.C(n_169),
.D(n_164),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_199),
.A2(n_187),
.B(n_174),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_217),
.B(n_225),
.Y(n_257)
);

AND2x6_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_199),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_161),
.B(n_187),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_216),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_234),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_220),
.A2(n_179),
.B1(n_181),
.B2(n_177),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_233),
.A2(n_238),
.B1(n_221),
.B2(n_231),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_216),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_204),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_235),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_220),
.A2(n_174),
.B1(n_193),
.B2(n_183),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_222),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_249),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_217),
.A2(n_174),
.B1(n_166),
.B2(n_173),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_241),
.A2(n_245),
.B1(n_252),
.B2(n_255),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_178),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_207),
.Y(n_243)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_243),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_244),
.A2(n_228),
.B(n_231),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_208),
.A2(n_170),
.B1(n_163),
.B2(n_190),
.Y(n_245)
);

AND2x6_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_215),
.Y(n_246)
);

AOI322xp5_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_209),
.A3(n_219),
.B1(n_223),
.B2(n_228),
.C1(n_230),
.C2(n_257),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_210),
.B(n_214),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_247),
.B(n_251),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_169),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_248),
.B(n_257),
.Y(n_275)
);

AO22x1_ASAP7_75t_SL g249 ( 
.A1(n_206),
.A2(n_197),
.B1(n_211),
.B2(n_226),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_212),
.Y(n_250)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_202),
.B(n_205),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_206),
.A2(n_201),
.B1(n_211),
.B2(n_227),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_205),
.B(n_225),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_253),
.B(n_254),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_222),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_229),
.A2(n_224),
.B1(n_203),
.B2(n_227),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_203),
.A2(n_229),
.B1(n_221),
.B2(n_213),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_209),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_263),
.Y(n_280)
);

NAND3xp33_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_236),
.C(n_232),
.Y(n_283)
);

OA22x2_ASAP7_75t_L g263 ( 
.A1(n_238),
.A2(n_212),
.B1(n_213),
.B2(n_219),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_277),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_236),
.A2(n_209),
.B(n_230),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_245),
.B(n_244),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_240),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_271),
.Y(n_279)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_239),
.Y(n_272)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_273),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_274),
.B(n_241),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_275),
.B(n_246),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_256),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_276),
.A2(n_237),
.B1(n_233),
.B2(n_234),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_282),
.A2(n_284),
.B1(n_258),
.B2(n_261),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_283),
.A2(n_294),
.B(n_259),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_276),
.A2(n_277),
.B1(n_267),
.B2(n_270),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_249),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_290),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_288),
.A2(n_268),
.B(n_264),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_250),
.Y(n_289)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_289),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_249),
.Y(n_290)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_271),
.Y(n_291)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_252),
.Y(n_292)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_248),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_266),
.C(n_269),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_296),
.B(n_278),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_305),
.C(n_307),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_298),
.A2(n_303),
.B1(n_309),
.B2(n_294),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_300),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_284),
.A2(n_278),
.B1(n_262),
.B2(n_265),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_265),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_306),
.B(n_279),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_282),
.A2(n_266),
.B1(n_269),
.B2(n_272),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_285),
.A2(n_263),
.B1(n_273),
.B2(n_290),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_310),
.A2(n_280),
.B1(n_287),
.B2(n_292),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_293),
.C(n_288),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_297),
.C(n_305),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_313),
.A2(n_316),
.B(n_318),
.Y(n_321)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_301),
.Y(n_314)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_314),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_299),
.B(n_279),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_317),
.Y(n_323)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_302),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_303),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_319),
.B(n_310),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_320),
.B(n_298),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_324),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_312),
.C(n_315),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_325),
.B(n_327),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_304),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_316),
.A2(n_306),
.B(n_300),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_311),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_328),
.Y(n_335)
);

OAI21xp33_ASAP7_75t_L g332 ( 
.A1(n_323),
.A2(n_320),
.B(n_304),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_332),
.B(n_334),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_321),
.B(n_317),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_319),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_336),
.Y(n_341)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_329),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_314),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_L g340 ( 
.A1(n_337),
.A2(n_308),
.B(n_322),
.C(n_291),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_339),
.A2(n_330),
.B(n_338),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_340),
.B(n_342),
.Y(n_344)
);

AOI322xp5_ASAP7_75t_L g343 ( 
.A1(n_341),
.A2(n_338),
.A3(n_318),
.B1(n_280),
.B2(n_286),
.C1(n_295),
.C2(n_326),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_343),
.B(n_281),
.Y(n_345)
);

AO21x1_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_344),
.B(n_281),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_346),
.B(n_309),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_347),
.A2(n_295),
.B(n_286),
.Y(n_348)
);


endmodule