module fake_jpeg_29449_n_420 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_420);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_420;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_4),
.B(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_50),
.B(n_55),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_63),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g52 ( 
.A(n_25),
.B(n_0),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_88),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_54),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_58),
.Y(n_153)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_14),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_67),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_16),
.B(n_13),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_21),
.B(n_13),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_70),
.B(n_71),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_21),
.B(n_23),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_77),
.Y(n_125)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

BUFx10_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_80),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_25),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_82),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_23),
.B(n_13),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_90),
.Y(n_110)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

NAND2x1_ASAP7_75t_L g88 ( 
.A(n_25),
.B(n_0),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_95),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_36),
.B(n_11),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_36),
.B(n_10),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_91),
.B(n_94),
.Y(n_143)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_18),
.B(n_0),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_34),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_69),
.A2(n_35),
.B1(n_29),
.B2(n_47),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_107),
.A2(n_118),
.B1(n_121),
.B2(n_123),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_93),
.A2(n_29),
.B1(n_44),
.B2(n_47),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_70),
.B(n_32),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_119),
.B(n_135),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_84),
.A2(n_29),
.B1(n_44),
.B2(n_30),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_30),
.B1(n_42),
.B2(n_38),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_59),
.A2(n_33),
.B1(n_42),
.B2(n_38),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_127),
.A2(n_134),
.B1(n_148),
.B2(n_150),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_52),
.A2(n_46),
.B(n_37),
.C(n_18),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_96),
.B(n_64),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g133 ( 
.A1(n_88),
.A2(n_46),
.B(n_37),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_133),
.B(n_58),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_57),
.A2(n_45),
.B1(n_40),
.B2(n_32),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_73),
.B(n_45),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_73),
.B(n_40),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_149),
.Y(n_172)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_65),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_76),
.A2(n_41),
.B1(n_3),
.B2(n_6),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_159),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_106),
.B(n_79),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_156),
.B(n_115),
.C(n_152),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_124),
.Y(n_157)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_167),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_132),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_160),
.Y(n_222)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_161),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_106),
.B(n_89),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_165),
.Y(n_205)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_164),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_106),
.B(n_110),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_129),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_103),
.Y(n_168)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_89),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_169),
.B(n_178),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_128),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_170),
.Y(n_199)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

OA22x2_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_87),
.B1(n_80),
.B2(n_82),
.Y(n_173)
);

OA21x2_ASAP7_75t_L g229 ( 
.A1(n_173),
.A2(n_186),
.B(n_190),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_102),
.B(n_41),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_174),
.B(n_185),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_125),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_82),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_75),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_184),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_120),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_182),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_116),
.B(n_75),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_112),
.B(n_41),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_150),
.A2(n_53),
.B(n_61),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_111),
.B(n_80),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_189),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_114),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_100),
.B(n_78),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_134),
.A2(n_54),
.B(n_3),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_113),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_191),
.Y(n_223)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_131),
.Y(n_192)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_103),
.Y(n_195)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_173),
.A2(n_147),
.B1(n_99),
.B2(n_139),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_206),
.A2(n_214),
.B1(n_186),
.B2(n_163),
.Y(n_235)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_165),
.A2(n_104),
.B(n_115),
.C(n_141),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_208),
.B(n_184),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_147),
.B1(n_99),
.B2(n_139),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_173),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_173),
.Y(n_231)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_154),
.Y(n_225)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_156),
.C(n_162),
.Y(n_232)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_154),
.Y(n_230)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_230),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_231),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_232),
.B(n_244),
.Y(n_276)
);

AO22x1_ASAP7_75t_L g233 ( 
.A1(n_229),
.A2(n_208),
.B1(n_190),
.B2(n_203),
.Y(n_233)
);

AO22x1_ASAP7_75t_SL g260 ( 
.A1(n_233),
.A2(n_255),
.B1(n_198),
.B2(n_210),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_235),
.A2(n_233),
.B1(n_249),
.B2(n_255),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_223),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_236),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_191),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_237),
.B(n_245),
.Y(n_266)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_189),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_240),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_220),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_241),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_242),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_203),
.A2(n_155),
.B(n_187),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_199),
.B(n_167),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_202),
.B(n_166),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_246),
.Y(n_282)
);

BUFx8_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_181),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_250),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_229),
.A2(n_156),
.B1(n_175),
.B2(n_170),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_249),
.A2(n_197),
.B1(n_182),
.B2(n_219),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_169),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_178),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_252),
.Y(n_274)
);

MAJx2_ASAP7_75t_L g253 ( 
.A(n_196),
.B(n_205),
.C(n_227),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_258),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_SL g255 ( 
.A1(n_229),
.A2(n_214),
.B(n_205),
.C(n_201),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_228),
.Y(n_256)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_172),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_260),
.B(n_263),
.Y(n_288)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_261),
.Y(n_287)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_265),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_272),
.B1(n_278),
.B2(n_284),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_233),
.A2(n_236),
.B(n_240),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_273),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_235),
.A2(n_197),
.B1(n_212),
.B2(n_210),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_255),
.A2(n_207),
.B1(n_200),
.B2(n_224),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_255),
.A2(n_109),
.B1(n_216),
.B2(n_200),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_254),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_255),
.A2(n_209),
.B1(n_198),
.B2(n_207),
.Y(n_278)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_254),
.Y(n_283)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_283),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_244),
.A2(n_209),
.B1(n_193),
.B2(n_176),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_258),
.Y(n_286)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_286),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_283),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_289),
.B(n_296),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_290),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_251),
.Y(n_291)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_291),
.Y(n_318)
);

A2O1A1Ixp33_ASAP7_75t_L g292 ( 
.A1(n_270),
.A2(n_250),
.B(n_239),
.C(n_248),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_292),
.A2(n_256),
.B(n_268),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_247),
.Y(n_293)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_293),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_294),
.A2(n_211),
.B1(n_183),
.B2(n_157),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_253),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_297),
.C(n_267),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_232),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_257),
.C(n_234),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_264),
.B(n_257),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_299),
.Y(n_315)
);

XNOR2x1_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_247),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_284),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_301),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_277),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_294),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_247),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_304),
.B1(n_279),
.B2(n_275),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_275),
.A2(n_256),
.B1(n_234),
.B2(n_238),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_264),
.B(n_226),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_271),
.Y(n_320)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_281),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_308),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_309),
.B(n_329),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_285),
.A2(n_260),
.B1(n_263),
.B2(n_281),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_311),
.A2(n_314),
.B1(n_325),
.B2(n_288),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_290),
.A2(n_260),
.B1(n_279),
.B2(n_259),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_312),
.B(n_310),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_302),
.A2(n_268),
.B1(n_271),
.B2(n_267),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_321),
.C(n_326),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_300),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_204),
.C(n_225),
.Y(n_321)
);

AO21x1_ASAP7_75t_L g339 ( 
.A1(n_323),
.A2(n_324),
.B(n_288),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_302),
.A2(n_241),
.B1(n_222),
.B2(n_160),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_297),
.B(n_204),
.C(n_230),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_300),
.A2(n_228),
.B(n_213),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_327),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_296),
.B(n_211),
.C(n_183),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_320),
.Y(n_343)
);

INVxp33_ASAP7_75t_SL g330 ( 
.A(n_299),
.Y(n_330)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_330),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_319),
.B(n_305),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_333),
.B(n_334),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_300),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_338),
.C(n_346),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_315),
.B(n_292),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_339),
.B(n_343),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_340),
.A2(n_345),
.B1(n_324),
.B2(n_329),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_306),
.Y(n_342)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_342),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_306),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_344),
.B(n_349),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_313),
.A2(n_307),
.B1(n_287),
.B2(n_308),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_315),
.B(n_298),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_321),
.B(n_287),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_347),
.B(n_350),
.C(n_307),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_348),
.A2(n_140),
.B1(n_157),
.B2(n_177),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_317),
.B(n_316),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_328),
.B(n_314),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_324),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_168),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_354),
.A2(n_338),
.B1(n_347),
.B2(n_346),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_SL g355 ( 
.A(n_337),
.B(n_322),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_355),
.B(n_356),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_348),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_351),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_358),
.B(n_363),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_322),
.Y(n_359)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_359),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_325),
.C(n_195),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_361),
.B(n_367),
.C(n_334),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_336),
.A2(n_140),
.B1(n_144),
.B2(n_138),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_333),
.B(n_192),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_364),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_365),
.B(n_161),
.Y(n_379)
);

XNOR2x1_ASAP7_75t_L g372 ( 
.A(n_366),
.B(n_335),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_341),
.B(n_179),
.C(n_164),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_368),
.B(n_370),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_369),
.B(n_372),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_357),
.A2(n_339),
.B(n_332),
.Y(n_371)
);

AOI21x1_ASAP7_75t_L g388 ( 
.A1(n_371),
.A2(n_151),
.B(n_105),
.Y(n_388)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_362),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_374),
.B(n_375),
.Y(n_383)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_365),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_377),
.B(n_353),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_379),
.B(n_361),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_358),
.B(n_142),
.C(n_141),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_380),
.B(n_367),
.C(n_353),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_374),
.B(n_352),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_386),
.Y(n_400)
);

NOR2x1_ASAP7_75t_L g384 ( 
.A(n_371),
.B(n_360),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_384),
.A2(n_388),
.B(n_379),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_385),
.B(n_387),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_373),
.B(n_124),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_390),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_378),
.B(n_160),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_391),
.B(n_392),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_369),
.B(n_131),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_381),
.A2(n_380),
.B(n_375),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_393),
.A2(n_386),
.B(n_389),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_383),
.B(n_377),
.Y(n_394)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_394),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_389),
.B(n_376),
.C(n_372),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_395),
.B(n_153),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_399),
.B(n_401),
.Y(n_405)
);

AOI21x1_ASAP7_75t_L g401 ( 
.A1(n_384),
.A2(n_376),
.B(n_151),
.Y(n_401)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_403),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_400),
.A2(n_388),
.B(n_138),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_404),
.A2(n_406),
.B(n_407),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_396),
.B(n_105),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_395),
.B(n_108),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_408),
.A2(n_122),
.B1(n_153),
.B2(n_108),
.Y(n_412)
);

O2A1O1Ixp33_ASAP7_75t_SL g409 ( 
.A1(n_405),
.A2(n_398),
.B(n_397),
.C(n_396),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_409),
.A2(n_2),
.B(n_6),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_412),
.Y(n_413)
);

NOR3xp33_ASAP7_75t_L g414 ( 
.A(n_411),
.B(n_402),
.C(n_407),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_414),
.A2(n_415),
.B1(n_410),
.B2(n_9),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_416),
.B(n_417),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_413),
.B(n_122),
.C(n_2),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_418),
.B(n_9),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_419),
.B(n_9),
.Y(n_420)
);


endmodule