module fake_jpeg_13974_n_67 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_67);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_67;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_66;

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx10_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

INVx13_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx13_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx11_ASAP7_75t_SL g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_18),
.C(n_21),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_19),
.B(n_20),
.Y(n_22)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_9),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_12),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_23),
.B(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_27),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_21),
.B1(n_16),
.B2(n_19),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_16),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_18),
.B1(n_17),
.B2(n_21),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_33),
.A2(n_34),
.B1(n_35),
.B2(n_16),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_18),
.B1(n_17),
.B2(n_21),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_16),
.B1(n_19),
.B2(n_9),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_4),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_8),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_45),
.Y(n_51)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_32),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_48),
.Y(n_52)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_42),
.C(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_55),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_34),
.B(n_9),
.C(n_11),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_45),
.B1(n_20),
.B2(n_15),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_19),
.C(n_16),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_9),
.B(n_11),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_20),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_58),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_61),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_60),
.C(n_58),
.Y(n_64)
);

MAJx2_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_63),
.C(n_61),
.Y(n_65)
);

AOI322xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_5),
.A3(n_6),
.B1(n_10),
.B2(n_11),
.C1(n_59),
.C2(n_50),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_5),
.Y(n_67)
);


endmodule