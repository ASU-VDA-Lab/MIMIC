module fake_jpeg_31349_n_297 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_297);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_46),
.Y(n_74)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_18),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_62),
.Y(n_84)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_35),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

HAxp5_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_0),
.CON(n_54),
.SN(n_54)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_55),
.Y(n_93)
);

BUFx12f_ASAP7_75t_SL g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_22),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_39),
.Y(n_68)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVxp67_ASAP7_75t_SL g62 ( 
.A(n_26),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_36),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_39),
.B1(n_38),
.B2(n_19),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_66),
.A2(n_90),
.B1(n_98),
.B2(n_5),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_1),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_57),
.B(n_28),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_69),
.B(n_78),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_39),
.B1(n_31),
.B2(n_34),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_70),
.A2(n_81),
.B1(n_33),
.B2(n_2),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_19),
.B1(n_29),
.B2(n_20),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_43),
.B1(n_36),
.B2(n_33),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_49),
.B(n_28),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_63),
.B1(n_51),
.B2(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_34),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_91),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_88),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_31),
.B1(n_21),
.B2(n_24),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_32),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_32),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_96),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_24),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_101),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_45),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_60),
.A2(n_19),
.B1(n_20),
.B2(n_29),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_48),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_100),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_20),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_40),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_102),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_52),
.B(n_16),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_103),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_52),
.B(n_40),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_104),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_66),
.A2(n_20),
.B1(n_30),
.B2(n_23),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_105),
.A2(n_133),
.B1(n_136),
.B2(n_139),
.Y(n_147)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_68),
.B(n_1),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_108),
.B(n_8),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_111),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_30),
.B(n_23),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_112),
.A2(n_131),
.B(n_84),
.Y(n_149)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_33),
.B1(n_56),
.B2(n_3),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_117),
.B(n_119),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_93),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_127),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_95),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_132),
.Y(n_142)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_130),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_3),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_76),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_135),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_73),
.A2(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_83),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_141),
.B(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

NAND2xp33_ASAP7_75t_SL g144 ( 
.A(n_114),
.B(n_101),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_144),
.A2(n_134),
.B(n_122),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_149),
.Y(n_187)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_74),
.A3(n_94),
.B1(n_98),
.B2(n_77),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_164),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_77),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_158),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_133),
.A2(n_73),
.B1(n_99),
.B2(n_86),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_162),
.B1(n_87),
.B2(n_128),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_108),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_76),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_117),
.A2(n_99),
.B1(n_72),
.B2(n_86),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_97),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_72),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_166),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_129),
.B(n_11),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_138),
.B(n_11),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_12),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_165),
.C(n_141),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_195),
.C(n_145),
.Y(n_203)
);

AO22x1_ASAP7_75t_L g173 ( 
.A1(n_144),
.A2(n_163),
.B1(n_150),
.B2(n_140),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_SL g217 ( 
.A1(n_173),
.A2(n_12),
.B(n_13),
.C(n_16),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_147),
.A2(n_123),
.B1(n_137),
.B2(n_87),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_174),
.A2(n_152),
.B1(n_155),
.B2(n_151),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_163),
.A2(n_109),
.B1(n_106),
.B2(n_132),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_182),
.B1(n_194),
.B2(n_197),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_163),
.A2(n_112),
.B(n_131),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g219 ( 
.A1(n_177),
.A2(n_179),
.B1(n_190),
.B2(n_173),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_131),
.B1(n_139),
.B2(n_113),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_159),
.A2(n_107),
.B1(n_120),
.B2(n_130),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_143),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_185),
.B(n_189),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_119),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_145),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_188),
.B(n_152),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_142),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_126),
.B1(n_135),
.B2(n_125),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_142),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_192),
.B(n_196),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_161),
.A2(n_115),
.B(n_121),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_193),
.A2(n_146),
.B(n_153),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_85),
.B1(n_124),
.B2(n_14),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_85),
.C(n_15),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_166),
.A2(n_154),
.B1(n_148),
.B2(n_160),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_198),
.B(n_186),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_169),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_199),
.B(n_212),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_207),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_213),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_186),
.B(n_180),
.Y(n_231)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_146),
.C(n_153),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_216),
.C(n_187),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_207),
.B1(n_204),
.B2(n_211),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_152),
.Y(n_212)
);

AOI322xp5_ASAP7_75t_L g214 ( 
.A1(n_173),
.A2(n_178),
.A3(n_184),
.B1(n_188),
.B2(n_183),
.C1(n_192),
.C2(n_189),
.Y(n_214)
);

AOI221xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_217),
.B1(n_197),
.B2(n_184),
.C(n_170),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_151),
.C(n_155),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_218),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_190),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_170),
.A2(n_178),
.B1(n_177),
.B2(n_182),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_220),
.A2(n_179),
.B1(n_196),
.B2(n_195),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_201),
.A2(n_193),
.B(n_176),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_232),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_240),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_210),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_225),
.B(n_221),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_235),
.C(n_221),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_229),
.Y(n_245)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_217),
.A2(n_181),
.B(n_191),
.Y(n_232)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_216),
.C(n_203),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_239),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_220),
.Y(n_237)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_204),
.Y(n_238)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_238),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_206),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_219),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_247),
.C(n_248),
.Y(n_266)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

AOI21xp33_ASAP7_75t_L g246 ( 
.A1(n_230),
.A2(n_217),
.B(n_213),
.Y(n_246)
);

NOR3xp33_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_228),
.C(n_232),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_227),
.C(n_234),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_219),
.C(n_215),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_219),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_229),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_215),
.C(n_205),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_252),
.B(n_239),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_222),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_259),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_262),
.B(n_263),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_241),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_242),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_267),
.C(n_248),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_228),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_261),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_250),
.A2(n_231),
.B(n_223),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_254),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_265),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_238),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_270),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_252),
.C(n_253),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_256),
.A2(n_240),
.B1(n_245),
.B2(n_244),
.Y(n_271)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_271),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_264),
.A2(n_229),
.B1(n_245),
.B2(n_249),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_262),
.Y(n_277)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_277),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_266),
.B(n_257),
.Y(n_278)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_278),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_266),
.C(n_222),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_279),
.B(n_270),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_272),
.A2(n_226),
.B(n_236),
.Y(n_281)
);

OAI21x1_ASAP7_75t_SL g287 ( 
.A1(n_281),
.A2(n_271),
.B(n_275),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_226),
.B(n_274),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_276),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_288),
.Y(n_291)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_287),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_286),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_292),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_280),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_289),
.A2(n_284),
.B(n_282),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_294),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_291),
.B1(n_293),
.B2(n_292),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_281),
.Y(n_297)
);


endmodule