module fake_jpeg_2638_n_228 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_228);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_26),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_13),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_11),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_8),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_14),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_52),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_82),
.B(n_84),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_21),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_0),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_57),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_81),
.A2(n_70),
.B1(n_73),
.B2(n_63),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_91),
.A2(n_95),
.B1(n_69),
.B2(n_55),
.Y(n_107)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_65),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_63),
.B1(n_61),
.B2(n_70),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_64),
.B1(n_73),
.B2(n_67),
.Y(n_96)
);

AOI22x1_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_100),
.B1(n_69),
.B2(n_55),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_99),
.B(n_58),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_64),
.B1(n_66),
.B2(n_56),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_102),
.B(n_104),
.Y(n_137)
);

BUFx24_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_62),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_106),
.B(n_114),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_109),
.Y(n_123)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_115),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_112),
.B(n_117),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_76),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_90),
.Y(n_117)
);

CKINVDCx6p67_ASAP7_75t_R g118 ( 
.A(n_100),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_118),
.Y(n_122)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_120),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_75),
.B(n_77),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_89),
.C(n_85),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_136),
.C(n_139),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_118),
.B(n_89),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_127),
.B(n_132),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_118),
.A2(n_80),
.B1(n_77),
.B2(n_72),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_134),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_24),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_131),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_25),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_108),
.B(n_0),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_27),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_107),
.A2(n_80),
.B1(n_72),
.B2(n_54),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_140),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g136 ( 
.A1(n_103),
.A2(n_54),
.B(n_87),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_74),
.B(n_2),
.C(n_4),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_87),
.B(n_59),
.Y(n_139)
);

NOR3xp33_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_1),
.C(n_5),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_20),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_87),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_159),
.Y(n_170)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_147),
.Y(n_181)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_152),
.Y(n_183)
);

OAI21x1_ASAP7_75t_R g177 ( 
.A1(n_150),
.A2(n_156),
.B(n_37),
.Y(n_177)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_22),
.B1(n_46),
.B2(n_45),
.Y(n_151)
);

AOI22x1_ASAP7_75t_L g182 ( 
.A1(n_151),
.A2(n_157),
.B1(n_10),
.B2(n_12),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_125),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_1),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_154),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_5),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_49),
.B(n_41),
.C(n_40),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_6),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_7),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_165),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_166),
.Y(n_179)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_164),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_136),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_38),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_9),
.Y(n_167)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_123),
.C(n_135),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_162),
.C(n_151),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_163),
.A2(n_128),
.B1(n_11),
.B2(n_12),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_169),
.A2(n_182),
.B1(n_187),
.B2(n_16),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_146),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_173),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_166),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_184),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_144),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_163),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_188),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_181),
.B(n_161),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_199),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_191),
.C(n_197),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_151),
.C(n_157),
.Y(n_191)
);

FAx1_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_156),
.CI(n_148),
.CON(n_193),
.SN(n_193)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_193),
.B(n_178),
.Y(n_203)
);

OAI21x1_ASAP7_75t_SL g196 ( 
.A1(n_170),
.A2(n_15),
.B(n_16),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_196),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_175),
.B(n_36),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_187),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_208),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_203),
.B(n_190),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_174),
.B1(n_168),
.B2(n_169),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_206),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_195),
.A2(n_174),
.B1(n_176),
.B2(n_182),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_192),
.A2(n_177),
.B1(n_180),
.B2(n_172),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_185),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_211),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_204),
.A2(n_193),
.B(n_198),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_201),
.A2(n_191),
.B(n_31),
.Y(n_212)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

NOR2xp67_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_215),
.Y(n_220)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_209),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_209),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_218),
.C(n_220),
.Y(n_222)
);

A2O1A1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_217),
.A2(n_210),
.B(n_213),
.C(n_17),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_222),
.Y(n_223)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_223),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_224),
.A2(n_219),
.B1(n_23),
.B2(n_28),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_32),
.C(n_33),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_17),
.B(n_19),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_19),
.Y(n_228)
);


endmodule