module fake_jpeg_10744_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_10),
.A2(n_3),
.B(n_4),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_21),
.B(n_22),
.Y(n_30)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_20),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_2),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_3),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_5),
.Y(n_27)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_26),
.B1(n_7),
.B2(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_7),
.C(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_32),
.B1(n_19),
.B2(n_26),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_22),
.B1(n_17),
.B2(n_16),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_7),
.C(n_6),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_38),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_34),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_30),
.B1(n_33),
.B2(n_32),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_37),
.Y(n_41)
);

AOI21x1_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_42),
.B(n_40),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_38),
.C(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_34),
.Y(n_45)
);

BUFx24_ASAP7_75t_SL g46 ( 
.A(n_45),
.Y(n_46)
);


endmodule