module fake_jpeg_11796_n_101 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_101);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_7),
.B(n_34),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_0),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_50),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_0),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_53),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_1),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_59),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_51),
.A2(n_43),
.B1(n_38),
.B2(n_40),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_43),
.B1(n_38),
.B2(n_47),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_54),
.B(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_2),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_3),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_68),
.B1(n_75),
.B2(n_14),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_69),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_43),
.B1(n_38),
.B2(n_36),
.Y(n_68)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_4),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_58),
.A2(n_39),
.B(n_35),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_6),
.B(n_12),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_5),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_35),
.B1(n_8),
.B2(n_10),
.Y(n_75)
);

AO22x1_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_92)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_15),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_83),
.C(n_84),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_65),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_16),
.B(n_17),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_89),
.A2(n_90),
.B1(n_91),
.B2(n_78),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_76),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_80),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_98),
.A2(n_92),
.B(n_88),
.Y(n_99)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_99),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_96),
.Y(n_101)
);


endmodule