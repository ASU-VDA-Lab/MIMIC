module fake_jpeg_11882_n_517 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_517);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_517;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_12),
.B(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_53),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_55),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_57),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_32),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_59),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_108)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_31),
.B(n_3),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_64),
.B(n_95),
.Y(n_142)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_67),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_21),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_21),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_29),
.Y(n_113)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g128 ( 
.A(n_87),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx11_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_93),
.Y(n_145)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_31),
.B(n_3),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVx5_ASAP7_75t_SL g140 ( 
.A(n_97),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_99),
.B(n_100),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_106),
.B(n_125),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_108),
.A2(n_123),
.B1(n_42),
.B2(n_36),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_111),
.B(n_113),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_50),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_129),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_61),
.A2(n_48),
.B1(n_44),
.B2(n_38),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_80),
.B(n_34),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_94),
.Y(n_129)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_82),
.B(n_46),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_143),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_46),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_71),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_147),
.B(n_152),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_75),
.B(n_50),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_92),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_156),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_96),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_157),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_20),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_159),
.B(n_172),
.Y(n_214)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

INVx3_ASAP7_75t_SL g162 ( 
.A(n_140),
.Y(n_162)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_162),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_152),
.A2(n_100),
.B1(n_99),
.B2(n_88),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_165),
.A2(n_204),
.B1(n_154),
.B2(n_103),
.Y(n_211)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_110),
.Y(n_166)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_166),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_116),
.B(n_141),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_169),
.B(n_29),
.Y(n_248)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_171),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_42),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_173),
.Y(n_238)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_102),
.A2(n_83),
.B1(n_87),
.B2(n_86),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_175),
.A2(n_187),
.B1(n_205),
.B2(n_135),
.Y(n_247)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_176),
.Y(n_244)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_177),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_84),
.B1(n_77),
.B2(n_62),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_178),
.A2(n_181),
.B1(n_188),
.B2(n_195),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_185),
.Y(n_241)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_124),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_193),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_102),
.A2(n_49),
.B1(n_41),
.B2(n_25),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_145),
.A2(n_74),
.B1(n_48),
.B2(n_41),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_194),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_122),
.B(n_36),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_208),
.Y(n_218)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_138),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_191),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_103),
.A2(n_51),
.B1(n_76),
.B2(n_72),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_192),
.A2(n_135),
.B(n_134),
.Y(n_221)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_115),
.A2(n_41),
.B1(n_33),
.B2(n_20),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_139),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_130),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_115),
.A2(n_37),
.B1(n_40),
.B2(n_33),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_198),
.A2(n_128),
.B1(n_153),
.B2(n_107),
.Y(n_209)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_132),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_202),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_104),
.A2(n_40),
.B(n_37),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_117),
.Y(n_230)
);

INVx5_ASAP7_75t_SL g202 ( 
.A(n_140),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_148),
.B(n_81),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_206),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_158),
.A2(n_44),
.B1(n_98),
.B2(n_45),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_154),
.A2(n_49),
.B1(n_65),
.B2(n_73),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_144),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_133),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_207),
.B(n_126),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_107),
.B(n_4),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_209),
.A2(n_234),
.B1(n_237),
.B2(n_242),
.Y(n_270)
);

OA22x2_ASAP7_75t_L g274 ( 
.A1(n_211),
.A2(n_175),
.B1(n_185),
.B2(n_170),
.Y(n_274)
);

INVxp33_ASAP7_75t_L g254 ( 
.A(n_217),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_221),
.A2(n_247),
.B1(n_135),
.B2(n_78),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_169),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_248),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_172),
.B(n_144),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_232),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_230),
.B(n_161),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_159),
.B(n_118),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_181),
.A2(n_128),
.B1(n_105),
.B2(n_146),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_204),
.A2(n_118),
.B1(n_112),
.B2(n_153),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_235),
.A2(n_240),
.B1(n_160),
.B2(n_173),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_197),
.A2(n_120),
.B1(n_49),
.B2(n_146),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_208),
.A2(n_120),
.B1(n_150),
.B2(n_126),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_190),
.A2(n_28),
.B1(n_29),
.B2(n_78),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_164),
.B(n_28),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_245),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_28),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_246),
.Y(n_283)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_249),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_221),
.A2(n_167),
.B(n_180),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_251),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_218),
.B(n_174),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_252),
.B(n_259),
.Y(n_287)
);

AND2x6_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_202),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_253),
.B(n_265),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_258),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_211),
.A2(n_175),
.B1(n_192),
.B2(n_179),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_257),
.A2(n_275),
.B1(n_282),
.B2(n_219),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_226),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_201),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_226),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_260),
.B(n_264),
.Y(n_299)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_227),
.Y(n_261)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_261),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_214),
.B(n_203),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_262),
.B(n_233),
.Y(n_306)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_263),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_226),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_207),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_225),
.B(n_199),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_267),
.B(n_269),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_214),
.B(n_203),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_233),
.C(n_246),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_228),
.B(n_166),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_229),
.Y(n_271)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_271),
.Y(n_301)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_229),
.Y(n_272)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_272),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_232),
.B(n_176),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_273),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_270),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_235),
.A2(n_175),
.B1(n_179),
.B2(n_177),
.Y(n_275)
);

A2O1A1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_218),
.A2(n_182),
.B(n_162),
.C(n_186),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_276),
.A2(n_280),
.B(n_231),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_237),
.A2(n_209),
.B1(n_227),
.B2(n_213),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_277),
.A2(n_213),
.B1(n_215),
.B2(n_222),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_212),
.B(n_206),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_278),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_246),
.Y(n_279)
);

NAND3xp33_ASAP7_75t_SL g316 ( 
.A(n_279),
.B(n_258),
.C(n_260),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_233),
.Y(n_281)
);

INVx11_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_220),
.B(n_193),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_284),
.A2(n_223),
.B(n_254),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_242),
.B(n_29),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_285),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_268),
.C(n_262),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_288),
.A2(n_259),
.B1(n_274),
.B2(n_281),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_249),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_239),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_256),
.A2(n_240),
.B1(n_239),
.B2(n_241),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_296),
.A2(n_263),
.B1(n_271),
.B2(n_272),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_257),
.A2(n_275),
.B1(n_282),
.B2(n_266),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_297),
.A2(n_270),
.B1(n_256),
.B2(n_280),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_303),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_304),
.A2(n_316),
.B(n_319),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_306),
.B(n_244),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_307),
.B(n_251),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_283),
.A2(n_231),
.B1(n_238),
.B2(n_215),
.Y(n_309)
);

OAI21xp33_ASAP7_75t_SL g342 ( 
.A1(n_309),
.A2(n_319),
.B(n_291),
.Y(n_342)
);

INVx8_ASAP7_75t_L g310 ( 
.A(n_269),
.Y(n_310)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_310),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_284),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_312),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_278),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_265),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_250),
.Y(n_338)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_261),
.Y(n_315)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_315),
.Y(n_325)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_276),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_318),
.Y(n_333)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_266),
.Y(n_320)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_320),
.Y(n_330)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_321),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_322),
.B(n_353),
.C(n_302),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_323),
.A2(n_340),
.B1(n_342),
.B2(n_348),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_326),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_287),
.B(n_252),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_329),
.B(n_343),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_331),
.A2(n_295),
.B1(n_305),
.B2(n_301),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_276),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_332),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_267),
.Y(n_334)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_334),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_264),
.Y(n_335)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_335),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_308),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_336),
.B(n_310),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_279),
.Y(n_337)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_337),
.Y(n_368)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_338),
.Y(n_362)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_294),
.Y(n_339)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_339),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_289),
.B(n_262),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_341),
.B(n_347),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_250),
.Y(n_343)
);

INVx11_ASAP7_75t_L g344 ( 
.A(n_291),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_344),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_312),
.B(n_255),
.Y(n_345)
);

NAND3xp33_ASAP7_75t_L g382 ( 
.A(n_345),
.B(n_182),
.C(n_5),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_290),
.A2(n_253),
.B(n_283),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_346),
.A2(n_298),
.B(n_302),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_289),
.B(n_283),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_297),
.A2(n_253),
.B1(n_274),
.B2(n_285),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_288),
.A2(n_274),
.B1(n_210),
.B2(n_222),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_349),
.A2(n_304),
.B1(n_296),
.B2(n_295),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_351),
.B(n_286),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_317),
.B(n_274),
.Y(n_352)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_352),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_306),
.B(n_244),
.C(n_236),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_333),
.A2(n_298),
.B1(n_290),
.B2(n_304),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_356),
.A2(n_381),
.B1(n_340),
.B2(n_327),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_357),
.B(n_331),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_322),
.B(n_293),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_358),
.B(n_367),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_337),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_363),
.B(n_385),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_365),
.A2(n_313),
.B1(n_210),
.B2(n_238),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_375),
.C(n_378),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_338),
.B(n_308),
.Y(n_369)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_369),
.Y(n_393)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_372),
.Y(n_395)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_339),
.Y(n_373)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_373),
.Y(n_398)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_374),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_351),
.B(n_299),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_346),
.B(n_305),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_323),
.A2(n_301),
.B1(n_292),
.B2(n_294),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_380),
.A2(n_324),
.B1(n_332),
.B2(n_327),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_352),
.A2(n_292),
.B1(n_300),
.B2(n_315),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_382),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_345),
.B(n_236),
.Y(n_383)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_383),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_328),
.B(n_313),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_321),
.Y(n_386)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_386),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_328),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_387),
.B(n_334),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_389),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_390),
.A2(n_416),
.B1(n_371),
.B2(n_380),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_370),
.A2(n_332),
.B(n_354),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_397),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_368),
.B(n_330),
.Y(n_394)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_394),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_370),
.A2(n_354),
.B(n_326),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_SL g402 ( 
.A(n_367),
.B(n_353),
.C(n_335),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_402),
.B(n_365),
.C(n_373),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_366),
.B(n_341),
.C(n_347),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_409),
.C(n_412),
.Y(n_417)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_405),
.Y(n_433)
);

XNOR2x1_ASAP7_75t_L g418 ( 
.A(n_406),
.B(n_411),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_355),
.A2(n_336),
.B1(n_330),
.B2(n_324),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_410),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_368),
.B(n_325),
.Y(n_408)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_408),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_357),
.B(n_348),
.C(n_325),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_355),
.A2(n_350),
.B1(n_349),
.B2(n_344),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_358),
.B(n_171),
.C(n_168),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_375),
.B(n_191),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_413),
.B(n_364),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_384),
.A2(n_163),
.B1(n_183),
.B2(n_6),
.Y(n_414)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_414),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_361),
.Y(n_415)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_415),
.Y(n_439)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_361),
.Y(n_416)
);

FAx1_ASAP7_75t_L g419 ( 
.A(n_392),
.B(n_356),
.CI(n_376),
.CON(n_419),
.SN(n_419)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_419),
.A2(n_408),
.B(n_394),
.Y(n_449)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_421),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_400),
.B(n_378),
.C(n_362),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_424),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_423),
.B(n_427),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_400),
.B(n_381),
.C(n_386),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_403),
.B(n_360),
.C(n_364),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_429),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_390),
.B(n_376),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_409),
.B(n_399),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_428),
.B(n_406),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_399),
.B(n_359),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_413),
.B(n_371),
.C(n_359),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_430),
.B(n_434),
.C(n_417),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_432),
.B(n_407),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_412),
.B(n_379),
.C(n_377),
.Y(n_434)
);

INVx3_ASAP7_75t_SL g438 ( 
.A(n_395),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_438),
.A2(n_396),
.B1(n_401),
.B2(n_388),
.Y(n_440)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_440),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_441),
.A2(n_442),
.B(n_445),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_425),
.A2(n_397),
.B(n_389),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_420),
.A2(n_402),
.B(n_416),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_424),
.B(n_391),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_446),
.B(n_447),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_439),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_449),
.B(n_419),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_426),
.B(n_393),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_450),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_433),
.A2(n_388),
.B1(n_404),
.B2(n_398),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_452),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_453),
.B(n_4),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_418),
.B(n_410),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_455),
.B(n_457),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_417),
.B(n_404),
.C(n_379),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_456),
.B(n_458),
.C(n_428),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_434),
.B(n_136),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_422),
.B(n_136),
.C(n_101),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_474),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_448),
.A2(n_435),
.B1(n_431),
.B2(n_437),
.Y(n_463)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_463),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_452),
.B(n_430),
.C(n_418),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_465),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_456),
.B(n_427),
.C(n_438),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_445),
.A2(n_436),
.B1(n_419),
.B2(n_136),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_466),
.B(n_473),
.Y(n_478)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_467),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_SL g469 ( 
.A1(n_447),
.A2(n_101),
.B1(n_73),
.B2(n_29),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_469),
.B(n_471),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_443),
.A2(n_101),
.B(n_54),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_444),
.B(n_85),
.C(n_21),
.Y(n_473)
);

BUFx24_ASAP7_75t_SL g475 ( 
.A(n_442),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_475),
.B(n_454),
.C(n_6),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_462),
.B(n_453),
.C(n_455),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_476),
.B(n_483),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_472),
.A2(n_458),
.B(n_449),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_470),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_484),
.A2(n_473),
.B1(n_474),
.B2(n_11),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_485),
.B(n_486),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_464),
.B(n_454),
.C(n_7),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g487 ( 
.A1(n_459),
.A2(n_5),
.B(n_7),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_487),
.B(n_488),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_465),
.B(n_7),
.C(n_8),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_460),
.B(n_15),
.C(n_9),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_489),
.B(n_463),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_477),
.B(n_468),
.Y(n_491)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_491),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_496),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_461),
.C(n_467),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_493),
.B(n_497),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_481),
.B(n_8),
.C(n_10),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_486),
.B(n_478),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_498),
.B(n_499),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_488),
.B(n_8),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_493),
.B(n_480),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_503),
.B(n_504),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_490),
.A2(n_482),
.B(n_489),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_498),
.B(n_479),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_506),
.A2(n_479),
.B(n_495),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_501),
.B(n_497),
.C(n_494),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_507),
.B(n_509),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_505),
.Y(n_509)
);

FAx1_ASAP7_75t_SL g511 ( 
.A(n_510),
.B(n_505),
.CI(n_500),
.CON(n_511),
.SN(n_511)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_511),
.B(n_512),
.Y(n_513)
);

AO21x1_ASAP7_75t_L g514 ( 
.A1(n_513),
.A2(n_508),
.B(n_511),
.Y(n_514)
);

OAI321xp33_ASAP7_75t_L g515 ( 
.A1(n_514),
.A2(n_502),
.A3(n_11),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_14),
.C(n_10),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_11),
.Y(n_517)
);


endmodule