module fake_jpeg_1757_n_369 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_369);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_369;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_5),
.B(n_6),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_55),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_56),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_58),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_53),
.B(n_8),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_59),
.B(n_65),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_63),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_7),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_66),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_67),
.B(n_77),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_32),
.B(n_11),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_68),
.B(n_71),
.Y(n_125)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_70),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_1),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_72),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_73),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_2),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_74),
.B(n_80),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_2),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_78),
.Y(n_182)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_21),
.Y(n_79)
);

CKINVDCx12_ASAP7_75t_R g135 ( 
.A(n_79),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_22),
.B(n_41),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_36),
.Y(n_82)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_43),
.A2(n_2),
.B(n_4),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_83),
.A2(n_77),
.B(n_65),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_31),
.B(n_12),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_84),
.B(n_90),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_44),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_91),
.Y(n_124)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_39),
.B(n_12),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_44),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_19),
.B(n_12),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_103),
.Y(n_129)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_31),
.B(n_14),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_97),
.B(n_98),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_41),
.B(n_14),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_17),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_99),
.B(n_109),
.Y(n_151)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_100),
.Y(n_164)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_102),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_45),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_40),
.B(n_17),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_105),
.B(n_107),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_106),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_47),
.Y(n_107)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_47),
.B(n_17),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_20),
.Y(n_110)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_51),
.B(n_0),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_112),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_51),
.B(n_20),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_35),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_121),
.B(n_161),
.Y(n_203)
);

OA22x2_ASAP7_75t_L g127 ( 
.A1(n_82),
.A2(n_35),
.B1(n_26),
.B2(n_28),
.Y(n_127)
);

AO22x1_ASAP7_75t_SL g222 ( 
.A1(n_127),
.A2(n_160),
.B1(n_131),
.B2(n_115),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_60),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_128),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_65),
.A2(n_30),
.B1(n_37),
.B2(n_52),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_130),
.A2(n_167),
.B1(n_153),
.B2(n_151),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_93),
.B(n_37),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_132),
.B(n_143),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_64),
.A2(n_24),
.B1(n_52),
.B2(n_50),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_24),
.B1(n_50),
.B2(n_99),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_98),
.A2(n_109),
.B1(n_90),
.B2(n_102),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_108),
.A2(n_72),
.B1(n_55),
.B2(n_58),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_141),
.A2(n_154),
.B1(n_170),
.B2(n_180),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_112),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_66),
.C(n_73),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_150),
.B(n_160),
.C(n_142),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_88),
.A2(n_87),
.B1(n_75),
.B2(n_101),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_169),
.Y(n_186)
);

OA22x2_ASAP7_75t_L g160 ( 
.A1(n_69),
.A2(n_75),
.B1(n_55),
.B2(n_56),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_94),
.B(n_77),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_67),
.A2(n_85),
.B1(n_91),
.B2(n_83),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_81),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_82),
.A2(n_23),
.B1(n_95),
.B2(n_96),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_59),
.B(n_103),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_172),
.B(n_173),
.Y(n_224)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_60),
.Y(n_173)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_173),
.Y(n_227)
);

BUFx16f_ASAP7_75t_L g178 ( 
.A(n_55),
.Y(n_178)
);

INVx6_ASAP7_75t_SL g213 ( 
.A(n_178),
.Y(n_213)
);

CKINVDCx12_ASAP7_75t_R g179 ( 
.A(n_79),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_179),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_83),
.A2(n_74),
.B1(n_68),
.B2(n_71),
.Y(n_180)
);

AOI21xp33_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_160),
.B(n_115),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_161),
.A2(n_123),
.B1(n_155),
.B2(n_159),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_183),
.Y(n_267)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_149),
.B(n_148),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_185),
.B(n_188),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_187),
.A2(n_194),
.B1(n_202),
.B2(n_228),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_129),
.B(n_168),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_124),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_189),
.B(n_190),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_121),
.A2(n_122),
.B(n_140),
.C(n_125),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_138),
.B(n_175),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_198),
.Y(n_241)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_133),
.B1(n_118),
.B2(n_127),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

AND2x2_ASAP7_75t_SL g262 ( 
.A(n_197),
.B(n_207),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_120),
.B(n_163),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_200),
.B(n_211),
.Y(n_242)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_139),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_116),
.A2(n_162),
.B1(n_119),
.B2(n_166),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_144),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_204),
.B(n_215),
.Y(n_259)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_145),
.B(n_127),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_210),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_117),
.B(n_158),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_144),
.B(n_177),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_208),
.Y(n_264)
);

NOR3xp33_ASAP7_75t_SL g249 ( 
.A(n_209),
.B(n_203),
.C(n_199),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_164),
.B(n_119),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_152),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_128),
.A2(n_141),
.B(n_170),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_237),
.C(n_233),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_152),
.B(n_114),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_216),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_135),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_114),
.B(n_165),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g217 ( 
.A(n_156),
.B(n_171),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_218),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_146),
.B(n_182),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_131),
.B(n_134),
.Y(n_219)
);

NAND2x1_ASAP7_75t_SL g265 ( 
.A(n_219),
.B(n_222),
.Y(n_265)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_166),
.Y(n_220)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_134),
.Y(n_221)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_162),
.B(n_147),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_229),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_235),
.Y(n_258)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_126),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_113),
.A2(n_180),
.B1(n_137),
.B2(n_181),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_113),
.A2(n_126),
.B(n_167),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_176),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_180),
.A2(n_181),
.B1(n_136),
.B2(n_133),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_231),
.A2(n_196),
.B1(n_225),
.B2(n_206),
.Y(n_243)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_155),
.Y(n_232)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_160),
.Y(n_233)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_233),
.Y(n_261)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_178),
.Y(n_234)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_234),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_143),
.B(n_129),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_143),
.B(n_129),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_191),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_125),
.B(n_180),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_155),
.Y(n_238)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_240),
.B(n_251),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_243),
.A2(n_207),
.B1(n_195),
.B2(n_219),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_229),
.A2(n_187),
.B1(n_237),
.B2(n_231),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_257),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_213),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_212),
.A2(n_222),
.B1(n_223),
.B2(n_210),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_203),
.A2(n_197),
.B1(n_202),
.B2(n_222),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_186),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_258),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_263),
.B(n_268),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_198),
.B(n_191),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_191),
.B(n_193),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_269),
.B(n_205),
.Y(n_286)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_270),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_272),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_243),
.A2(n_238),
.B1(n_232),
.B2(n_184),
.Y(n_273)
);

AOI22x1_ASAP7_75t_L g307 ( 
.A1(n_273),
.A2(n_275),
.B1(n_288),
.B2(n_289),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_239),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_277),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_251),
.A2(n_230),
.B1(n_217),
.B2(n_208),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_276),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_259),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_279),
.B(n_285),
.Y(n_317)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_253),
.Y(n_280)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_280),
.Y(n_314)
);

O2A1O1Ixp33_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_190),
.B(n_213),
.C(n_226),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_281),
.B(n_287),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_208),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_284),
.C(n_264),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_286),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_207),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_191),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_253),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_244),
.A2(n_245),
.B1(n_262),
.B2(n_247),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_244),
.A2(n_201),
.B1(n_219),
.B2(n_221),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_290),
.B(n_294),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_252),
.B(n_227),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_295),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_240),
.A2(n_234),
.B(n_227),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_293),
.A2(n_265),
.B(n_267),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_245),
.A2(n_246),
.B1(n_261),
.B2(n_257),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_266),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_249),
.B(n_242),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_283),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_297),
.B(n_303),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_274),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_299),
.B(n_316),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_273),
.Y(n_302)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_302),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_255),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_305),
.A2(n_315),
.B(n_296),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_278),
.A2(n_265),
.B1(n_267),
.B2(n_256),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_275),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_311),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_241),
.C(n_266),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_293),
.A2(n_291),
.B(n_278),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_281),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_318),
.A2(n_330),
.B1(n_333),
.B2(n_313),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_307),
.A2(n_291),
.B1(n_294),
.B2(n_288),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_319),
.A2(n_322),
.B1(n_309),
.B2(n_302),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_298),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_324),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_307),
.A2(n_284),
.B1(n_272),
.B2(n_280),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_314),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_325),
.B(n_326),
.Y(n_339)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_300),
.Y(n_326)
);

OAI32xp33_ASAP7_75t_L g327 ( 
.A1(n_307),
.A2(n_295),
.A3(n_287),
.B1(n_290),
.B2(n_271),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_327),
.A2(n_331),
.B(n_305),
.Y(n_342)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_300),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_239),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_250),
.Y(n_337)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_313),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_334),
.Y(n_348)
);

A2O1A1Ixp33_ASAP7_75t_SL g335 ( 
.A1(n_321),
.A2(n_316),
.B(n_306),
.C(n_308),
.Y(n_335)
);

OA22x2_ASAP7_75t_L g346 ( 
.A1(n_335),
.A2(n_321),
.B1(n_329),
.B2(n_308),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_337),
.B(n_338),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_323),
.B(n_311),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_320),
.A2(n_317),
.B1(n_304),
.B2(n_301),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_341),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_322),
.B(n_315),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_342),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_310),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_343),
.B(n_345),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_344),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_331),
.B(n_297),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_346),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_335),
.A2(n_318),
.B1(n_309),
.B2(n_327),
.Y(n_350)
);

INVxp33_ASAP7_75t_L g356 ( 
.A(n_350),
.Y(n_356)
);

XNOR2x1_ASAP7_75t_L g354 ( 
.A(n_351),
.B(n_345),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_354),
.A2(n_353),
.B(n_347),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_349),
.B(n_301),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_355),
.B(n_358),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_352),
.B(n_336),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_352),
.B(n_339),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_359),
.B(n_312),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_357),
.Y(n_360)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_360),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_362),
.B(n_363),
.Y(n_364)
);

AOI221xp5_ASAP7_75t_L g366 ( 
.A1(n_365),
.A2(n_361),
.B1(n_350),
.B2(n_319),
.C(n_356),
.Y(n_366)
);

AO21x1_ASAP7_75t_L g367 ( 
.A1(n_366),
.A2(n_357),
.B(n_348),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_367),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_368),
.B(n_364),
.Y(n_369)
);


endmodule