module fake_jpeg_9508_n_273 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_273);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx8_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_37),
.Y(n_68)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_39),
.Y(n_64)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVxp67_ASAP7_75t_SL g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_32),
.B1(n_28),
.B2(n_17),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_49),
.B1(n_54),
.B2(n_57),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_51),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_32),
.B1(n_28),
.B2(n_17),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_33),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_32),
.B1(n_17),
.B2(n_25),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_34),
.C(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_59),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_18),
.B1(n_21),
.B2(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_33),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_63),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_33),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_35),
.A2(n_30),
.B1(n_18),
.B2(n_31),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_39),
.B1(n_35),
.B2(n_24),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_22),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_22),
.Y(n_84)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_74),
.Y(n_108)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_27),
.B1(n_23),
.B2(n_42),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_76),
.A2(n_77),
.B1(n_39),
.B2(n_64),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_35),
.B1(n_39),
.B2(n_26),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_81),
.Y(n_111)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_86),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_85),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_47),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_61),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_67),
.Y(n_101)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_96),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_56),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_SL g126 ( 
.A(n_94),
.B(n_97),
.C(n_36),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_85),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_63),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_105),
.Y(n_118)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_99),
.B(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_68),
.C(n_49),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_114),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_55),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_85),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_112),
.A2(n_90),
.B1(n_80),
.B2(n_64),
.Y(n_116)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_100),
.A2(n_78),
.B1(n_75),
.B2(n_50),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_121),
.B1(n_137),
.B2(n_112),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_116),
.A2(n_92),
.B1(n_48),
.B2(n_106),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_130),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_119),
.A2(n_125),
.B(n_126),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_120),
.B(n_127),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_78),
.B1(n_64),
.B2(n_70),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_58),
.C(n_16),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_129),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_60),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_58),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_0),
.Y(n_132)
);

NOR2x1_ASAP7_75t_SL g146 ( 
.A(n_132),
.B(n_19),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_69),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_133),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_69),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_134),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_24),
.B(n_26),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_109),
.B(n_19),
.Y(n_154)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_138),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_91),
.A2(n_89),
.B1(n_48),
.B2(n_27),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_89),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_48),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_141),
.A2(n_116),
.B1(n_128),
.B2(n_129),
.Y(n_171)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_94),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_151),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_99),
.C(n_97),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_148),
.C(n_160),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_153),
.C(n_0),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_123),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_147),
.B(n_154),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_114),
.C(n_107),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_104),
.Y(n_149)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_87),
.Y(n_150)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_87),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_157),
.Y(n_167)
);

NOR2xp67_ASAP7_75t_SL g153 ( 
.A(n_119),
.B(n_44),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_153),
.B1(n_156),
.B2(n_146),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_22),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_144),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_115),
.A2(n_92),
.B1(n_106),
.B2(n_44),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_161),
.A2(n_127),
.B1(n_135),
.B2(n_137),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_118),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_151),
.Y(n_177)
);

OAI32xp33_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_19),
.A3(n_27),
.B1(n_23),
.B2(n_22),
.Y(n_164)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_164),
.Y(n_169)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_149),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_177),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_119),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_173),
.C(n_178),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_171),
.A2(n_174),
.B1(n_181),
.B2(n_188),
.Y(n_192)
);

OAI31xp33_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_121),
.A3(n_125),
.B(n_128),
.Y(n_172)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_125),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_179),
.A2(n_29),
.B(n_2),
.Y(n_207)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_185),
.Y(n_201)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_15),
.C(n_14),
.Y(n_204)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_186),
.A2(n_189),
.B1(n_187),
.B2(n_176),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_130),
.C(n_66),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_161),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_141),
.A2(n_130),
.B1(n_29),
.B2(n_98),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_168),
.C(n_182),
.Y(n_210)
);

NOR4xp25_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_157),
.C(n_147),
.D(n_143),
.Y(n_191)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_154),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_193),
.B(n_207),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_194),
.A2(n_198),
.B(n_203),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_155),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_205),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_169),
.A2(n_140),
.B1(n_142),
.B2(n_159),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_197),
.A2(n_12),
.B1(n_62),
.B2(n_72),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_167),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_164),
.Y(n_199)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_174),
.C(n_46),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_163),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_204),
.A2(n_206),
.B(n_3),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_46),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_0),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_172),
.B1(n_182),
.B2(n_175),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_209),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_220),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_211),
.A2(n_226),
.B(n_194),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_29),
.C(n_72),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_222),
.Y(n_233)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_208),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_217),
.A2(n_221),
.B(n_203),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_36),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_201),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_1),
.C(n_2),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_1),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_190),
.Y(n_234)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_204),
.Y(n_231)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_195),
.A2(n_10),
.B(n_5),
.Y(n_226)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_216),
.Y(n_229)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_236),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_218),
.A2(n_192),
.B1(n_212),
.B2(n_214),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_235),
.A2(n_224),
.B1(n_226),
.B2(n_7),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_214),
.B(n_193),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_206),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_238),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_199),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_219),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_243),
.C(n_7),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_220),
.C(n_223),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_6),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_229),
.A2(n_232),
.B(n_228),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_247),
.A2(n_248),
.B(n_6),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_236),
.A2(n_3),
.B(n_6),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_233),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_252),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_230),
.B(n_234),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_254),
.C(n_243),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_7),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_255),
.B(n_256),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_8),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_8),
.Y(n_257)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_257),
.Y(n_258)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_260),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_257),
.B(n_241),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_249),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_266),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_249),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_258),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_259),
.C(n_258),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_269),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_264),
.B(n_268),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_271),
.A2(n_263),
.B(n_9),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_9),
.Y(n_273)
);


endmodule