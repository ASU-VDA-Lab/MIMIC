module fake_jpeg_20102_n_286 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_286);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_286;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_26),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_60),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_26),
.B1(n_21),
.B2(n_31),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_37),
.B1(n_42),
.B2(n_41),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_26),
.B1(n_21),
.B2(n_31),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_50),
.A2(n_57),
.B1(n_37),
.B2(n_42),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_22),
.C(n_29),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_21),
.B1(n_31),
.B2(n_27),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_19),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_63),
.A2(n_44),
.B(n_29),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_37),
.B1(n_38),
.B2(n_42),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_64),
.A2(n_69),
.B1(n_76),
.B2(n_80),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_65),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_37),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_67),
.A2(n_81),
.B1(n_90),
.B2(n_92),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_68),
.B(n_18),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_27),
.B1(n_41),
.B2(n_42),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_60),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_73),
.B(n_99),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_27),
.B1(n_32),
.B2(n_25),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_98),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_41),
.B1(n_40),
.B2(n_36),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_52),
.B(n_24),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_84),
.B(n_87),
.Y(n_113)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_86),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_24),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_47),
.A2(n_36),
.B1(n_40),
.B2(n_62),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_88),
.A2(n_89),
.B1(n_96),
.B2(n_101),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_47),
.A2(n_19),
.B1(n_25),
.B2(n_32),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_47),
.A2(n_34),
.B1(n_28),
.B2(n_23),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_56),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_97),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_53),
.A2(n_34),
.B1(n_28),
.B2(n_23),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_30),
.B(n_33),
.C(n_35),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_93),
.A2(n_94),
.B(n_30),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_53),
.A2(n_30),
.B1(n_33),
.B2(n_18),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_56),
.A2(n_40),
.B1(n_36),
.B2(n_35),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_46),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_40),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_61),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_61),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_100),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_48),
.A2(n_36),
.B1(n_17),
.B2(n_18),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_111),
.B(n_112),
.Y(n_146)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_29),
.C(n_44),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_128),
.Y(n_132)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_118),
.B(n_79),
.Y(n_153)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_18),
.B1(n_17),
.B2(n_30),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_126),
.A2(n_68),
.B1(n_80),
.B2(n_88),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_64),
.B1(n_63),
.B2(n_81),
.Y(n_138)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_73),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_134),
.B(n_135),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_129),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_71),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_136),
.B(n_143),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_126),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_139),
.A2(n_144),
.B1(n_150),
.B2(n_121),
.Y(n_178)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_67),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_120),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_30),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_63),
.B1(n_75),
.B2(n_78),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_153),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_72),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_148),
.B(n_152),
.Y(n_177)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_116),
.A2(n_81),
.B1(n_67),
.B2(n_94),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_103),
.Y(n_152)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_105),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_107),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_104),
.B(n_117),
.Y(n_156)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_157),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_158),
.B(n_173),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_147),
.A2(n_116),
.B1(n_119),
.B2(n_109),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_163),
.B1(n_175),
.B2(n_178),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_176),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_128),
.C(n_123),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_150),
.C(n_138),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_108),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_93),
.Y(n_193)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_146),
.Y(n_173)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_179),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_147),
.A2(n_119),
.B1(n_108),
.B2(n_124),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_106),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_145),
.A2(n_102),
.B1(n_107),
.B2(n_75),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_181),
.A2(n_155),
.B1(n_149),
.B2(n_140),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_130),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_183),
.B(n_184),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_137),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_172),
.C(n_168),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_176),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_198),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_161),
.A2(n_139),
.B1(n_144),
.B2(n_133),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_191),
.A2(n_197),
.B1(n_205),
.B2(n_208),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_193),
.B(n_33),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_196),
.B1(n_204),
.B2(n_159),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_162),
.A2(n_142),
.B1(n_137),
.B2(n_130),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_142),
.B1(n_100),
.B2(n_99),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_82),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_177),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_200),
.B(n_201),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_167),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_160),
.B(n_15),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_202),
.B(n_14),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_86),
.B(n_95),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_203),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_183),
.A2(n_85),
.B1(n_78),
.B2(n_83),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_163),
.A2(n_185),
.B1(n_167),
.B2(n_180),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_171),
.A2(n_14),
.B1(n_1),
.B2(n_2),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_179),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_210),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_187),
.A2(n_182),
.B1(n_164),
.B2(n_168),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_194),
.B1(n_204),
.B2(n_189),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_186),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_214),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_208),
.B(n_182),
.Y(n_214)
);

XNOR2x1_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_33),
.Y(n_215)
);

XNOR2x1_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_222),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_198),
.C(n_188),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_190),
.B(n_159),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_219),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_220),
.A2(n_224),
.B1(n_33),
.B2(n_20),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_195),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_223),
.B(n_227),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_172),
.B1(n_174),
.B2(n_2),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_20),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_226),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_20),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_220),
.A2(n_191),
.B(n_197),
.C(n_187),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_225),
.B(n_226),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_240),
.C(n_239),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_217),
.A2(n_203),
.B1(n_205),
.B2(n_192),
.Y(n_231)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_233),
.A2(n_224),
.B1(n_225),
.B2(n_215),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g234 ( 
.A(n_221),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_234),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_0),
.C(n_1),
.Y(n_240)
);

NAND2xp33_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_1),
.Y(n_241)
);

NAND2xp33_ASAP7_75t_SL g247 ( 
.A(n_241),
.B(n_3),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_2),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_244),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_3),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_252),
.C(n_237),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_248),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_230),
.B(n_227),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_249),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_221),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_236),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_253),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_222),
.C(n_5),
.Y(n_252)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_257),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_240),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_261),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_254),
.A2(n_234),
.B(n_235),
.Y(n_263)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_263),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_246),
.A2(n_256),
.B(n_245),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_264),
.A2(n_246),
.B(n_249),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_237),
.C(n_228),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_255),
.Y(n_272)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_267),
.Y(n_276)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_260),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_269),
.B(n_271),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_257),
.A2(n_253),
.B(n_228),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_272),
.A2(n_228),
.B1(n_7),
.B2(n_8),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_269),
.A2(n_259),
.B(n_262),
.Y(n_273)
);

AOI21xp33_ASAP7_75t_L g279 ( 
.A1(n_273),
.A2(n_266),
.B(n_10),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_277),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_4),
.B1(n_7),
.B2(n_9),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_276),
.A2(n_275),
.B(n_270),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_4),
.Y(n_282)
);

NAND2x1_ASAP7_75t_SL g281 ( 
.A(n_279),
.B(n_273),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_281),
.A2(n_282),
.B(n_280),
.Y(n_283)
);

O2A1O1Ixp33_ASAP7_75t_SL g284 ( 
.A1(n_283),
.A2(n_281),
.B(n_11),
.C(n_12),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_10),
.B(n_11),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_285),
.B(n_10),
.Y(n_286)
);


endmodule