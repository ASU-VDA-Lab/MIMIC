module fake_jpeg_11538_n_40 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_40);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_40;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_15),
.B(n_19),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_21),
.B(n_23),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_19),
.B1(n_14),
.B2(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_28),
.B1(n_0),
.B2(n_1),
.Y(n_30)
);

XOR2x2_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_6),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_0),
.C(n_1),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_17),
.B1(n_18),
.B2(n_2),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_20),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_29),
.B(n_30),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_32),
.C(n_24),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_35),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_24),
.C(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_36),
.B1(n_20),
.B2(n_10),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_3),
.Y(n_40)
);


endmodule