module fake_aes_4028_n_30 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
OAI21x1_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_4), .B(n_7), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
CKINVDCx6p67_ASAP7_75t_R g15 ( .A(n_10), .Y(n_15) );
CKINVDCx8_ASAP7_75t_R g16 ( .A(n_0), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_11), .Y(n_17) );
AND2x4_ASAP7_75t_L g18 ( .A(n_5), .B(n_0), .Y(n_18) );
AOI22xp33_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_15), .B1(n_17), .B2(n_14), .Y(n_19) );
BUFx3_ASAP7_75t_L g20 ( .A(n_14), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
OAI322xp33_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_17), .A3(n_16), .B1(n_19), .B2(n_18), .C1(n_20), .C2(n_15), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
AOI222xp33_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_18), .B1(n_20), .B2(n_13), .C1(n_16), .C2(n_5), .Y(n_25) );
OAI21xp33_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_24), .B(n_13), .Y(n_26) );
OAI22xp33_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_27) );
XNOR2x1_ASAP7_75t_SL g28 ( .A(n_27), .B(n_1), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
AOI322xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_26), .A3(n_3), .B1(n_4), .B2(n_6), .C1(n_2), .C2(n_9), .Y(n_30) );
endmodule