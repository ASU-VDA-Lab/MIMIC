module fake_jpeg_1953_n_617 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_617);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_617;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx8_ASAP7_75t_SL g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_14),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_32),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g192 ( 
.A(n_59),
.Y(n_192)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_27),
.B(n_9),
.Y(n_62)
);

NAND2x1p5_ASAP7_75t_L g179 ( 
.A(n_62),
.B(n_66),
.Y(n_179)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g137 ( 
.A(n_63),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_64),
.Y(n_156)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_65),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_27),
.B(n_9),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_67),
.Y(n_160)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_69),
.Y(n_190)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_71),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_26),
.B(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_72),
.B(n_125),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_73),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_74),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_75),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_80),
.Y(n_154)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_81),
.Y(n_186)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_82),
.Y(n_142)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_83),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_84),
.Y(n_155)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_86),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_87),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_88),
.Y(n_185)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_89),
.Y(n_176)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_93),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_94),
.Y(n_202)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_95),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_96),
.Y(n_194)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_98),
.Y(n_204)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_100),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_101),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_102),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_103),
.Y(n_215)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

BUFx16f_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_105),
.Y(n_189)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_21),
.Y(n_108)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_40),
.Y(n_109)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_109),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_23),
.Y(n_110)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_110),
.Y(n_209)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_23),
.Y(n_111)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_112),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_29),
.Y(n_114)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_114),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_115),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_33),
.Y(n_116)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_116),
.Y(n_213)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_20),
.Y(n_117)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_33),
.Y(n_118)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_33),
.Y(n_119)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_34),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_127),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_33),
.Y(n_121)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_121),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_33),
.Y(n_122)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_122),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_123),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_50),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_124),
.Y(n_195)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_36),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_126),
.B(n_53),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_21),
.Y(n_127)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_50),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_24),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_62),
.A2(n_56),
.B1(n_55),
.B2(n_37),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_129),
.A2(n_150),
.B1(n_162),
.B2(n_167),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_80),
.A2(n_46),
.B1(n_52),
.B2(n_47),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_143),
.A2(n_147),
.B1(n_168),
.B2(n_173),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_145),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_69),
.A2(n_46),
.B1(n_52),
.B2(n_47),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_66),
.A2(n_43),
.B1(n_55),
.B2(n_28),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_76),
.B(n_56),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_161),
.B(n_163),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_61),
.A2(n_37),
.B1(n_43),
.B2(n_28),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_49),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_164),
.B(n_0),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_64),
.A2(n_49),
.B1(n_45),
.B2(n_53),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_107),
.A2(n_45),
.B1(n_21),
.B2(n_30),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_105),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_171),
.B(n_183),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_90),
.A2(n_93),
.B1(n_104),
.B2(n_99),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_63),
.A2(n_21),
.B1(n_30),
.B2(n_24),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_175),
.A2(n_184),
.B1(n_219),
.B2(n_41),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_123),
.B(n_25),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_71),
.A2(n_21),
.B1(n_25),
.B2(n_39),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_124),
.B(n_11),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_187),
.B(n_198),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_108),
.B(n_11),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_114),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_201),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_116),
.B(n_12),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_73),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_206),
.B1(n_214),
.B2(n_122),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_74),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_118),
.B(n_13),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_208),
.B(n_218),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_67),
.A2(n_41),
.B1(n_39),
.B2(n_20),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_119),
.B(n_12),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_101),
.A2(n_41),
.B1(n_39),
.B2(n_34),
.Y(n_219)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_130),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_220),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_221),
.Y(n_350)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_132),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_222),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_192),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_223),
.B(n_235),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_224),
.A2(n_251),
.B1(n_280),
.B2(n_281),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_137),
.Y(n_226)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_226),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

BUFx4f_ASAP7_75t_L g311 ( 
.A(n_227),
.Y(n_311)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_137),
.Y(n_228)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_228),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_154),
.Y(n_229)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_229),
.Y(n_300)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_230),
.Y(n_302)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_151),
.Y(n_231)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_231),
.Y(n_304)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_157),
.Y(n_232)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_232),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_179),
.B(n_121),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_233),
.B(n_263),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_188),
.Y(n_235)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_130),
.Y(n_236)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_236),
.Y(n_322)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_165),
.Y(n_237)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_237),
.Y(n_324)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_169),
.Y(n_238)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_238),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_239),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_172),
.B(n_109),
.C(n_100),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_240),
.B(n_279),
.C(n_184),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_205),
.A2(n_98),
.B1(n_96),
.B2(n_88),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_241),
.A2(n_211),
.B1(n_160),
.B2(n_158),
.Y(n_338)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_177),
.Y(n_242)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_242),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_243),
.Y(n_308)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_141),
.Y(n_245)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_245),
.Y(n_333)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_141),
.Y(n_246)
);

INVx4_ASAP7_75t_SL g335 ( 
.A(n_246),
.Y(n_335)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_178),
.Y(n_247)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_247),
.Y(n_348)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_193),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_248),
.Y(n_330)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_191),
.Y(n_249)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_249),
.Y(n_351)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_196),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_250),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_154),
.A2(n_87),
.B1(n_84),
.B2(n_78),
.Y(n_251)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_203),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_253),
.B(n_255),
.Y(n_319)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_213),
.Y(n_255)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_186),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_257),
.B(n_259),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_148),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_258),
.Y(n_346)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_139),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_179),
.A2(n_77),
.B1(n_75),
.B2(n_34),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_260),
.A2(n_264),
.B1(n_270),
.B2(n_272),
.Y(n_305)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_186),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_261),
.B(n_262),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_140),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_133),
.B(n_10),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_136),
.A2(n_42),
.B1(n_10),
.B2(n_12),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_138),
.B(n_8),
.Y(n_265)
);

NOR3xp33_ASAP7_75t_L g327 ( 
.A(n_265),
.B(n_271),
.C(n_276),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_148),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_266),
.B(n_268),
.Y(n_331)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_159),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_159),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_269),
.B(n_273),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_206),
.A2(n_42),
.B1(n_8),
.B2(n_13),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_193),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_147),
.A2(n_219),
.B1(n_143),
.B2(n_168),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_166),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_135),
.A2(n_42),
.B1(n_7),
.B2(n_13),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_274),
.A2(n_277),
.B1(n_283),
.B2(n_289),
.Y(n_326)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_152),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_275),
.B(n_278),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_165),
.A2(n_42),
.B1(n_13),
.B2(n_5),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_174),
.B(n_170),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_146),
.B(n_142),
.C(n_210),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_176),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_135),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_149),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_282),
.A2(n_286),
.B1(n_288),
.B2(n_292),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_149),
.A2(n_42),
.B1(n_15),
.B2(n_6),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_189),
.B(n_6),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_284),
.B(n_287),
.Y(n_341)
);

A2O1A1Ixp33_ASAP7_75t_L g285 ( 
.A1(n_181),
.A2(n_6),
.B(n_7),
.C(n_15),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_285),
.A2(n_209),
.B(n_199),
.Y(n_321)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_182),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_188),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_156),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_155),
.A2(n_6),
.B1(n_15),
.B2(n_16),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_195),
.B(n_15),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_290),
.B(n_291),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_131),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_217),
.Y(n_292)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_217),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_294),
.A2(n_296),
.B1(n_131),
.B2(n_215),
.Y(n_320)
);

AO22x2_ASAP7_75t_SL g295 ( 
.A1(n_197),
.A2(n_1),
.B1(n_4),
.B2(n_17),
.Y(n_295)
);

OA22x2_ASAP7_75t_L g314 ( 
.A1(n_295),
.A2(n_194),
.B1(n_204),
.B2(n_185),
.Y(n_314)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_156),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_234),
.A2(n_243),
.B(n_175),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_298),
.A2(n_347),
.B(n_248),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_301),
.B(n_349),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_240),
.B(n_144),
.C(n_207),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_309),
.B(n_310),
.C(n_334),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_279),
.B(n_144),
.C(n_153),
.Y(n_310)
);

NAND2xp33_ASAP7_75t_SL g312 ( 
.A(n_276),
.B(n_209),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_312),
.A2(n_321),
.B(n_340),
.Y(n_368)
);

OAI22xp33_ASAP7_75t_L g313 ( 
.A1(n_234),
.A2(n_173),
.B1(n_204),
.B2(n_155),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_313),
.A2(n_336),
.B1(n_345),
.B2(n_326),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_314),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_320),
.Y(n_375)
);

AOI32xp33_ASAP7_75t_L g328 ( 
.A1(n_252),
.A2(n_180),
.A3(n_199),
.B1(n_202),
.B2(n_134),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_328),
.B(n_237),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_244),
.B(n_180),
.C(n_197),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_256),
.A2(n_158),
.B1(n_185),
.B2(n_194),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_338),
.A2(n_297),
.B1(n_301),
.B2(n_326),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_225),
.A2(n_211),
.B(n_160),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_L g345 ( 
.A1(n_256),
.A2(n_17),
.B1(n_251),
.B2(n_295),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_285),
.A2(n_17),
.B(n_278),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_231),
.B(n_17),
.C(n_238),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_349),
.B(n_352),
.C(n_347),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_267),
.B(n_254),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_241),
.A2(n_257),
.B1(n_261),
.B2(n_286),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_353),
.A2(n_226),
.B1(n_229),
.B2(n_275),
.Y(n_355)
);

OAI32xp33_ASAP7_75t_L g354 ( 
.A1(n_293),
.A2(n_295),
.A3(n_250),
.B1(n_255),
.B2(n_253),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_354),
.B(n_277),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_355),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_321),
.A2(n_264),
.B(n_246),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_356),
.A2(n_360),
.B(n_397),
.Y(n_410)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_311),
.Y(n_357)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_357),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_358),
.B(n_391),
.Y(n_415)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_311),
.Y(n_359)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_359),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_308),
.A2(n_294),
.B1(n_292),
.B2(n_271),
.Y(n_360)
);

OAI21xp33_ASAP7_75t_L g421 ( 
.A1(n_362),
.A2(n_372),
.B(n_330),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_339),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_363),
.B(n_364),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_329),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_299),
.B(n_245),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_365),
.B(n_385),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_298),
.A2(n_282),
.B1(n_281),
.B2(n_296),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_366),
.A2(n_377),
.B1(n_382),
.B2(n_386),
.Y(n_406)
);

XOR2x2_ASAP7_75t_SL g367 ( 
.A(n_341),
.B(n_344),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_367),
.B(n_385),
.Y(n_423)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_311),
.Y(n_369)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_369),
.Y(n_403)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_324),
.Y(n_370)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_370),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_340),
.B(n_268),
.Y(n_371)
);

CKINVDCx14_ASAP7_75t_R g419 ( 
.A(n_371),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_SL g373 ( 
.A(n_344),
.B(n_273),
.C(n_269),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_373),
.B(n_384),
.C(n_389),
.Y(n_411)
);

AOI22x1_ASAP7_75t_L g374 ( 
.A1(n_308),
.A2(n_220),
.B1(n_236),
.B2(n_288),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_374),
.A2(n_396),
.B1(n_335),
.B2(n_324),
.Y(n_408)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_319),
.Y(n_376)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_376),
.Y(n_428)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_319),
.Y(n_378)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_378),
.Y(n_435)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_319),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_379),
.B(n_380),
.Y(n_418)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_307),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_325),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_381),
.B(n_387),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_338),
.A2(n_354),
.B1(n_305),
.B2(n_336),
.Y(n_382)
);

XNOR2x1_ASAP7_75t_L g407 ( 
.A(n_383),
.B(n_395),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_309),
.B(n_310),
.C(n_334),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_299),
.B(n_352),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_303),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_307),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_388),
.B(n_392),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_341),
.B(n_316),
.C(n_342),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_323),
.B(n_312),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_315),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_393),
.B(n_394),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_305),
.A2(n_314),
.B1(n_323),
.B2(n_328),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_314),
.A2(n_327),
.B1(n_317),
.B2(n_322),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_331),
.A2(n_351),
.B(n_302),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_314),
.A2(n_302),
.B1(n_348),
.B2(n_318),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_398),
.B(n_343),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_350),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_399),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_358),
.A2(n_322),
.B1(n_348),
.B2(n_318),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_405),
.A2(n_398),
.B1(n_382),
.B2(n_428),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_L g450 ( 
.A1(n_408),
.A2(n_390),
.B1(n_396),
.B2(n_379),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_362),
.A2(n_332),
.B(n_300),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_409),
.A2(n_425),
.B(n_431),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_395),
.B(n_351),
.C(n_346),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_412),
.B(n_413),
.C(n_416),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_361),
.B(n_346),
.C(n_333),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_361),
.B(n_304),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_414),
.B(n_371),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_384),
.B(n_333),
.C(n_306),
.Y(n_416)
);

OAI21xp33_ASAP7_75t_L g459 ( 
.A1(n_421),
.A2(n_378),
.B(n_375),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_423),
.B(n_373),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_365),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_424),
.B(n_429),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_368),
.A2(n_300),
.B(n_325),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_367),
.B(n_306),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_427),
.B(n_436),
.C(n_397),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_363),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_368),
.A2(n_343),
.B(n_350),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_433),
.B(n_376),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_389),
.B(n_311),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_434),
.B(n_337),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_383),
.B(n_330),
.C(n_304),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_437),
.B(n_448),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_419),
.A2(n_371),
.B(n_356),
.Y(n_438)
);

AO21x1_ASAP7_75t_L g496 ( 
.A1(n_438),
.A2(n_447),
.B(n_465),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_417),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_439),
.B(n_445),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_405),
.A2(n_394),
.B1(n_377),
.B2(n_371),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_442),
.A2(n_450),
.B1(n_451),
.B2(n_462),
.Y(n_475)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_417),
.Y(n_443)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_443),
.Y(n_481)
);

CKINVDCx14_ASAP7_75t_R g487 ( 
.A(n_444),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_402),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_418),
.Y(n_446)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_446),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_419),
.A2(n_371),
.B(n_391),
.Y(n_447)
);

OA22x2_ASAP7_75t_L g448 ( 
.A1(n_406),
.A2(n_390),
.B1(n_374),
.B2(n_386),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_449),
.B(n_456),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_426),
.A2(n_366),
.B1(n_387),
.B2(n_364),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_402),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_453),
.B(n_467),
.Y(n_484)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_418),
.Y(n_454)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_454),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_407),
.B(n_414),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_455),
.B(n_463),
.C(n_416),
.Y(n_477)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_430),
.Y(n_457)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_457),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_414),
.Y(n_474)
);

OAI211xp5_ASAP7_75t_L g489 ( 
.A1(n_459),
.A2(n_447),
.B(n_445),
.C(n_453),
.Y(n_489)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_430),
.Y(n_460)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_460),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_433),
.Y(n_461)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_461),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_SL g462 ( 
.A1(n_400),
.A2(n_399),
.B1(n_370),
.B2(n_381),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_407),
.B(n_388),
.C(n_380),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_406),
.A2(n_360),
.B1(n_374),
.B2(n_393),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_464),
.A2(n_468),
.B1(n_408),
.B2(n_428),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_410),
.A2(n_392),
.B(n_357),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_424),
.B(n_359),
.Y(n_466)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_466),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_429),
.B(n_369),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_415),
.A2(n_337),
.B1(n_335),
.B2(n_350),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_469),
.B(n_470),
.Y(n_500)
);

FAx1_ASAP7_75t_SL g470 ( 
.A(n_423),
.B(n_335),
.CI(n_337),
.CON(n_470),
.SN(n_470)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_474),
.B(n_449),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_442),
.A2(n_426),
.B1(n_415),
.B2(n_410),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_476),
.A2(n_479),
.B1(n_491),
.B2(n_457),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_477),
.B(n_497),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_438),
.A2(n_431),
.B(n_427),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g518 ( 
.A(n_478),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_437),
.A2(n_425),
.B1(n_409),
.B2(n_434),
.Y(n_479)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_482),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_452),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_483),
.B(n_492),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_446),
.B(n_404),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_488),
.B(n_493),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_489),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_461),
.A2(n_411),
.B1(n_435),
.B2(n_404),
.Y(n_491)
);

AOI32xp33_ASAP7_75t_L g492 ( 
.A1(n_452),
.A2(n_411),
.A3(n_435),
.B1(n_413),
.B2(n_422),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_467),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_455),
.B(n_412),
.C(n_436),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_498),
.C(n_458),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_463),
.B(n_420),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_440),
.B(n_422),
.C(n_420),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_440),
.B(n_401),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_501),
.B(n_469),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_SL g502 ( 
.A(n_471),
.B(n_456),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_502),
.B(n_512),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_506),
.B(n_516),
.C(n_523),
.Y(n_534)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_480),
.Y(n_507)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_507),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_508),
.A2(n_515),
.B1(n_517),
.B2(n_482),
.Y(n_531)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_480),
.Y(n_509)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_509),
.Y(n_539)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_484),
.Y(n_510)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_510),
.Y(n_545)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_484),
.Y(n_511)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_511),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_471),
.B(n_454),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_513),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_497),
.B(n_460),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_514),
.B(n_521),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_475),
.A2(n_439),
.B1(n_444),
.B2(n_464),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_501),
.B(n_443),
.C(n_465),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_475),
.A2(n_472),
.B1(n_479),
.B2(n_476),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_487),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_473),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_522),
.B(n_524),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_477),
.B(n_466),
.C(n_441),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_SL g524 ( 
.A(n_474),
.B(n_451),
.Y(n_524)
);

FAx1_ASAP7_75t_SL g525 ( 
.A(n_498),
.B(n_470),
.CI(n_441),
.CON(n_525),
.SN(n_525)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_525),
.B(n_478),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_526),
.B(n_527),
.C(n_491),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_494),
.B(n_468),
.C(n_470),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_496),
.Y(n_528)
);

CKINVDCx14_ASAP7_75t_R g538 ( 
.A(n_528),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_530),
.B(n_536),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_531),
.A2(n_504),
.B1(n_517),
.B2(n_526),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_510),
.B(n_473),
.Y(n_533)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_533),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_520),
.B(n_485),
.C(n_486),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_537),
.B(n_547),
.C(n_523),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_511),
.B(n_490),
.Y(n_541)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_541),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_518),
.A2(n_472),
.B1(n_500),
.B2(n_499),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_542),
.A2(n_546),
.B1(n_548),
.B2(n_515),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_503),
.B(n_486),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_543),
.B(n_516),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_505),
.A2(n_472),
.B1(n_499),
.B2(n_485),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_520),
.B(n_481),
.C(n_495),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_504),
.A2(n_495),
.B1(n_496),
.B2(n_448),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_550),
.B(n_555),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_538),
.A2(n_508),
.B(n_519),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_551),
.A2(n_559),
.B(n_448),
.Y(n_581)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_552),
.Y(n_569)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_553),
.Y(n_573)
);

CKINVDCx16_ASAP7_75t_R g555 ( 
.A(n_532),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_540),
.B(n_527),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_556),
.B(n_561),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_534),
.B(n_506),
.C(n_524),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_557),
.B(n_564),
.C(n_536),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_530),
.A2(n_549),
.B(n_545),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_537),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_560),
.B(n_563),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_540),
.B(n_514),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_562),
.A2(n_535),
.B1(n_529),
.B2(n_548),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_543),
.B(n_525),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_534),
.B(n_512),
.C(n_513),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_533),
.B(n_525),
.Y(n_566)
);

AOI21x1_ASAP7_75t_L g578 ( 
.A1(n_566),
.A2(n_544),
.B(n_535),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_554),
.B(n_547),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_567),
.B(n_572),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_561),
.B(n_531),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_568),
.B(n_552),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_570),
.B(n_564),
.C(n_556),
.Y(n_585)
);

NOR2xp67_ASAP7_75t_L g571 ( 
.A(n_553),
.B(n_541),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_L g591 ( 
.A1(n_571),
.A2(n_578),
.B(n_575),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_554),
.B(n_539),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_550),
.B(n_563),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_574),
.B(n_566),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_559),
.A2(n_546),
.B1(n_542),
.B2(n_551),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_577),
.A2(n_579),
.B1(n_448),
.B2(n_403),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_581),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_568),
.B(n_557),
.C(n_562),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_582),
.B(n_584),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_585),
.B(n_588),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_587),
.B(n_575),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_570),
.B(n_558),
.C(n_565),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_580),
.B(n_565),
.Y(n_589)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_589),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_590),
.Y(n_597)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_591),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_576),
.B(n_502),
.C(n_448),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_592),
.B(n_586),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_573),
.B(n_401),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_593),
.A2(n_578),
.B(n_581),
.Y(n_599)
);

OAI21x1_ASAP7_75t_L g603 ( 
.A1(n_594),
.A2(n_599),
.B(n_601),
.Y(n_603)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_598),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_583),
.B(n_569),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_600),
.B(n_588),
.Y(n_604)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_604),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_595),
.B(n_582),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_605),
.B(n_607),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_596),
.B(n_602),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_594),
.A2(n_587),
.B(n_579),
.Y(n_608)
);

AOI21x1_ASAP7_75t_SL g610 ( 
.A1(n_608),
.A2(n_601),
.B(n_577),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_SL g612 ( 
.A1(n_610),
.A2(n_603),
.B(n_606),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_SL g614 ( 
.A1(n_612),
.A2(n_613),
.B(n_611),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_609),
.B(n_597),
.C(n_576),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_614),
.A2(n_592),
.B(n_403),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_615),
.B(n_432),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g617 ( 
.A(n_616),
.B(n_432),
.Y(n_617)
);


endmodule