module real_aes_1895_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_756;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_0), .B(n_121), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_1), .A2(n_130), .B(n_135), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_2), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_3), .B(n_137), .Y(n_176) );
INVx1_ASAP7_75t_L g128 ( .A(n_4), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_5), .B(n_137), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_6), .B(n_148), .Y(n_510) );
INVx1_ASAP7_75t_L g530 ( .A(n_7), .Y(n_530) );
CKINVDCx16_ASAP7_75t_R g457 ( .A(n_8), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_9), .Y(n_543) );
NAND2xp33_ASAP7_75t_L g199 ( .A(n_10), .B(n_139), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_11), .A2(n_37), .B1(n_432), .B2(n_433), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_11), .Y(n_433) );
INVx2_ASAP7_75t_L g118 ( .A(n_12), .Y(n_118) );
AOI221x1_ASAP7_75t_L g223 ( .A1(n_13), .A2(n_27), .B1(n_121), .B2(n_130), .C(n_224), .Y(n_223) );
CKINVDCx16_ASAP7_75t_R g444 ( .A(n_14), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_15), .B(n_121), .Y(n_195) );
AO21x2_ASAP7_75t_L g192 ( .A1(n_16), .A2(n_193), .B(n_194), .Y(n_192) );
INVx1_ASAP7_75t_L g519 ( .A(n_17), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_18), .B(n_141), .Y(n_227) );
XOR2xp5_ASAP7_75t_L g472 ( .A(n_19), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_20), .B(n_137), .Y(n_152) );
AO21x1_ASAP7_75t_L g171 ( .A1(n_21), .A2(n_121), .B(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g448 ( .A(n_22), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_23), .A2(n_59), .B1(n_474), .B2(n_475), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g475 ( .A(n_23), .Y(n_475) );
INVx1_ASAP7_75t_L g517 ( .A(n_24), .Y(n_517) );
INVx1_ASAP7_75t_SL g584 ( .A(n_25), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_26), .B(n_122), .Y(n_504) );
NAND2x1_ASAP7_75t_L g216 ( .A(n_28), .B(n_137), .Y(n_216) );
AOI33xp33_ASAP7_75t_L g562 ( .A1(n_29), .A2(n_55), .A3(n_492), .B1(n_501), .B2(n_563), .B3(n_564), .Y(n_562) );
NAND2x1_ASAP7_75t_L g162 ( .A(n_30), .B(n_139), .Y(n_162) );
INVx1_ASAP7_75t_L g538 ( .A(n_31), .Y(n_538) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_32), .A2(n_90), .B(n_118), .Y(n_117) );
OR2x2_ASAP7_75t_L g143 ( .A(n_32), .B(n_90), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_33), .B(n_528), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_34), .B(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_35), .B(n_137), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_36), .B(n_139), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_37), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_38), .A2(n_130), .B(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g127 ( .A(n_39), .B(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g131 ( .A(n_39), .B(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g500 ( .A(n_39), .Y(n_500) );
OR2x6_ASAP7_75t_L g446 ( .A(n_40), .B(n_447), .Y(n_446) );
AOI221xp5_ASAP7_75t_L g103 ( .A1(n_41), .A2(n_104), .B1(n_452), .B2(n_459), .C(n_468), .Y(n_103) );
OAI22xp5_ASAP7_75t_SL g434 ( .A1(n_41), .A2(n_89), .B1(n_435), .B2(n_436), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_41), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_42), .B(n_831), .Y(n_830) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_43), .B(n_121), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_44), .B(n_528), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_45), .A2(n_116), .B1(n_148), .B2(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_46), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_47), .B(n_122), .Y(n_585) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_48), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_49), .B(n_139), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_50), .B(n_193), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_51), .B(n_122), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_52), .A2(n_130), .B(n_161), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_53), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_54), .B(n_139), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_56), .B(n_122), .Y(n_555) );
INVx1_ASAP7_75t_L g124 ( .A(n_57), .Y(n_124) );
INVx1_ASAP7_75t_L g134 ( .A(n_57), .Y(n_134) );
AND2x2_ASAP7_75t_L g556 ( .A(n_58), .B(n_141), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_59), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g527 ( .A1(n_60), .A2(n_76), .B1(n_498), .B2(n_528), .C(n_529), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_61), .B(n_528), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_62), .B(n_137), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_63), .B(n_116), .Y(n_545) );
AOI21xp5_ASAP7_75t_SL g573 ( .A1(n_64), .A2(n_498), .B(n_574), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_65), .A2(n_130), .B(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g513 ( .A(n_66), .Y(n_513) );
AO21x1_ASAP7_75t_L g173 ( .A1(n_67), .A2(n_130), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g120 ( .A(n_68), .B(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g554 ( .A(n_69), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_70), .B(n_121), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_71), .A2(n_498), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g188 ( .A(n_72), .B(n_142), .Y(n_188) );
INVx1_ASAP7_75t_L g126 ( .A(n_73), .Y(n_126) );
INVx1_ASAP7_75t_L g132 ( .A(n_73), .Y(n_132) );
AND2x2_ASAP7_75t_L g166 ( .A(n_74), .B(n_115), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_75), .B(n_528), .Y(n_565) );
AND2x2_ASAP7_75t_L g586 ( .A(n_77), .B(n_115), .Y(n_586) );
INVx1_ASAP7_75t_L g514 ( .A(n_78), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_79), .A2(n_498), .B(n_583), .Y(n_582) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_80), .A2(n_498), .B(n_503), .C(n_508), .Y(n_497) );
OAI22xp5_ASAP7_75t_SL g470 ( .A1(n_81), .A2(n_471), .B1(n_472), .B2(n_476), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_81), .Y(n_476) );
INVx1_ASAP7_75t_L g449 ( .A(n_82), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_83), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g114 ( .A(n_84), .B(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_85), .B(n_121), .Y(n_154) );
AND2x2_ASAP7_75t_SL g571 ( .A(n_86), .B(n_115), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_87), .A2(n_498), .B1(n_560), .B2(n_561), .Y(n_559) );
AND2x2_ASAP7_75t_L g172 ( .A(n_88), .B(n_148), .Y(n_172) );
CKINVDCx16_ASAP7_75t_R g436 ( .A(n_89), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_91), .B(n_139), .Y(n_153) );
AND2x2_ASAP7_75t_L g219 ( .A(n_92), .B(n_115), .Y(n_219) );
INVx1_ASAP7_75t_L g575 ( .A(n_93), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_94), .B(n_137), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_95), .A2(n_130), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_96), .B(n_139), .Y(n_225) );
AND2x2_ASAP7_75t_L g566 ( .A(n_97), .B(n_115), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_98), .B(n_137), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_99), .A2(n_536), .B(n_537), .C(n_539), .Y(n_535) );
BUFx2_ASAP7_75t_L g458 ( .A(n_100), .Y(n_458) );
BUFx2_ASAP7_75t_SL g465 ( .A(n_100), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_101), .A2(n_130), .B(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_102), .B(n_122), .Y(n_576) );
OAI21x1_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_439), .B(n_450), .Y(n_104) );
AOI22xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_434), .B1(n_437), .B2(n_438), .Y(n_105) );
INVx2_ASAP7_75t_L g437 ( .A(n_106), .Y(n_437) );
XNOR2x1_ASAP7_75t_L g106 ( .A(n_107), .B(n_431), .Y(n_106) );
INVx2_ASAP7_75t_L g829 ( .A(n_107), .Y(n_829) );
AND2x4_ASAP7_75t_L g107 ( .A(n_108), .B(n_316), .Y(n_107) );
NOR3xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_271), .C(n_300), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g109 ( .A(n_110), .B(n_244), .Y(n_109) );
AOI221xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_167), .B1(n_189), .B2(n_201), .C(n_205), .Y(n_110) );
INVx3_ASAP7_75t_SL g361 ( .A(n_111), .Y(n_361) );
AND2x2_ASAP7_75t_SL g111 ( .A(n_112), .B(n_144), .Y(n_111) );
NAND2x1p5_ASAP7_75t_L g207 ( .A(n_112), .B(n_157), .Y(n_207) );
INVx4_ASAP7_75t_L g242 ( .A(n_112), .Y(n_242) );
AND2x2_ASAP7_75t_L g264 ( .A(n_112), .B(n_158), .Y(n_264) );
AND2x2_ASAP7_75t_L g270 ( .A(n_112), .B(n_209), .Y(n_270) );
INVx5_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g239 ( .A(n_113), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_113), .B(n_157), .Y(n_315) );
AND2x2_ASAP7_75t_L g320 ( .A(n_113), .B(n_158), .Y(n_320) );
AND2x2_ASAP7_75t_L g332 ( .A(n_113), .B(n_192), .Y(n_332) );
NOR2x1_ASAP7_75t_SL g371 ( .A(n_113), .B(n_209), .Y(n_371) );
OR2x6_ASAP7_75t_L g113 ( .A(n_114), .B(n_119), .Y(n_113) );
INVx3_ASAP7_75t_L g187 ( .A(n_115), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_115), .A2(n_187), .B1(n_435), .B2(n_535), .Y(n_534) );
INVx4_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_116), .B(n_542), .Y(n_541) );
INVx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx4f_ASAP7_75t_L g193 ( .A(n_117), .Y(n_193) );
AND2x2_ASAP7_75t_SL g142 ( .A(n_118), .B(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g148 ( .A(n_118), .B(n_143), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_129), .B(n_141), .Y(n_119) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_127), .Y(n_121) );
INVx1_ASAP7_75t_L g515 ( .A(n_122), .Y(n_515) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_125), .Y(n_122) );
AND2x6_ASAP7_75t_L g139 ( .A(n_123), .B(n_132), .Y(n_139) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x4_ASAP7_75t_L g137 ( .A(n_125), .B(n_134), .Y(n_137) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx5_ASAP7_75t_L g140 ( .A(n_127), .Y(n_140) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_127), .Y(n_539) );
AND2x2_ASAP7_75t_L g133 ( .A(n_128), .B(n_134), .Y(n_133) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_128), .Y(n_493) );
AND2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
BUFx3_ASAP7_75t_L g495 ( .A(n_131), .Y(n_495) );
INVx2_ASAP7_75t_L g502 ( .A(n_132), .Y(n_502) );
AND2x4_ASAP7_75t_L g498 ( .A(n_133), .B(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g492 ( .A(n_134), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_138), .B(n_140), .Y(n_135) );
INVxp67_ASAP7_75t_L g520 ( .A(n_137), .Y(n_520) );
INVxp67_ASAP7_75t_L g518 ( .A(n_139), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_140), .A2(n_152), .B(n_153), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_140), .A2(n_162), .B(n_163), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_140), .A2(n_175), .B(n_176), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_140), .A2(n_184), .B(n_185), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_140), .A2(n_198), .B(n_199), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_140), .A2(n_216), .B(n_217), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_140), .A2(n_225), .B(n_226), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_140), .A2(n_504), .B(n_505), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_140), .B(n_148), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_SL g529 ( .A1(n_140), .A2(n_507), .B(n_530), .C(n_531), .Y(n_529) );
O2A1O1Ixp33_ASAP7_75t_L g553 ( .A1(n_140), .A2(n_507), .B(n_554), .C(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g560 ( .A(n_140), .Y(n_560) );
O2A1O1Ixp33_ASAP7_75t_L g574 ( .A1(n_140), .A2(n_507), .B(n_575), .C(n_576), .Y(n_574) );
O2A1O1Ixp33_ASAP7_75t_SL g583 ( .A1(n_140), .A2(n_507), .B(n_584), .C(n_585), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_141), .Y(n_165) );
OA21x2_ASAP7_75t_L g222 ( .A1(n_141), .A2(n_223), .B(n_227), .Y(n_222) );
OA21x2_ASAP7_75t_L g267 ( .A1(n_141), .A2(n_223), .B(n_227), .Y(n_267) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g200 ( .A(n_144), .Y(n_200) );
AND2x2_ASAP7_75t_L g304 ( .A(n_144), .B(n_253), .Y(n_304) );
AND2x2_ASAP7_75t_L g401 ( .A(n_144), .B(n_332), .Y(n_401) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_157), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g233 ( .A(n_146), .Y(n_233) );
INVx2_ASAP7_75t_L g255 ( .A(n_146), .Y(n_255) );
AO21x2_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_149), .B(n_155), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_147), .B(n_156), .Y(n_155) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_147), .A2(n_149), .B(n_155), .Y(n_209) );
INVx1_ASAP7_75t_SL g147 ( .A(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_148), .B(n_178), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_148), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_148), .A2(n_573), .B(n_577), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_154), .Y(n_149) );
AND2x2_ASAP7_75t_L g230 ( .A(n_157), .B(n_191), .Y(n_230) );
INVx2_ASAP7_75t_L g234 ( .A(n_157), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_157), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g333 ( .A(n_157), .B(n_298), .Y(n_333) );
OR2x2_ASAP7_75t_L g380 ( .A(n_157), .B(n_192), .Y(n_380) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_158), .Y(n_330) );
AO21x2_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_165), .B(n_166), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_164), .Y(n_159) );
AO21x2_ASAP7_75t_L g579 ( .A1(n_165), .A2(n_580), .B(n_586), .Y(n_579) );
AND2x2_ASAP7_75t_L g377 ( .A(n_167), .B(n_258), .Y(n_377) );
AND2x2_ASAP7_75t_L g427 ( .A(n_167), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OR2x2_ASAP7_75t_L g303 ( .A(n_168), .B(n_247), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_169), .B(n_179), .Y(n_168) );
AND2x2_ASAP7_75t_L g236 ( .A(n_169), .B(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g266 ( .A(n_169), .B(n_267), .Y(n_266) );
AND2x4_ASAP7_75t_L g287 ( .A(n_169), .B(n_267), .Y(n_287) );
AND2x4_ASAP7_75t_L g322 ( .A(n_169), .B(n_310), .Y(n_322) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g203 ( .A(n_170), .Y(n_203) );
OAI21x1_ASAP7_75t_SL g170 ( .A1(n_171), .A2(n_173), .B(n_177), .Y(n_170) );
INVx1_ASAP7_75t_L g178 ( .A(n_172), .Y(n_178) );
AND2x2_ASAP7_75t_L g249 ( .A(n_179), .B(n_202), .Y(n_249) );
AND2x2_ASAP7_75t_L g335 ( .A(n_179), .B(n_267), .Y(n_335) );
AND2x2_ASAP7_75t_L g346 ( .A(n_179), .B(n_211), .Y(n_346) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g210 ( .A(n_180), .B(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g277 ( .A(n_180), .B(n_212), .Y(n_277) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_187), .B(n_188), .Y(n_180) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_181), .A2(n_187), .B(n_188), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_182), .B(n_186), .Y(n_181) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_187), .A2(n_213), .B(n_219), .Y(n_212) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_187), .A2(n_213), .B(n_219), .Y(n_237) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_187), .A2(n_550), .B(n_556), .Y(n_549) );
AO21x2_ASAP7_75t_L g603 ( .A1(n_187), .A2(n_550), .B(n_556), .Y(n_603) );
INVx2_ASAP7_75t_SL g189 ( .A(n_190), .Y(n_189) );
OR2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_200), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_191), .B(n_242), .Y(n_299) );
AND2x2_ASAP7_75t_L g343 ( .A(n_191), .B(n_209), .Y(n_343) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_192), .B(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g253 ( .A(n_192), .Y(n_253) );
BUFx3_ASAP7_75t_L g262 ( .A(n_192), .Y(n_262) );
AND2x2_ASAP7_75t_L g285 ( .A(n_192), .B(n_255), .Y(n_285) );
INVx2_ASAP7_75t_SL g508 ( .A(n_193), .Y(n_508) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_193), .A2(n_527), .B(n_532), .Y(n_526) );
OAI322xp33_ASAP7_75t_L g205 ( .A1(n_200), .A2(n_206), .A3(n_210), .B1(n_220), .B2(n_228), .C1(n_235), .C2(n_240), .Y(n_205) );
INVx1_ASAP7_75t_L g366 ( .A(n_200), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_201), .B(n_241), .Y(n_240) );
AND2x4_ASAP7_75t_L g279 ( .A(n_201), .B(n_221), .Y(n_279) );
INVx2_ASAP7_75t_L g324 ( .A(n_201), .Y(n_324) );
AND2x2_ASAP7_75t_L g340 ( .A(n_201), .B(n_282), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_201), .B(n_358), .Y(n_388) );
AND2x4_ASAP7_75t_L g201 ( .A(n_202), .B(n_204), .Y(n_201) );
AND2x2_ASAP7_75t_SL g291 ( .A(n_202), .B(n_267), .Y(n_291) );
OR2x2_ASAP7_75t_L g312 ( .A(n_202), .B(n_229), .Y(n_312) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
BUFx2_ASAP7_75t_L g284 ( .A(n_203), .Y(n_284) );
INVx2_ASAP7_75t_L g229 ( .A(n_204), .Y(n_229) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_204), .Y(n_231) );
OR2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
INVx2_ASAP7_75t_L g274 ( .A(n_207), .Y(n_274) );
INVxp67_ASAP7_75t_SL g294 ( .A(n_208), .Y(n_294) );
INVx1_ASAP7_75t_L g392 ( .A(n_208), .Y(n_392) );
INVxp67_ASAP7_75t_SL g407 ( .A(n_208), .Y(n_407) );
NAND2x1_ASAP7_75t_L g417 ( .A(n_210), .B(n_221), .Y(n_417) );
INVx1_ASAP7_75t_L g424 ( .A(n_210), .Y(n_424) );
BUFx2_ASAP7_75t_L g258 ( .A(n_211), .Y(n_258) );
AND2x2_ASAP7_75t_L g334 ( .A(n_211), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
BUFx3_ASAP7_75t_L g243 ( .A(n_212), .Y(n_243) );
INVxp67_ASAP7_75t_L g247 ( .A(n_212), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_218), .Y(n_213) );
NAND3xp33_ASAP7_75t_L g235 ( .A(n_220), .B(n_236), .C(n_238), .Y(n_235) );
INVx1_ASAP7_75t_SL g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_SL g256 ( .A(n_221), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_221), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g408 ( .A(n_221), .B(n_357), .Y(n_408) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g310 ( .A(n_222), .Y(n_310) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_222), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B1(n_231), .B2(n_232), .Y(n_228) );
AND2x4_ASAP7_75t_SL g357 ( .A(n_229), .B(n_237), .Y(n_357) );
AND2x2_ASAP7_75t_L g370 ( .A(n_230), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_231), .Y(n_372) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
INVx2_ASAP7_75t_L g329 ( .A(n_233), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_233), .B(n_242), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_234), .B(n_252), .Y(n_251) );
AND3x2_ASAP7_75t_L g269 ( .A(n_234), .B(n_262), .C(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g293 ( .A(n_234), .Y(n_293) );
AND2x2_ASAP7_75t_L g406 ( .A(n_234), .B(n_407), .Y(n_406) );
BUFx2_ASAP7_75t_L g282 ( .A(n_237), .Y(n_282) );
INVx1_ASAP7_75t_L g360 ( .A(n_237), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_238), .B(n_261), .Y(n_399) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_239), .B(n_343), .Y(n_348) );
AND2x4_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
AND2x2_ASAP7_75t_L g339 ( .A(n_242), .B(n_285), .Y(n_339) );
INVx1_ASAP7_75t_SL g290 ( .A(n_243), .Y(n_290) );
AND2x2_ASAP7_75t_L g398 ( .A(n_243), .B(n_310), .Y(n_398) );
AND2x2_ASAP7_75t_L g419 ( .A(n_243), .B(n_291), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_250), .B1(n_256), .B2(n_259), .C(n_265), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
INVx1_ASAP7_75t_L g411 ( .A(n_247), .Y(n_411) );
AOI21xp33_ASAP7_75t_SL g265 ( .A1(n_248), .A2(n_266), .B(n_268), .Y(n_265) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g257 ( .A(n_249), .B(n_258), .Y(n_257) );
AOI222xp33_ASAP7_75t_L g280 ( .A1(n_249), .A2(n_281), .B1(n_283), .B2(n_288), .C1(n_292), .C2(n_295), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_249), .B(n_398), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g301 ( .A1(n_250), .A2(n_279), .B1(n_302), .B2(n_304), .Y(n_301) );
INVx1_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
INVx1_ASAP7_75t_L g286 ( .A(n_253), .Y(n_286) );
AND2x2_ASAP7_75t_L g405 ( .A(n_253), .B(n_371), .Y(n_405) );
OAI32xp33_ASAP7_75t_L g409 ( .A1(n_253), .A2(n_278), .A3(n_330), .B1(n_338), .B2(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g414 ( .A(n_253), .B(n_264), .Y(n_414) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g298 ( .A(n_255), .Y(n_298) );
OAI21xp5_ASAP7_75t_SL g305 ( .A1(n_256), .A2(n_306), .B(n_313), .Y(n_305) );
INVx1_ASAP7_75t_L g369 ( .A(n_258), .Y(n_369) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
AND2x2_ASAP7_75t_L g273 ( .A(n_261), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx2_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g281 ( .A(n_264), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g354 ( .A(n_264), .B(n_285), .Y(n_354) );
INVx1_ASAP7_75t_SL g425 ( .A(n_266), .Y(n_425) );
AND2x2_ASAP7_75t_L g359 ( .A(n_267), .B(n_360), .Y(n_359) );
OAI222xp33_ASAP7_75t_L g412 ( .A1(n_268), .A2(n_321), .B1(n_400), .B2(n_413), .C1(n_415), .C2(n_417), .Y(n_412) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g385 ( .A(n_270), .B(n_386), .Y(n_385) );
OAI21xp33_ASAP7_75t_SL g271 ( .A1(n_272), .A2(n_275), .B(n_280), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_274), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
INVx1_ASAP7_75t_L g353 ( .A(n_276), .Y(n_353) );
INVx1_ASAP7_75t_L g321 ( .A(n_277), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_277), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g375 ( .A(n_282), .Y(n_375) );
AO22x1_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B1(n_286), .B2(n_287), .Y(n_283) );
OAI322xp33_ASAP7_75t_L g395 ( .A1(n_284), .A2(n_345), .A3(n_348), .B1(n_396), .B2(n_397), .C1(n_399), .C2(n_400), .Y(n_395) );
AND2x2_ASAP7_75t_SL g319 ( .A(n_285), .B(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g314 ( .A(n_286), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_287), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g416 ( .A(n_287), .B(n_346), .Y(n_416) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g396 ( .A(n_290), .Y(n_396) );
INVx1_ASAP7_75t_SL g325 ( .A(n_291), .Y(n_325) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
OR2x2_ASAP7_75t_L g327 ( .A(n_299), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g365 ( .A(n_299), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_305), .Y(n_300) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_311), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g338 ( .A(n_309), .B(n_324), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_309), .B(n_346), .Y(n_345) );
BUFx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g368 ( .A(n_312), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NOR2x1_ASAP7_75t_L g316 ( .A(n_317), .B(n_381), .Y(n_316) );
NAND4xp25_ASAP7_75t_L g317 ( .A(n_318), .B(n_336), .C(n_349), .D(n_362), .Y(n_317) );
AOI322xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_321), .A3(n_322), .B1(n_323), .B2(n_326), .C1(n_331), .C2(n_334), .Y(n_318) );
AOI211xp5_ASAP7_75t_L g418 ( .A1(n_319), .A2(n_419), .B(n_420), .C(n_423), .Y(n_418) );
AND2x2_ASAP7_75t_L g430 ( .A(n_320), .B(n_407), .Y(n_430) );
INVx1_ASAP7_75t_L g352 ( .A(n_322), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_322), .B(n_357), .Y(n_394) );
NAND2xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_330), .B(n_343), .Y(n_410) );
AND2x4_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
AOI222xp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_339), .B1(n_340), .B2(n_341), .C1(n_344), .C2(n_347), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g349 ( .A1(n_339), .A2(n_350), .B1(n_353), .B2(n_354), .C(n_355), .Y(n_349) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AOI21xp33_ASAP7_75t_SL g355 ( .A1(n_356), .A2(n_358), .B(n_361), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_367), .B1(n_370), .B2(n_372), .C(n_373), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g422 ( .A(n_371), .Y(n_422) );
AOI21xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_376), .B(n_378), .Y(n_373) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx2_ASAP7_75t_L g386 ( .A(n_380), .Y(n_386) );
OR2x2_ASAP7_75t_L g421 ( .A(n_380), .B(n_422), .Y(n_421) );
NAND3xp33_ASAP7_75t_L g381 ( .A(n_382), .B(n_402), .C(n_418), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_395), .Y(n_382) );
OAI21xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_387), .B(n_389), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_393), .Y(n_389) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_408), .B1(n_409), .B2(n_411), .C(n_412), .Y(n_402) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NOR2x1_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_417), .B(n_421), .Y(n_420) );
O2A1O1Ixp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B(n_426), .C(n_429), .Y(n_423) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g438 ( .A(n_434), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVxp67_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx2_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_443), .Y(n_451) );
BUFx2_ASAP7_75t_L g467 ( .A(n_443), .Y(n_467) );
BUFx2_ASAP7_75t_L g838 ( .A(n_443), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
CKINVDCx16_ASAP7_75t_R g826 ( .A(n_444), .Y(n_826) );
OR2x2_ASAP7_75t_L g832 ( .A(n_444), .B(n_446), .Y(n_832) );
O2A1O1Ixp33_ASAP7_75t_SL g468 ( .A1(n_445), .A2(n_469), .B(n_830), .C(n_833), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
CKINVDCx9p33_ASAP7_75t_R g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_SL g455 ( .A(n_456), .B(n_458), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_456), .A2(n_463), .B(n_466), .Y(n_462) );
INVx2_ASAP7_75t_L g837 ( .A(n_456), .Y(n_837) );
NAND2xp5_ASAP7_75t_SL g836 ( .A(n_458), .B(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
CKINVDCx11_ASAP7_75t_R g463 ( .A(n_464), .Y(n_463) );
CKINVDCx8_ASAP7_75t_R g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
XNOR2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_477), .Y(n_469) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp33_ASAP7_75t_SL g477 ( .A(n_478), .B(n_827), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_826), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_760), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_482), .B(n_683), .Y(n_481) );
NAND3xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_630), .C(n_663), .Y(n_482) );
AOI211xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_587), .B(n_596), .C(n_620), .Y(n_483) );
OAI21xp33_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_522), .B(n_567), .Y(n_484) );
OR2x2_ASAP7_75t_L g640 ( .A(n_485), .B(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g795 ( .A(n_485), .B(n_796), .Y(n_795) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AOI22xp33_ASAP7_75t_SL g685 ( .A1(n_486), .A2(n_686), .B1(n_690), .B2(n_692), .Y(n_685) );
AND2x2_ASAP7_75t_L g722 ( .A(n_486), .B(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_509), .Y(n_486) );
INVx1_ASAP7_75t_L g619 ( .A(n_487), .Y(n_619) );
AND2x4_ASAP7_75t_L g636 ( .A(n_487), .B(n_617), .Y(n_636) );
INVx2_ASAP7_75t_L g658 ( .A(n_487), .Y(n_658) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_487), .Y(n_741) );
AND2x2_ASAP7_75t_L g812 ( .A(n_487), .B(n_570), .Y(n_812) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_497), .Y(n_487) );
NOR3xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_494), .C(n_496), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x4_ASAP7_75t_L g528 ( .A(n_491), .B(n_495), .Y(n_528) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
OR2x6_ASAP7_75t_L g507 ( .A(n_492), .B(n_502), .Y(n_507) );
INVxp33_ASAP7_75t_L g563 ( .A(n_492), .Y(n_563) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVxp67_ASAP7_75t_L g544 ( .A(n_498), .Y(n_544) );
NOR2x1p5_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g564 ( .A(n_501), .Y(n_564) );
INVx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_507), .A2(n_513), .B1(n_514), .B2(n_515), .Y(n_512) );
INVxp67_ASAP7_75t_L g536 ( .A(n_507), .Y(n_536) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_508), .A2(n_558), .B(n_566), .Y(n_557) );
AO21x2_ASAP7_75t_L g601 ( .A1(n_508), .A2(n_558), .B(n_566), .Y(n_601) );
AND2x2_ASAP7_75t_L g578 ( .A(n_509), .B(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g606 ( .A(n_509), .Y(n_606) );
INVx3_ASAP7_75t_L g617 ( .A(n_509), .Y(n_617) );
AND2x4_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
OAI21xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_516), .B(n_521), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_515), .B(n_538), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B1(n_519), .B2(n_520), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g806 ( .A1(n_522), .A2(n_807), .B1(n_809), .B2(n_811), .Y(n_806) );
NAND2xp5_ASAP7_75t_SL g817 ( .A(n_522), .B(n_818), .Y(n_817) );
INVx2_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_547), .Y(n_523) );
INVx3_ASAP7_75t_L g590 ( .A(n_524), .Y(n_590) );
AND2x2_ASAP7_75t_L g598 ( .A(n_524), .B(n_599), .Y(n_598) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_524), .Y(n_628) );
NAND2x1_ASAP7_75t_SL g822 ( .A(n_524), .B(n_589), .Y(n_822) );
AND2x4_ASAP7_75t_L g524 ( .A(n_525), .B(n_533), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g595 ( .A(n_526), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_526), .B(n_601), .Y(n_613) );
AND2x2_ASAP7_75t_L g626 ( .A(n_526), .B(n_533), .Y(n_626) );
AND2x4_ASAP7_75t_L g633 ( .A(n_526), .B(n_634), .Y(n_633) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_526), .Y(n_682) );
INVxp67_ASAP7_75t_L g689 ( .A(n_526), .Y(n_689) );
INVx1_ASAP7_75t_L g694 ( .A(n_526), .Y(n_694) );
INVx1_ASAP7_75t_L g546 ( .A(n_528), .Y(n_546) );
INVx1_ASAP7_75t_L g593 ( .A(n_533), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_533), .B(n_603), .Y(n_612) );
INVx2_ASAP7_75t_L g680 ( .A(n_533), .Y(n_680) );
INVx1_ASAP7_75t_L g719 ( .A(n_533), .Y(n_719) );
OR2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_540), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_544), .B1(n_545), .B2(n_546), .Y(n_540) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g649 ( .A(n_547), .B(n_626), .Y(n_649) );
AND2x2_ASAP7_75t_L g717 ( .A(n_547), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g731 ( .A(n_547), .B(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_547), .B(n_746), .Y(n_745) );
AND2x4_ASAP7_75t_L g547 ( .A(n_548), .B(n_557), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NOR2x1_ASAP7_75t_L g594 ( .A(n_549), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g687 ( .A(n_549), .B(n_680), .Y(n_687) );
AND2x2_ASAP7_75t_L g778 ( .A(n_549), .B(n_600), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g589 ( .A(n_557), .Y(n_589) );
INVx2_ASAP7_75t_L g634 ( .A(n_557), .Y(n_634) );
AND2x2_ASAP7_75t_L g679 ( .A(n_557), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_559), .B(n_565), .Y(n_558) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_578), .Y(n_568) );
AND2x2_ASAP7_75t_L g721 ( .A(n_569), .B(n_722), .Y(n_721) );
OR2x6_ASAP7_75t_L g780 ( .A(n_569), .B(n_781), .Y(n_780) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx4_ASAP7_75t_L g610 ( .A(n_570), .Y(n_610) );
AND2x4_ASAP7_75t_L g618 ( .A(n_570), .B(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g653 ( .A(n_570), .B(n_579), .Y(n_653) );
INVx2_ASAP7_75t_L g702 ( .A(n_570), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g751 ( .A(n_570), .B(n_676), .Y(n_751) );
AND2x2_ASAP7_75t_L g788 ( .A(n_570), .B(n_606), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_570), .B(n_671), .Y(n_796) );
OR2x6_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
AND2x2_ASAP7_75t_L g629 ( .A(n_578), .B(n_618), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_578), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_SL g768 ( .A(n_578), .B(n_656), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_578), .B(n_669), .Y(n_790) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_579), .Y(n_608) );
AND2x2_ASAP7_75t_L g616 ( .A(n_579), .B(n_617), .Y(n_616) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_579), .Y(n_639) );
INVx2_ASAP7_75t_L g642 ( .A(n_579), .Y(n_642) );
INVx1_ASAP7_75t_L g675 ( .A(n_579), .Y(n_675) );
INVx1_ASAP7_75t_L g723 ( .A(n_579), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
NAND2xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_591), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_589), .B(n_592), .Y(n_665) );
OR2x2_ASAP7_75t_L g737 ( .A(n_589), .B(n_738), .Y(n_737) );
AND4x1_ASAP7_75t_SL g783 ( .A(n_589), .B(n_765), .C(n_784), .D(n_785), .Y(n_783) );
OR2x2_ASAP7_75t_L g807 ( .A(n_590), .B(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g644 ( .A(n_593), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_593), .B(n_602), .Y(n_794) );
AND2x2_ASAP7_75t_L g819 ( .A(n_594), .B(n_679), .Y(n_819) );
OAI32xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_604), .A3(n_609), .B1(n_611), .B2(n_614), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g692 ( .A(n_599), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g792 ( .A(n_599), .B(n_746), .Y(n_792) );
AND2x4_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
AND2x2_ASAP7_75t_L g688 ( .A(n_600), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g774 ( .A(n_600), .Y(n_774) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_601), .B(n_603), .Y(n_808) );
INVx3_ASAP7_75t_L g625 ( .A(n_602), .Y(n_625) );
NAND2x1p5_ASAP7_75t_L g803 ( .A(n_602), .B(n_730), .Y(n_803) );
INVx3_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_603), .Y(n_662) );
AND2x2_ASAP7_75t_L g681 ( .A(n_603), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g815 ( .A(n_605), .Y(n_815) );
NAND2x1_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_L g655 ( .A(n_606), .Y(n_655) );
NOR2x1_ASAP7_75t_L g756 ( .A(n_606), .B(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_609), .B(n_715), .Y(n_714) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g647 ( .A(n_610), .B(n_615), .Y(n_647) );
AND2x4_ASAP7_75t_L g669 ( .A(n_610), .B(n_619), .Y(n_669) );
AND2x4_ASAP7_75t_SL g740 ( .A(n_610), .B(n_741), .Y(n_740) );
NOR2x1_ASAP7_75t_L g766 ( .A(n_610), .B(n_691), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_611), .A2(n_734), .B1(n_737), .B2(n_739), .Y(n_733) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx2_ASAP7_75t_SL g753 ( .A(n_612), .Y(n_753) );
INVx2_ASAP7_75t_L g645 ( .A(n_613), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_618), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_616), .B(n_622), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_616), .A2(n_752), .B1(n_755), .B2(n_758), .Y(n_754) );
INVx1_ASAP7_75t_L g676 ( .A(n_617), .Y(n_676) );
AND2x2_ASAP7_75t_L g699 ( .A(n_617), .B(n_658), .Y(n_699) );
INVx2_ASAP7_75t_L g622 ( .A(n_618), .Y(n_622) );
OAI21xp5_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_623), .B(n_627), .Y(n_620) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_624), .A2(n_696), .B1(n_700), .B2(n_701), .Y(n_695) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_625), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_625), .B(n_693), .Y(n_709) );
INVx1_ASAP7_75t_L g713 ( .A(n_625), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
NOR3xp33_ASAP7_75t_L g630 ( .A(n_631), .B(n_646), .C(n_650), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_635), .B1(n_640), .B2(n_643), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g660 ( .A(n_633), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g700 ( .A(n_633), .B(n_687), .Y(n_700) );
AND2x2_ASAP7_75t_L g752 ( .A(n_633), .B(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g769 ( .A(n_633), .B(n_719), .Y(n_769) );
AND2x2_ASAP7_75t_L g824 ( .A(n_633), .B(n_718), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx4_ASAP7_75t_L g691 ( .A(n_636), .Y(n_691) );
AND2x2_ASAP7_75t_L g701 ( .A(n_636), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
BUFx2_ASAP7_75t_L g706 ( .A(n_639), .Y(n_706) );
AND2x2_ASAP7_75t_L g715 ( .A(n_639), .B(n_699), .Y(n_715) );
INVx1_ASAP7_75t_L g750 ( .A(n_641), .Y(n_750) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g671 ( .A(n_642), .Y(n_671) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_644), .B(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_645), .B(n_713), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_654), .B(n_659), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_652), .B(n_691), .Y(n_800) );
INVx2_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
AOI21xp33_ASAP7_75t_SL g663 ( .A1(n_655), .A2(n_664), .B(n_666), .Y(n_663) );
AND2x2_ASAP7_75t_L g810 ( .A(n_655), .B(n_669), .Y(n_810) );
AND2x4_ASAP7_75t_L g673 ( .A(n_656), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_SL g707 ( .A(n_656), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g789 ( .A(n_656), .B(n_723), .Y(n_789) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AOI21xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_672), .B(n_677), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_669), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_669), .B(n_674), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_670), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g732 ( .A(n_670), .Y(n_732) );
INVx1_ASAP7_75t_L g736 ( .A(n_670), .Y(n_736) );
AND2x2_ASAP7_75t_L g820 ( .A(n_670), .B(n_788), .Y(n_820) );
AND2x2_ASAP7_75t_L g823 ( .A(n_670), .B(n_740), .Y(n_823) );
INVx3_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AND2x4_ASAP7_75t_SL g674 ( .A(n_675), .B(n_676), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_675), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x4_ASAP7_75t_L g678 ( .A(n_679), .B(n_681), .Y(n_678) );
INVx1_ASAP7_75t_L g802 ( .A(n_679), .Y(n_802) );
AND2x2_ASAP7_75t_L g693 ( .A(n_680), .B(n_694), .Y(n_693) );
NAND4xp75_ASAP7_75t_L g683 ( .A(n_684), .B(n_703), .C(n_724), .D(n_742), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_695), .Y(n_684) );
AND2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
NAND2x1p5_ASAP7_75t_L g773 ( .A(n_687), .B(n_774), .Y(n_773) );
NAND2x1p5_ASAP7_75t_L g759 ( .A(n_688), .B(n_753), .Y(n_759) );
NAND2xp5_ASAP7_75t_R g775 ( .A(n_691), .B(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g825 ( .A(n_691), .Y(n_825) );
INVx2_ASAP7_75t_L g738 ( .A(n_693), .Y(n_738) );
BUFx3_ASAP7_75t_L g730 ( .A(n_694), .Y(n_730) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
BUFx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g781 ( .A(n_699), .Y(n_781) );
AND2x2_ASAP7_75t_L g735 ( .A(n_701), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g757 ( .A(n_702), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_708), .B(n_710), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_706), .B(n_740), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_707), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_709), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_714), .B1(n_716), .B2(n_720), .Y(n_710) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
OA21x2_ASAP7_75t_L g725 ( .A1(n_718), .A2(n_726), .B(n_727), .Y(n_725) );
INVx1_ASAP7_75t_L g746 ( .A(n_718), .Y(n_746) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g777 ( .A(n_719), .B(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g785 ( .A(n_719), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_720), .B(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g755 ( .A(n_723), .B(n_756), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_731), .B(n_733), .Y(n_724) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OR2x2_ASAP7_75t_L g772 ( .A(n_729), .B(n_773), .Y(n_772) );
INVx3_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_736), .Y(n_784) );
INVx2_ASAP7_75t_SL g776 ( .A(n_740), .Y(n_776) );
AND2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_754), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_747), .B1(n_749), .B2(n_752), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g805 ( .A(n_749), .Y(n_805) );
NOR2x1_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx3_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_761), .B(n_797), .Y(n_760) );
NAND3xp33_ASAP7_75t_L g761 ( .A(n_762), .B(n_770), .C(n_782), .Y(n_761) );
NOR2x1_ASAP7_75t_L g762 ( .A(n_763), .B(n_767), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
BUFx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
AND2x2_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
AOI22xp33_ASAP7_75t_SL g770 ( .A1(n_771), .A2(n_775), .B1(n_777), .B2(n_779), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
NOR3xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_786), .C(n_793), .Y(n_782) );
AOI21xp33_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_790), .B(n_791), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_798), .B(n_816), .Y(n_797) );
NOR3xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_806), .C(n_813), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_801), .B1(n_804), .B2(n_805), .Y(n_799) );
OR2x2_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
NOR3xp33_ASAP7_75t_L g813 ( .A(n_807), .B(n_812), .C(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVxp67_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
AOI222xp33_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_820), .B1(n_821), .B2(n_823), .C1(n_824), .C2(n_825), .Y(n_816) );
INVx1_ASAP7_75t_SL g818 ( .A(n_819), .Y(n_818) );
INVx2_ASAP7_75t_SL g821 ( .A(n_822), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_826), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_828), .B(n_829), .Y(n_827) );
INVx3_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx2_ASAP7_75t_SL g833 ( .A(n_834), .Y(n_833) );
AND2x2_ASAP7_75t_L g834 ( .A(n_835), .B(n_838), .Y(n_834) );
INVxp67_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
endmodule