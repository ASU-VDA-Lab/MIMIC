module fake_jpeg_21807_n_248 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx24_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_29),
.B(n_31),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_7),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_35),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_7),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_23),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_26),
.B1(n_23),
.B2(n_24),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_32),
.A2(n_26),
.B1(n_23),
.B2(n_24),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_48)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_24),
.B1(n_26),
.B2(n_21),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_29),
.B(n_14),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_35),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_21),
.B1(n_20),
.B2(n_22),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_33),
.B1(n_27),
.B2(n_19),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_22),
.B1(n_20),
.B2(n_19),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_56),
.A2(n_37),
.B1(n_15),
.B2(n_28),
.Y(n_60)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_58),
.Y(n_81)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_70),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_64),
.B1(n_67),
.B2(n_51),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_33),
.B1(n_22),
.B2(n_20),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_15),
.B1(n_22),
.B2(n_28),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_33),
.B1(n_14),
.B2(n_27),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_33),
.B(n_13),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_40),
.B(n_46),
.C(n_47),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_56),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_71),
.B(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_31),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_91),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_85),
.B1(n_86),
.B2(n_93),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_80),
.A2(n_82),
.B(n_84),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_40),
.B(n_45),
.C(n_48),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_39),
.C(n_55),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_52),
.B1(n_50),
.B2(n_38),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_49),
.B(n_53),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_64),
.B(n_9),
.Y(n_118)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_65),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_61),
.B(n_18),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_63),
.A2(n_52),
.B1(n_50),
.B2(n_38),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_42),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_18),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_95),
.B(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_62),
.B(n_1),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_97),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_101),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_92),
.B(n_71),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_103),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_76),
.B1(n_59),
.B2(n_58),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_112),
.B1(n_114),
.B2(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_107),
.Y(n_127)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_106),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_75),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_116),
.Y(n_134)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_110),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_57),
.B1(n_64),
.B2(n_73),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_83),
.B(n_64),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_113),
.A2(n_82),
.B(n_78),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_79),
.A2(n_64),
.B1(n_73),
.B2(n_74),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_95),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_118),
.A2(n_87),
.B(n_80),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_115),
.A2(n_83),
.B(n_84),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_131),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_100),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_125),
.B(n_110),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_138),
.B1(n_112),
.B2(n_114),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_115),
.B(n_85),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_130),
.Y(n_145)
);

AOI32xp33_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_80),
.A3(n_82),
.B1(n_91),
.B2(n_96),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_135),
.Y(n_153)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_140),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_133),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_149),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_111),
.C(n_104),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_156),
.C(n_122),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_172)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_152),
.B(n_119),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_155),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_104),
.C(n_108),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_99),
.B1(n_107),
.B2(n_113),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_124),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_131),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_126),
.A2(n_139),
.B1(n_136),
.B2(n_130),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_138),
.A2(n_113),
.B1(n_78),
.B2(n_101),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_151),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_167),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_105),
.C(n_100),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_137),
.B1(n_121),
.B2(n_135),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_166),
.A2(n_160),
.B1(n_148),
.B2(n_150),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_134),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_169),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_134),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_171),
.A2(n_177),
.B1(n_41),
.B2(n_90),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_179),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_123),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_145),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_119),
.Y(n_175)
);

AND3x1_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_8),
.C(n_12),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_113),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_149),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_178),
.A2(n_41),
.B1(n_2),
.B2(n_3),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_105),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_182),
.Y(n_202)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_146),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_176),
.A2(n_150),
.B1(n_144),
.B2(n_156),
.Y(n_183)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_159),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_188),
.C(n_167),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_144),
.B1(n_157),
.B2(n_105),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_177),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_192),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_42),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_193),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_172),
.B(n_8),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_166),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_168),
.B(n_165),
.Y(n_196)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_200),
.B(n_201),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_209),
.C(n_185),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_178),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_206),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_170),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_208),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_164),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_168),
.C(n_162),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_213),
.Y(n_226)
);

OAI321xp33_ASAP7_75t_L g211 ( 
.A1(n_198),
.A2(n_194),
.A3(n_175),
.B1(n_193),
.B2(n_168),
.C(n_170),
.Y(n_211)
);

AOI21x1_ASAP7_75t_SL g223 ( 
.A1(n_211),
.A2(n_197),
.B(n_199),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_182),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_202),
.C(n_205),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_215),
.A2(n_220),
.B(n_11),
.Y(n_229)
);

AOI31xp33_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_180),
.A3(n_170),
.B(n_162),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_218),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_1),
.C(n_2),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_203),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_229),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_214),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_224),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_216),
.B(n_8),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_13),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_228),
.Y(n_231)
);

AOI322xp5_ASAP7_75t_L g234 ( 
.A1(n_227),
.A2(n_210),
.A3(n_220),
.B1(n_215),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_13),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_234),
.A2(n_221),
.B1(n_10),
.B2(n_11),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_226),
.B(n_10),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_235),
.A2(n_236),
.B(n_231),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_2),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_237),
.Y(n_241)
);

AOI21x1_ASAP7_75t_SL g243 ( 
.A1(n_238),
.A2(n_239),
.B(n_240),
.Y(n_243)
);

NOR3xp33_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_3),
.C(n_4),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_4),
.B(n_5),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_240),
.A2(n_230),
.B(n_236),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_5),
.C(n_6),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_245),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_241),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_246),
.A2(n_243),
.B(n_5),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g248 ( 
.A(n_247),
.Y(n_248)
);


endmodule