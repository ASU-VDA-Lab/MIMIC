module real_aes_16977_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_1034;
wire n_549;
wire n_1328;
wire n_571;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1893;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_1883;
wire n_608;
wire n_760;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1346;
wire n_1383;
wire n_552;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1284;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_877;
wire n_424;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_1499;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1853;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_1856;
wire n_658;
wire n_676;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1908;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1899;
wire n_816;
wire n_1470;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1827;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_1226;
wire n_525;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1343;
wire n_719;
wire n_465;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1889;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1823;
wire n_1547;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1891;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1352;
wire n_1323;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g1860 ( .A(n_0), .Y(n_1860) );
AOI22xp33_ASAP7_75t_SL g1248 ( .A1(n_1), .A2(n_335), .B1(n_871), .B2(n_892), .Y(n_1248) );
INVxp67_ASAP7_75t_SL g1274 ( .A(n_1), .Y(n_1274) );
INVx1_ASAP7_75t_L g1423 ( .A(n_2), .Y(n_1423) );
AO22x1_ASAP7_75t_L g1454 ( .A1(n_2), .A2(n_246), .B1(n_451), .B2(n_1008), .Y(n_1454) );
INVx1_ASAP7_75t_L g391 ( .A(n_3), .Y(n_391) );
AND2x2_ASAP7_75t_L g417 ( .A(n_3), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g425 ( .A(n_3), .B(n_269), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_3), .B(n_401), .Y(n_616) );
INVx1_ASAP7_75t_L g1432 ( .A(n_4), .Y(n_1432) );
AOI22xp33_ASAP7_75t_L g1453 ( .A1(n_4), .A2(n_146), .B1(n_419), .B2(n_1019), .Y(n_1453) );
OAI211xp5_ASAP7_75t_SL g1881 ( .A1(n_5), .A2(n_1500), .B(n_1882), .C(n_1883), .Y(n_1881) );
INVx1_ASAP7_75t_L g1902 ( .A(n_5), .Y(n_1902) );
AOI22xp33_ASAP7_75t_SL g891 ( .A1(n_6), .A2(n_333), .B1(n_540), .B2(n_892), .Y(n_891) );
AOI221xp5_ASAP7_75t_L g913 ( .A1(n_6), .A2(n_278), .B1(n_855), .B2(n_914), .C(n_918), .Y(n_913) );
INVx1_ASAP7_75t_L g1067 ( .A(n_7), .Y(n_1067) );
OAI22xp5_ASAP7_75t_L g1142 ( .A1(n_8), .A2(n_235), .B1(n_509), .B2(n_1143), .Y(n_1142) );
AOI22xp33_ASAP7_75t_SL g1553 ( .A1(n_9), .A2(n_239), .B1(n_559), .B2(n_896), .Y(n_1553) );
INVxp67_ASAP7_75t_SL g1575 ( .A(n_9), .Y(n_1575) );
AOI221xp5_ASAP7_75t_L g843 ( .A1(n_10), .A2(n_324), .B1(n_437), .B2(n_456), .C(n_844), .Y(n_843) );
AOI22xp33_ASAP7_75t_SL g872 ( .A1(n_10), .A2(n_351), .B1(n_550), .B2(n_553), .Y(n_872) );
INVxp67_ASAP7_75t_SL g995 ( .A(n_11), .Y(n_995) );
AND4x1_ASAP7_75t_L g1041 ( .A(n_11), .B(n_997), .C(n_1000), .D(n_1021), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g1326 ( .A1(n_12), .A2(n_353), .B1(n_722), .B2(n_857), .Y(n_1326) );
INVx1_ASAP7_75t_L g1341 ( .A(n_12), .Y(n_1341) );
INVx2_ASAP7_75t_L g491 ( .A(n_13), .Y(n_491) );
OAI22xp5_ASAP7_75t_SL g1820 ( .A1(n_14), .A2(n_304), .B1(n_1304), .B2(n_1821), .Y(n_1820) );
OAI221xp5_ASAP7_75t_L g1831 ( .A1(n_14), .A2(n_304), .B1(n_415), .B2(n_976), .C(n_1832), .Y(n_1831) );
AOI22xp5_ASAP7_75t_L g1622 ( .A1(n_15), .A2(n_17), .B1(n_1593), .B2(n_1601), .Y(n_1622) );
INVx1_ASAP7_75t_L g1115 ( .A(n_16), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_18), .A2(n_323), .B1(n_722), .B2(n_723), .Y(n_727) );
INVx1_ASAP7_75t_L g755 ( .A(n_18), .Y(n_755) );
INVx1_ASAP7_75t_L g1530 ( .A(n_19), .Y(n_1530) );
INVx1_ASAP7_75t_L g1864 ( .A(n_20), .Y(n_1864) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_21), .A2(n_285), .B1(n_445), .B2(n_848), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_21), .A2(n_279), .B1(n_871), .B2(n_877), .Y(n_876) );
OAI22xp33_ASAP7_75t_L g1254 ( .A1(n_22), .A2(n_277), .B1(n_772), .B2(n_959), .Y(n_1254) );
INVx1_ASAP7_75t_L g1267 ( .A(n_22), .Y(n_1267) );
INVx1_ASAP7_75t_L g1113 ( .A(n_23), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1129 ( .A1(n_23), .A2(n_79), .B1(n_440), .B2(n_1130), .Y(n_1129) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_24), .A2(n_178), .B1(n_743), .B2(n_964), .Y(n_999) );
OAI211xp5_ASAP7_75t_L g1001 ( .A1(n_24), .A2(n_798), .B(n_1002), .C(n_1005), .Y(n_1001) );
INVx1_ASAP7_75t_L g732 ( .A(n_25), .Y(n_732) );
INVx1_ASAP7_75t_L g1201 ( .A(n_26), .Y(n_1201) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_27), .A2(n_325), .B1(n_743), .B2(n_964), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_28), .A2(n_104), .B1(n_926), .B2(n_1008), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_28), .A2(n_40), .B1(n_1030), .B2(n_1031), .Y(n_1032) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_29), .Y(n_386) );
AND2x2_ASAP7_75t_L g1594 ( .A(n_29), .B(n_384), .Y(n_1594) );
INVx1_ASAP7_75t_L g1830 ( .A(n_30), .Y(n_1830) );
AOI22xp33_ASAP7_75t_L g1661 ( .A1(n_31), .A2(n_209), .B1(n_1601), .B2(n_1662), .Y(n_1661) );
OAI211xp5_ASAP7_75t_SL g797 ( .A1(n_32), .A2(n_798), .B(n_799), .C(n_804), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_32), .A2(n_292), .B1(n_498), .B2(n_509), .Y(n_811) );
OAI22xp5_ASAP7_75t_SL g1504 ( .A1(n_33), .A2(n_310), .B1(n_624), .B2(n_629), .Y(n_1504) );
INVxp67_ASAP7_75t_SL g1534 ( .A(n_33), .Y(n_1534) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_34), .A2(n_237), .B1(n_550), .B2(n_950), .Y(n_954) );
AOI221xp5_ASAP7_75t_L g986 ( .A1(n_34), .A2(n_341), .B1(n_929), .B2(n_987), .C(n_989), .Y(n_986) );
CKINVDCx5p33_ASAP7_75t_R g1538 ( .A(n_35), .Y(n_1538) );
INVx1_ASAP7_75t_L g1151 ( .A(n_36), .Y(n_1151) );
OAI211xp5_ASAP7_75t_L g1159 ( .A1(n_36), .A2(n_716), .B(n_724), .C(n_1160), .Y(n_1159) );
INVxp67_ASAP7_75t_L g883 ( .A(n_37), .Y(n_883) );
CKINVDCx5p33_ASAP7_75t_R g998 ( .A(n_38), .Y(n_998) );
AOI22xp5_ASAP7_75t_L g856 ( .A1(n_39), .A2(n_351), .B1(n_848), .B2(n_857), .Y(n_856) );
AOI22xp5_ASAP7_75t_L g873 ( .A1(n_39), .A2(n_324), .B1(n_550), .B2(n_874), .Y(n_873) );
AOI221xp5_ASAP7_75t_L g1018 ( .A1(n_40), .A2(n_360), .B1(n_719), .B2(n_929), .C(n_1019), .Y(n_1018) );
CKINVDCx5p33_ASAP7_75t_R g612 ( .A(n_41), .Y(n_612) );
AOI21xp33_ASAP7_75t_L g432 ( .A1(n_42), .A2(n_433), .B(n_437), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_42), .A2(n_340), .B1(n_546), .B2(n_550), .Y(n_545) );
INVx1_ASAP7_75t_L g945 ( .A(n_43), .Y(n_945) );
OAI221xp5_ASAP7_75t_L g975 ( .A1(n_43), .A2(n_262), .B1(n_413), .B2(n_976), .C(n_980), .Y(n_975) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_44), .A2(n_129), .B1(n_454), .B2(n_458), .C(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g756 ( .A(n_44), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_45), .B(n_479), .Y(n_785) );
INVx1_ASAP7_75t_L g496 ( .A(n_46), .Y(n_496) );
AOI221xp5_ASAP7_75t_L g1171 ( .A1(n_47), .A2(n_328), .B1(n_437), .B2(n_1019), .C(n_1123), .Y(n_1171) );
INVxp67_ASAP7_75t_SL g1178 ( .A(n_47), .Y(n_1178) );
INVx1_ASAP7_75t_L g1156 ( .A(n_48), .Y(n_1156) );
OAI22xp5_ASAP7_75t_L g1172 ( .A1(n_48), .A2(n_228), .B1(n_798), .B2(n_1173), .Y(n_1172) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_49), .Y(n_592) );
OAI211xp5_ASAP7_75t_SL g646 ( .A1(n_50), .A2(n_639), .B(n_647), .C(n_650), .Y(n_646) );
INVx1_ASAP7_75t_L g696 ( .A(n_50), .Y(n_696) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_51), .Y(n_603) );
INVx1_ASAP7_75t_L g1329 ( .A(n_52), .Y(n_1329) );
AOI22xp33_ASAP7_75t_L g1551 ( .A1(n_53), .A2(n_303), .B1(n_762), .B2(n_899), .Y(n_1551) );
INVx1_ASAP7_75t_L g1568 ( .A(n_53), .Y(n_1568) );
OAI21xp5_ASAP7_75t_L g861 ( .A1(n_54), .A2(n_498), .B(n_862), .Y(n_861) );
NAND5xp2_ASAP7_75t_L g1358 ( .A(n_55), .B(n_1359), .C(n_1378), .D(n_1388), .E(n_1395), .Y(n_1358) );
INVx1_ASAP7_75t_L g1404 ( .A(n_55), .Y(n_1404) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_56), .A2(n_166), .B1(n_743), .B2(n_964), .Y(n_1257) );
OAI211xp5_ASAP7_75t_SL g1259 ( .A1(n_56), .A2(n_798), .B(n_1260), .C(n_1265), .Y(n_1259) );
INVx1_ASAP7_75t_L g1328 ( .A(n_57), .Y(n_1328) );
INVxp67_ASAP7_75t_SL g1170 ( .A(n_58), .Y(n_1170) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_58), .A2(n_158), .B1(n_1189), .B2(n_1190), .Y(n_1188) );
AOI22xp5_ASAP7_75t_L g1675 ( .A1(n_59), .A2(n_229), .B1(n_1593), .B2(n_1598), .Y(n_1675) );
AOI22xp5_ASAP7_75t_L g1608 ( .A1(n_60), .A2(n_356), .B1(n_1601), .B2(n_1609), .Y(n_1608) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_61), .Y(n_398) );
INVx1_ASAP7_75t_L g1003 ( .A(n_62), .Y(n_1003) );
OAI22xp33_ASAP7_75t_L g1024 ( .A1(n_62), .A2(n_114), .B1(n_772), .B2(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g466 ( .A(n_63), .Y(n_466) );
OAI22xp33_ASAP7_75t_L g562 ( .A1(n_63), .A2(n_327), .B1(n_563), .B2(n_569), .Y(n_562) );
XOR2xp5_ASAP7_75t_L g1240 ( .A(n_64), .B(n_1241), .Y(n_1240) );
AOI22xp5_ASAP7_75t_L g1676 ( .A1(n_64), .A2(n_336), .B1(n_1601), .B2(n_1662), .Y(n_1676) );
INVx1_ASAP7_75t_L g1546 ( .A(n_65), .Y(n_1546) );
AOI22xp5_ASAP7_75t_L g1629 ( .A1(n_66), .A2(n_148), .B1(n_1593), .B2(n_1598), .Y(n_1629) );
AOI22xp33_ASAP7_75t_SL g1249 ( .A1(n_67), .A2(n_308), .B1(n_899), .B2(n_1250), .Y(n_1249) );
AOI221xp5_ASAP7_75t_L g1277 ( .A1(n_67), .A2(n_272), .B1(n_731), .B2(n_1278), .C(n_1279), .Y(n_1277) );
INVx1_ASAP7_75t_L g1829 ( .A(n_68), .Y(n_1829) );
INVx1_ASAP7_75t_L g655 ( .A(n_69), .Y(n_655) );
OAI211xp5_ASAP7_75t_L g683 ( .A1(n_69), .A2(n_684), .B(n_686), .C(n_688), .Y(n_683) );
XOR2x2_ASAP7_75t_L g573 ( .A(n_70), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g740 ( .A(n_71), .Y(n_740) );
OAI332xp33_ASAP7_75t_SL g745 ( .A1(n_71), .A2(n_555), .A3(n_746), .B1(n_752), .B2(n_753), .B3(n_759), .C1(n_765), .C2(n_772), .Y(n_745) );
AOI221xp5_ASAP7_75t_L g800 ( .A1(n_72), .A2(n_130), .B1(n_457), .B2(n_801), .C(n_802), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_72), .A2(n_266), .B1(n_561), .B2(n_818), .Y(n_820) );
AOI221xp5_ASAP7_75t_L g1364 ( .A1(n_73), .A2(n_183), .B1(n_419), .B2(n_437), .C(n_1019), .Y(n_1364) );
AOI22xp33_ASAP7_75t_L g1382 ( .A1(n_73), .A2(n_253), .B1(n_550), .B2(n_1383), .Y(n_1382) );
INVx1_ASAP7_75t_L g1216 ( .A(n_74), .Y(n_1216) );
AOI22xp33_ASAP7_75t_L g1365 ( .A1(n_75), .A2(n_253), .B1(n_857), .B2(n_1008), .Y(n_1365) );
AOI22xp33_ASAP7_75t_L g1381 ( .A1(n_75), .A2(n_183), .B1(n_550), .B2(n_762), .Y(n_1381) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_76), .A2(n_175), .B1(n_888), .B2(n_899), .Y(n_898) );
AOI21xp33_ASAP7_75t_L g927 ( .A1(n_76), .A2(n_928), .B(n_929), .Y(n_927) );
AOI221xp5_ASAP7_75t_L g1006 ( .A1(n_77), .A2(n_359), .B1(n_458), .B2(n_928), .C(n_987), .Y(n_1006) );
AOI22xp33_ASAP7_75t_SL g1033 ( .A1(n_77), .A2(n_316), .B1(n_1034), .B2(n_1036), .Y(n_1033) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_78), .A2(n_832), .B1(n_833), .B2(n_879), .Y(n_831) );
INVxp67_ASAP7_75t_SL g879 ( .A(n_78), .Y(n_879) );
INVx1_ASAP7_75t_L g1101 ( .A(n_79), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_80), .A2(n_271), .B1(n_722), .B2(n_723), .Y(n_721) );
INVx1_ASAP7_75t_L g763 ( .A(n_80), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_81), .A2(n_110), .B1(n_440), .B2(n_445), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_81), .A2(n_251), .B1(n_559), .B2(n_561), .Y(n_558) );
AOI22xp33_ASAP7_75t_SL g1205 ( .A1(n_82), .A2(n_307), .B1(n_561), .B2(n_871), .Y(n_1205) );
AOI22xp33_ASAP7_75t_L g1229 ( .A1(n_82), .A2(n_322), .B1(n_848), .B2(n_1227), .Y(n_1229) );
AOI22xp33_ASAP7_75t_SL g1548 ( .A1(n_83), .A2(n_190), .B1(n_540), .B2(n_1346), .Y(n_1548) );
INVxp67_ASAP7_75t_SL g1574 ( .A(n_83), .Y(n_1574) );
INVx1_ASAP7_75t_L g734 ( .A(n_84), .Y(n_734) );
INVx1_ASAP7_75t_L g840 ( .A(n_85), .Y(n_840) );
CKINVDCx5p33_ASAP7_75t_R g902 ( .A(n_86), .Y(n_902) );
OAI21xp5_ASAP7_75t_SL g934 ( .A1(n_87), .A2(n_743), .B(n_935), .Y(n_934) );
CKINVDCx5p33_ASAP7_75t_R g1370 ( .A(n_88), .Y(n_1370) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_89), .A2(n_249), .B1(n_559), .B2(n_948), .Y(n_1060) );
AOI22xp33_ASAP7_75t_SL g1086 ( .A1(n_89), .A2(n_309), .B1(n_722), .B2(n_926), .Y(n_1086) );
AOI22xp33_ASAP7_75t_SL g955 ( .A1(n_90), .A2(n_368), .B1(n_871), .B2(n_956), .Y(n_955) );
AOI221xp5_ASAP7_75t_L g970 ( .A1(n_90), .A2(n_163), .B1(n_855), .B2(n_922), .C(n_971), .Y(n_970) );
CKINVDCx5p33_ASAP7_75t_R g600 ( .A(n_91), .Y(n_600) );
AOI22xp33_ASAP7_75t_SL g895 ( .A1(n_92), .A2(n_278), .B1(n_542), .B2(n_896), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_92), .A2(n_333), .B1(n_925), .B2(n_926), .Y(n_924) );
INVx1_ASAP7_75t_L g842 ( .A(n_93), .Y(n_842) );
OR2x2_ASAP7_75t_L g1154 ( .A(n_94), .B(n_479), .Y(n_1154) );
OAI221xp5_ASAP7_75t_L g1165 ( .A1(n_95), .A2(n_226), .B1(n_976), .B2(n_1166), .C(n_1167), .Y(n_1165) );
OAI322xp33_ASAP7_75t_L g1176 ( .A1(n_95), .A2(n_959), .A3(n_1117), .B1(n_1177), .B2(n_1180), .C1(n_1181), .C2(n_1185), .Y(n_1176) );
AOI22xp33_ASAP7_75t_SL g1059 ( .A1(n_96), .A2(n_242), .B1(n_1056), .B2(n_1058), .Y(n_1059) );
INVx1_ASAP7_75t_L g1081 ( .A(n_96), .Y(n_1081) );
OAI21xp5_ASAP7_75t_L g1237 ( .A1(n_97), .A2(n_743), .B(n_1238), .Y(n_1237) );
AOI22xp33_ASAP7_75t_SL g1507 ( .A1(n_98), .A2(n_176), .B1(n_451), .B2(n_1508), .Y(n_1507) );
INVxp67_ASAP7_75t_SL g1526 ( .A(n_98), .Y(n_1526) );
INVx1_ASAP7_75t_L g1805 ( .A(n_99), .Y(n_1805) );
AOI22xp33_ASAP7_75t_SL g1813 ( .A1(n_100), .A2(n_305), .B1(n_1296), .B2(n_1528), .Y(n_1813) );
AOI221xp5_ASAP7_75t_L g1825 ( .A1(n_100), .A2(n_109), .B1(n_433), .B2(n_855), .C(n_971), .Y(n_1825) );
INVx1_ASAP7_75t_L g1853 ( .A(n_101), .Y(n_1853) );
INVx1_ASAP7_75t_L g1885 ( .A(n_102), .Y(n_1885) );
INVx1_ASAP7_75t_L g1578 ( .A(n_103), .Y(n_1578) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_104), .A2(n_360), .B1(n_1030), .B2(n_1031), .Y(n_1029) );
AOI22xp5_ASAP7_75t_L g1616 ( .A1(n_105), .A2(n_365), .B1(n_1593), .B2(n_1598), .Y(n_1616) );
AOI22xp33_ASAP7_75t_L g1302 ( .A1(n_106), .A2(n_293), .B1(n_871), .B2(n_1296), .Y(n_1302) );
AOI221xp5_ASAP7_75t_L g1308 ( .A1(n_106), .A2(n_288), .B1(n_456), .B2(n_457), .C(n_802), .Y(n_1308) );
INVx1_ASAP7_75t_L g1807 ( .A(n_107), .Y(n_1807) );
INVx1_ASAP7_75t_L g1294 ( .A(n_108), .Y(n_1294) );
AOI22xp33_ASAP7_75t_L g1309 ( .A1(n_108), .A2(n_314), .B1(n_445), .B2(n_925), .Y(n_1309) );
AOI22xp33_ASAP7_75t_L g1819 ( .A1(n_109), .A2(n_205), .B1(n_1189), .B2(n_1346), .Y(n_1819) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_110), .A2(n_276), .B1(n_540), .B2(n_543), .Y(n_539) );
INVx1_ASAP7_75t_L g1112 ( .A(n_111), .Y(n_1112) );
AOI221xp5_ASAP7_75t_L g1122 ( .A1(n_111), .A2(n_243), .B1(n_914), .B2(n_929), .C(n_1123), .Y(n_1122) );
CKINVDCx5p33_ASAP7_75t_R g911 ( .A(n_112), .Y(n_911) );
XNOR2xp5_ASAP7_75t_L g1320 ( .A(n_113), .B(n_1321), .Y(n_1320) );
AOI22xp5_ASAP7_75t_SL g1617 ( .A1(n_113), .A2(n_240), .B1(n_1601), .B2(n_1609), .Y(n_1617) );
INVx1_ASAP7_75t_L g1004 ( .A(n_114), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1206 ( .A1(n_115), .A2(n_338), .B1(n_1207), .B2(n_1208), .Y(n_1206) );
AOI221xp5_ASAP7_75t_L g1230 ( .A1(n_115), .A2(n_362), .B1(n_795), .B2(n_1231), .C(n_1234), .Y(n_1230) );
OAI211xp5_ASAP7_75t_L g1368 ( .A1(n_116), .A2(n_620), .B(n_1082), .C(n_1369), .Y(n_1368) );
INVx1_ASAP7_75t_L g1400 ( .A(n_116), .Y(n_1400) );
INVx1_ASAP7_75t_L g1168 ( .A(n_117), .Y(n_1168) );
CKINVDCx5p33_ASAP7_75t_R g906 ( .A(n_118), .Y(n_906) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_118), .A2(n_139), .B1(n_931), .B2(n_932), .Y(n_930) );
XOR2xp5_ASAP7_75t_L g1800 ( .A(n_119), .B(n_1801), .Y(n_1800) );
AOI22xp33_ASAP7_75t_L g1513 ( .A1(n_120), .A2(n_250), .B1(n_451), .B2(n_463), .Y(n_1513) );
AOI22xp33_ASAP7_75t_L g1523 ( .A1(n_120), .A2(n_273), .B1(n_542), .B2(n_948), .Y(n_1523) );
INVx1_ASAP7_75t_L g791 ( .A(n_121), .Y(n_791) );
AOI21xp33_ASAP7_75t_L g1333 ( .A1(n_122), .A2(n_456), .B(n_795), .Y(n_1333) );
INVx1_ASAP7_75t_L g1340 ( .A(n_122), .Y(n_1340) );
AOI22xp33_ASAP7_75t_L g1213 ( .A1(n_123), .A2(n_322), .B1(n_871), .B2(n_948), .Y(n_1213) );
AOI221xp5_ASAP7_75t_L g1224 ( .A1(n_123), .A2(n_307), .B1(n_802), .B2(n_971), .C(n_1225), .Y(n_1224) );
INVx1_ASAP7_75t_L g1285 ( .A(n_124), .Y(n_1285) );
INVx1_ASAP7_75t_L g1496 ( .A(n_125), .Y(n_1496) );
OAI221xp5_ASAP7_75t_L g1009 ( .A1(n_126), .A2(n_290), .B1(n_413), .B2(n_1010), .C(n_1012), .Y(n_1009) );
INVx1_ASAP7_75t_L g1040 ( .A(n_126), .Y(n_1040) );
INVx1_ASAP7_75t_L g384 ( .A(n_127), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g1325 ( .A1(n_128), .A2(n_270), .B1(n_729), .B2(n_802), .C(n_852), .Y(n_1325) );
AOI22xp33_ASAP7_75t_L g1342 ( .A1(n_128), .A2(n_192), .B1(n_543), .B2(n_871), .Y(n_1342) );
INVx1_ASAP7_75t_L g771 ( .A(n_129), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_130), .A2(n_282), .B1(n_543), .B2(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g805 ( .A(n_131), .Y(n_805) );
OAI22xp33_ASAP7_75t_L g823 ( .A1(n_131), .A2(n_199), .B1(n_569), .B2(n_772), .Y(n_823) );
AOI22xp33_ASAP7_75t_SL g1253 ( .A1(n_132), .A2(n_306), .B1(n_561), .B2(n_871), .Y(n_1253) );
INVxp67_ASAP7_75t_SL g1276 ( .A(n_132), .Y(n_1276) );
AOI22xp33_ASAP7_75t_L g1549 ( .A1(n_133), .A2(n_200), .B1(n_762), .B2(n_1550), .Y(n_1549) );
INVx1_ASAP7_75t_L g1572 ( .A(n_133), .Y(n_1572) );
OAI22xp33_ASAP7_75t_L g1098 ( .A1(n_134), .A2(n_319), .B1(n_772), .B2(n_1025), .Y(n_1098) );
INVx1_ASAP7_75t_L g1133 ( .A(n_134), .Y(n_1133) );
AOI22xp5_ASAP7_75t_L g1613 ( .A1(n_135), .A2(n_345), .B1(n_1598), .B2(n_1609), .Y(n_1613) );
OAI222xp33_ASAP7_75t_L g1440 ( .A1(n_136), .A2(n_355), .B1(n_1441), .B2(n_1443), .C1(n_1445), .C2(n_1447), .Y(n_1440) );
INVx1_ASAP7_75t_L g1458 ( .A(n_136), .Y(n_1458) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_137), .Y(n_589) );
INVx1_ASAP7_75t_L g1869 ( .A(n_138), .Y(n_1869) );
CKINVDCx5p33_ASAP7_75t_R g904 ( .A(n_139), .Y(n_904) );
INVx1_ASAP7_75t_L g426 ( .A(n_140), .Y(n_426) );
INVx1_ASAP7_75t_L g1865 ( .A(n_141), .Y(n_1865) );
INVx1_ASAP7_75t_L g1867 ( .A(n_142), .Y(n_1867) );
OAI211xp5_ASAP7_75t_L g448 ( .A1(n_143), .A2(n_449), .B(n_452), .C(n_465), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_143), .A2(n_286), .B1(n_498), .B2(n_509), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g1889 ( .A1(n_144), .A2(n_154), .B1(n_661), .B2(n_665), .Y(n_1889) );
OAI22xp33_ASAP7_75t_L g1903 ( .A1(n_144), .A2(n_154), .B1(n_1904), .B2(n_1905), .Y(n_1903) );
OAI211xp5_ASAP7_75t_L g1498 ( .A1(n_145), .A2(n_1499), .B(n_1500), .C(n_1501), .Y(n_1498) );
INVxp33_ASAP7_75t_SL g1517 ( .A(n_145), .Y(n_1517) );
INVx1_ASAP7_75t_L g1428 ( .A(n_146), .Y(n_1428) );
CKINVDCx5p33_ASAP7_75t_R g1299 ( .A(n_147), .Y(n_1299) );
INVx1_ASAP7_75t_L g1103 ( .A(n_149), .Y(n_1103) );
AOI221xp5_ASAP7_75t_L g1126 ( .A1(n_149), .A2(n_301), .B1(n_1123), .B2(n_1127), .C(n_1128), .Y(n_1126) );
INVx1_ASAP7_75t_L g1888 ( .A(n_150), .Y(n_1888) );
OAI211xp5_ASAP7_75t_L g1896 ( .A1(n_150), .A2(n_1897), .B(n_1899), .C(n_1900), .Y(n_1896) );
INVx1_ASAP7_75t_L g850 ( .A(n_151), .Y(n_850) );
INVx1_ASAP7_75t_L g1856 ( .A(n_152), .Y(n_1856) );
INVx1_ASAP7_75t_L g1290 ( .A(n_153), .Y(n_1290) );
AOI21xp33_ASAP7_75t_L g1316 ( .A1(n_153), .A2(n_456), .B(n_929), .Y(n_1316) );
INVxp67_ASAP7_75t_SL g428 ( .A(n_155), .Y(n_428) );
AOI22xp33_ASAP7_75t_SL g552 ( .A1(n_155), .A2(n_298), .B1(n_550), .B2(n_553), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g1286 ( .A1(n_156), .A2(n_182), .B1(n_498), .B2(n_964), .Y(n_1286) );
OAI211xp5_ASAP7_75t_L g1306 ( .A1(n_156), .A2(n_449), .B(n_1307), .C(n_1310), .Y(n_1306) );
INVx1_ASAP7_75t_L g1542 ( .A(n_157), .Y(n_1542) );
OAI222xp33_ASAP7_75t_L g1565 ( .A1(n_157), .A2(n_224), .B1(n_716), .B2(n_1010), .C1(n_1566), .C2(n_1573), .Y(n_1565) );
AOI221xp5_ASAP7_75t_L g1164 ( .A1(n_158), .A2(n_238), .B1(n_802), .B2(n_971), .C(n_1019), .Y(n_1164) );
AOI221xp5_ASAP7_75t_L g851 ( .A1(n_159), .A2(n_279), .B1(n_852), .B2(n_853), .C(n_855), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_159), .A2(n_285), .B1(n_543), .B2(n_871), .Y(n_870) );
OAI22xp33_ASAP7_75t_L g1890 ( .A1(n_160), .A2(n_261), .B1(n_1891), .B2(n_1892), .Y(n_1890) );
OAI22xp33_ASAP7_75t_L g1894 ( .A1(n_160), .A2(n_261), .B1(n_679), .B2(n_1895), .Y(n_1894) );
INVx1_ASAP7_75t_L g1049 ( .A(n_161), .Y(n_1049) );
OAI221xp5_ASAP7_75t_L g1078 ( .A1(n_161), .A2(n_162), .B1(n_1011), .B2(n_1079), .C(n_1080), .Y(n_1078) );
INVx1_ASAP7_75t_L g1050 ( .A(n_162), .Y(n_1050) );
AOI22xp33_ASAP7_75t_SL g947 ( .A1(n_163), .A2(n_206), .B1(n_871), .B2(n_948), .Y(n_947) );
OA21x2_ASAP7_75t_L g1803 ( .A1(n_164), .A2(n_479), .B(n_1804), .Y(n_1803) );
CKINVDCx5p33_ASAP7_75t_R g654 ( .A(n_165), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_167), .A2(n_341), .B1(n_950), .B2(n_952), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_167), .A2(n_237), .B1(n_723), .B2(n_969), .Y(n_968) );
OAI22xp33_ASAP7_75t_L g668 ( .A1(n_168), .A2(n_320), .B1(n_669), .B2(n_670), .Y(n_668) );
OAI22xp33_ASAP7_75t_L g676 ( .A1(n_168), .A2(n_320), .B1(n_677), .B2(n_680), .Y(n_676) );
INVx1_ASAP7_75t_L g835 ( .A(n_169), .Y(n_835) );
INVx1_ASAP7_75t_L g1557 ( .A(n_170), .Y(n_1557) );
CKINVDCx5p33_ASAP7_75t_R g962 ( .A(n_171), .Y(n_962) );
OAI221xp5_ASAP7_75t_L g1330 ( .A1(n_172), .A2(n_363), .B1(n_1011), .B2(n_1079), .C(n_1331), .Y(n_1330) );
OAI22xp33_ASAP7_75t_L g1347 ( .A1(n_172), .A2(n_363), .B1(n_776), .B2(n_1304), .Y(n_1347) );
AO22x1_ASAP7_75t_L g887 ( .A1(n_173), .A2(n_214), .B1(n_822), .B2(n_888), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_173), .B(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g1394 ( .A(n_174), .Y(n_1394) );
AOI22xp33_ASAP7_75t_SL g919 ( .A1(n_175), .A2(n_214), .B1(n_723), .B2(n_848), .Y(n_919) );
INVx1_ASAP7_75t_L g1522 ( .A(n_176), .Y(n_1522) );
CKINVDCx5p33_ASAP7_75t_R g1256 ( .A(n_177), .Y(n_1256) );
OA22x2_ASAP7_75t_L g786 ( .A1(n_179), .A2(n_787), .B1(n_824), .B2(n_825), .Y(n_786) );
CKINVDCx16_ASAP7_75t_R g824 ( .A(n_179), .Y(n_824) );
OAI211xp5_ASAP7_75t_L g412 ( .A1(n_180), .A2(n_413), .B(n_421), .C(n_427), .Y(n_412) );
INVx1_ASAP7_75t_L g528 ( .A(n_180), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g1503 ( .A(n_181), .Y(n_1503) );
INVx1_ASAP7_75t_L g1424 ( .A(n_184), .Y(n_1424) );
AOI22xp33_ASAP7_75t_L g1474 ( .A1(n_184), .A2(n_281), .B1(n_857), .B2(n_1008), .Y(n_1474) );
INVx1_ASAP7_75t_L g810 ( .A(n_185), .Y(n_810) );
INVx1_ASAP7_75t_L g1239 ( .A(n_186), .Y(n_1239) );
INVx1_ASAP7_75t_L g1658 ( .A(n_187), .Y(n_1658) );
AOI22xp5_ASAP7_75t_SL g1628 ( .A1(n_188), .A2(n_198), .B1(n_1601), .B2(n_1609), .Y(n_1628) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_189), .A2(n_295), .B1(n_659), .B2(n_663), .Y(n_658) );
OAI22xp33_ASAP7_75t_L g697 ( .A1(n_189), .A2(n_295), .B1(n_698), .B2(n_701), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g1562 ( .A1(n_190), .A2(n_239), .B1(n_458), .B2(n_1278), .C(n_1279), .Y(n_1562) );
CKINVDCx5p33_ASAP7_75t_R g1502 ( .A(n_191), .Y(n_1502) );
AOI22xp33_ASAP7_75t_SL g1334 ( .A1(n_192), .A2(n_334), .B1(n_451), .B2(n_848), .Y(n_1334) );
OAI211xp5_ASAP7_75t_L g1323 ( .A1(n_193), .A2(n_449), .B(n_1324), .C(n_1327), .Y(n_1323) );
OAI22xp5_ASAP7_75t_L g1350 ( .A1(n_193), .A2(n_358), .B1(n_498), .B2(n_964), .Y(n_1350) );
INVx1_ASAP7_75t_L g1511 ( .A(n_194), .Y(n_1511) );
AOI22xp33_ASAP7_75t_SL g1055 ( .A1(n_195), .A2(n_311), .B1(n_1056), .B2(n_1058), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_195), .A2(n_242), .B1(n_445), .B2(n_1074), .Y(n_1073) );
INVx1_ASAP7_75t_L g1812 ( .A(n_196), .Y(n_1812) );
AOI221xp5_ASAP7_75t_L g1838 ( .A1(n_196), .A2(n_241), .B1(n_731), .B2(n_853), .C(n_1231), .Y(n_1838) );
OAI211xp5_ASAP7_75t_L g1360 ( .A1(n_197), .A2(n_1361), .B(n_1362), .C(n_1367), .Y(n_1360) );
NOR2xp33_ASAP7_75t_L g1377 ( .A(n_197), .B(n_509), .Y(n_1377) );
XNOR2x2_ASAP7_75t_L g939 ( .A(n_198), .B(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g808 ( .A(n_199), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g1563 ( .A1(n_200), .A2(n_303), .B1(n_969), .B2(n_1130), .Y(n_1563) );
INVx2_ASAP7_75t_L g1596 ( .A(n_201), .Y(n_1596) );
AND2x2_ASAP7_75t_L g1599 ( .A(n_201), .B(n_1597), .Y(n_1599) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_201), .B(n_315), .Y(n_1604) );
CKINVDCx5p33_ASAP7_75t_R g1175 ( .A(n_202), .Y(n_1175) );
INVx1_ASAP7_75t_L g1312 ( .A(n_203), .Y(n_1312) );
AOI22xp5_ASAP7_75t_SL g1621 ( .A1(n_204), .A2(n_274), .B1(n_1598), .B2(n_1603), .Y(n_1621) );
INVx1_ASAP7_75t_L g1837 ( .A(n_205), .Y(n_1837) );
INVxp67_ASAP7_75t_SL g982 ( .A(n_206), .Y(n_982) );
XNOR2xp5_ASAP7_75t_L g409 ( .A(n_207), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g1222 ( .A(n_208), .Y(n_1222) );
XOR2x2_ASAP7_75t_L g711 ( .A(n_209), .B(n_712), .Y(n_711) );
CKINVDCx5p33_ASAP7_75t_R g910 ( .A(n_210), .Y(n_910) );
AOI22xp5_ASAP7_75t_L g1600 ( .A1(n_211), .A2(n_343), .B1(n_1601), .B2(n_1603), .Y(n_1600) );
OAI22xp33_ASAP7_75t_L g958 ( .A1(n_212), .A2(n_284), .B1(n_563), .B2(n_959), .Y(n_958) );
INVx1_ASAP7_75t_L g973 ( .A(n_212), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_213), .A2(n_362), .B1(n_1031), .B2(n_1207), .Y(n_1209) );
AOI22xp33_ASAP7_75t_L g1226 ( .A1(n_213), .A2(n_338), .B1(n_722), .B2(n_1227), .Y(n_1226) );
AOI22xp5_ASAP7_75t_L g1607 ( .A1(n_215), .A2(n_280), .B1(n_1593), .B2(n_1598), .Y(n_1607) );
INVx1_ASAP7_75t_L g1485 ( .A(n_216), .Y(n_1485) );
INVx1_ASAP7_75t_L g1556 ( .A(n_217), .Y(n_1556) );
AOI22xp33_ASAP7_75t_L g1363 ( .A1(n_218), .A2(n_300), .B1(n_463), .B2(n_857), .Y(n_1363) );
AOI22xp33_ASAP7_75t_SL g1384 ( .A1(n_218), .A2(n_313), .B1(n_871), .B2(n_877), .Y(n_1384) );
AOI22xp33_ASAP7_75t_SL g1295 ( .A1(n_219), .A2(n_288), .B1(n_871), .B2(n_1296), .Y(n_1295) );
AOI22xp33_ASAP7_75t_SL g1317 ( .A1(n_219), .A2(n_293), .B1(n_848), .B2(n_926), .Y(n_1317) );
AOI21xp33_ASAP7_75t_L g794 ( .A1(n_220), .A2(n_729), .B(n_795), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_220), .A2(n_342), .B1(n_546), .B2(n_550), .Y(n_819) );
INVx1_ASAP7_75t_L g1107 ( .A(n_221), .Y(n_1107) );
OAI211xp5_ASAP7_75t_L g789 ( .A1(n_222), .A2(n_413), .B(n_790), .C(n_792), .Y(n_789) );
INVx1_ASAP7_75t_L g815 ( .A(n_222), .Y(n_815) );
INVx1_ASAP7_75t_L g1818 ( .A(n_223), .Y(n_1818) );
AOI22xp33_ASAP7_75t_L g1826 ( .A1(n_223), .A2(n_294), .B1(n_857), .B2(n_1827), .Y(n_1826) );
INVx1_ASAP7_75t_L g1543 ( .A(n_224), .Y(n_1543) );
AOI22xp5_ASAP7_75t_L g1614 ( .A1(n_225), .A2(n_299), .B1(n_1593), .B2(n_1601), .Y(n_1614) );
INVx1_ASAP7_75t_L g1150 ( .A(n_226), .Y(n_1150) );
CKINVDCx5p33_ASAP7_75t_R g1426 ( .A(n_227), .Y(n_1426) );
INVx1_ASAP7_75t_L g1153 ( .A(n_228), .Y(n_1153) );
CKINVDCx5p33_ASAP7_75t_R g1332 ( .A(n_230), .Y(n_1332) );
OAI22xp5_ASAP7_75t_L g1068 ( .A1(n_231), .A2(n_370), .B1(n_563), .B2(n_959), .Y(n_1068) );
INVx1_ASAP7_75t_L g1076 ( .A(n_231), .Y(n_1076) );
INVx1_ASAP7_75t_L g1191 ( .A(n_232), .Y(n_1191) );
CKINVDCx5p33_ASAP7_75t_R g1373 ( .A(n_233), .Y(n_1373) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_234), .B(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g519 ( .A(n_234), .Y(n_519) );
INVx1_ASAP7_75t_L g557 ( .A(n_234), .Y(n_557) );
OAI211xp5_ASAP7_75t_L g1124 ( .A1(n_235), .A2(n_449), .B(n_1125), .C(n_1132), .Y(n_1124) );
INVx1_ASAP7_75t_L g1436 ( .A(n_236), .Y(n_1436) );
NAND2xp33_ASAP7_75t_SL g1475 ( .A(n_236), .B(n_419), .Y(n_1475) );
INVx1_ASAP7_75t_L g1184 ( .A(n_238), .Y(n_1184) );
INVx1_ASAP7_75t_L g1817 ( .A(n_241), .Y(n_1817) );
INVx1_ASAP7_75t_L g1109 ( .A(n_243), .Y(n_1109) );
INVx1_ASAP7_75t_L g1163 ( .A(n_244), .Y(n_1163) );
OAI22xp5_ASAP7_75t_L g1376 ( .A1(n_245), .A2(n_321), .B1(n_429), .B2(n_620), .Y(n_1376) );
INVx1_ASAP7_75t_L g1398 ( .A(n_245), .Y(n_1398) );
AOI21xp5_ASAP7_75t_L g1437 ( .A1(n_246), .A2(n_556), .B(n_1035), .Y(n_1437) );
INVx1_ASAP7_75t_L g1479 ( .A(n_247), .Y(n_1479) );
BUFx3_ASAP7_75t_L g484 ( .A(n_248), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g1072 ( .A1(n_249), .A2(n_258), .B1(n_456), .B2(n_457), .C(n_802), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g1527 ( .A1(n_250), .A2(n_296), .B1(n_948), .B2(n_1528), .Y(n_1527) );
AOI221xp5_ASAP7_75t_L g453 ( .A1(n_251), .A2(n_276), .B1(n_454), .B2(n_457), .C(n_458), .Y(n_453) );
INVx1_ASAP7_75t_L g744 ( .A(n_252), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g1215 ( .A(n_254), .Y(n_1215) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_255), .A2(n_259), .B1(n_776), .B2(n_1096), .Y(n_1095) );
OAI221xp5_ASAP7_75t_L g1120 ( .A1(n_255), .A2(n_259), .B1(n_413), .B2(n_1010), .C(n_1121), .Y(n_1120) );
AOI22xp5_ASAP7_75t_L g1592 ( .A1(n_256), .A2(n_297), .B1(n_1593), .B2(n_1598), .Y(n_1592) );
INVx1_ASAP7_75t_L g1415 ( .A(n_257), .Y(n_1415) );
NOR2xp33_ASAP7_75t_L g1417 ( .A(n_257), .B(n_1418), .Y(n_1417) );
AOI22xp33_ASAP7_75t_SL g1054 ( .A1(n_258), .A2(n_309), .B1(n_540), .B2(n_948), .Y(n_1054) );
AOI21xp33_ASAP7_75t_L g1512 ( .A1(n_260), .A2(n_437), .B(n_456), .Y(n_1512) );
INVx1_ASAP7_75t_L g1521 ( .A(n_260), .Y(n_1521) );
INVx1_ASAP7_75t_L g944 ( .A(n_262), .Y(n_944) );
AOI22xp5_ASAP7_75t_L g1091 ( .A1(n_263), .A2(n_1092), .B1(n_1093), .B2(n_1144), .Y(n_1091) );
INVx1_ASAP7_75t_L g1144 ( .A(n_263), .Y(n_1144) );
INVx1_ASAP7_75t_L g1220 ( .A(n_264), .Y(n_1220) );
XOR2x2_ASAP7_75t_L g1491 ( .A(n_265), .B(n_1492), .Y(n_1491) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_266), .A2(n_282), .B1(n_440), .B2(n_445), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_267), .B(n_1045), .Y(n_1044) );
AOI22xp5_ASAP7_75t_L g1063 ( .A1(n_267), .A2(n_1064), .B1(n_1065), .B2(n_1087), .Y(n_1063) );
INVx1_ASAP7_75t_L g1089 ( .A(n_267), .Y(n_1089) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_268), .Y(n_582) );
BUFx3_ASAP7_75t_L g401 ( .A(n_269), .Y(n_401) );
INVx1_ASAP7_75t_L g418 ( .A(n_269), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g1345 ( .A1(n_270), .A2(n_334), .B1(n_871), .B2(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g749 ( .A(n_271), .Y(n_749) );
AOI22xp33_ASAP7_75t_SL g1252 ( .A1(n_272), .A2(n_326), .B1(n_899), .B2(n_1250), .Y(n_1252) );
NAND2xp5_ASAP7_75t_SL g1506 ( .A(n_273), .B(n_456), .Y(n_1506) );
AOI22xp33_ASAP7_75t_L g1844 ( .A1(n_274), .A2(n_1845), .B1(n_1847), .B2(n_1908), .Y(n_1844) );
XNOR2xp5_ASAP7_75t_L g1848 ( .A(n_274), .B(n_1849), .Y(n_1848) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_275), .A2(n_342), .B1(n_445), .B2(n_461), .Y(n_803) );
AOI22xp33_ASAP7_75t_SL g821 ( .A1(n_275), .A2(n_354), .B1(n_553), .B2(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g1266 ( .A(n_277), .Y(n_1266) );
INVx1_ASAP7_75t_L g1433 ( .A(n_281), .Y(n_1433) );
INVx1_ASAP7_75t_L g1862 ( .A(n_283), .Y(n_1862) );
INVx1_ASAP7_75t_L g974 ( .A(n_284), .Y(n_974) );
CKINVDCx5p33_ASAP7_75t_R g1062 ( .A(n_287), .Y(n_1062) );
INVx1_ASAP7_75t_L g1161 ( .A(n_289), .Y(n_1161) );
INVx1_ASAP7_75t_L g1038 ( .A(n_290), .Y(n_1038) );
INVx1_ASAP7_75t_L g1311 ( .A(n_291), .Y(n_1311) );
NAND2xp33_ASAP7_75t_SL g1814 ( .A(n_294), .B(n_1550), .Y(n_1814) );
NAND2xp5_ASAP7_75t_SL g1509 ( .A(n_296), .B(n_971), .Y(n_1509) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_298), .A2(n_340), .B1(n_445), .B2(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_SL g1380 ( .A1(n_300), .A2(n_373), .B1(n_871), .B2(n_1296), .Y(n_1380) );
INVx1_ASAP7_75t_L g1116 ( .A(n_301), .Y(n_1116) );
INVx1_ASAP7_75t_L g485 ( .A(n_302), .Y(n_485) );
INVx1_ASAP7_75t_L g515 ( .A(n_302), .Y(n_515) );
INVx1_ASAP7_75t_L g1834 ( .A(n_305), .Y(n_1834) );
AOI221xp5_ASAP7_75t_L g1261 ( .A1(n_306), .A2(n_335), .B1(n_458), .B2(n_1225), .C(n_1262), .Y(n_1261) );
AOI22xp33_ASAP7_75t_L g1264 ( .A1(n_308), .A2(n_326), .B1(n_722), .B2(n_1227), .Y(n_1264) );
OAI21xp33_ASAP7_75t_L g1515 ( .A1(n_310), .A2(n_569), .B(n_1516), .Y(n_1515) );
AOI21xp33_ASAP7_75t_L g1084 ( .A1(n_311), .A2(n_929), .B(n_1085), .Y(n_1084) );
CKINVDCx5p33_ASAP7_75t_R g1413 ( .A(n_312), .Y(n_1413) );
AOI221xp5_ASAP7_75t_SL g1366 ( .A1(n_313), .A2(n_373), .B1(n_419), .B2(n_855), .C(n_916), .Y(n_1366) );
INVx1_ASAP7_75t_L g1301 ( .A(n_314), .Y(n_1301) );
INVx1_ASAP7_75t_L g1597 ( .A(n_315), .Y(n_1597) );
AND2x2_ASAP7_75t_L g1602 ( .A(n_315), .B(n_1596), .Y(n_1602) );
INVxp67_ASAP7_75t_SL g1017 ( .A(n_316), .Y(n_1017) );
INVx1_ASAP7_75t_L g735 ( .A(n_317), .Y(n_735) );
INVx1_ASAP7_75t_L g860 ( .A(n_318), .Y(n_860) );
INVx1_ASAP7_75t_L g1134 ( .A(n_319), .Y(n_1134) );
INVx1_ASAP7_75t_L g1387 ( .A(n_321), .Y(n_1387) );
INVx1_ASAP7_75t_L g766 ( .A(n_323), .Y(n_766) );
OAI211xp5_ASAP7_75t_L g966 ( .A1(n_325), .A2(n_798), .B(n_967), .C(n_972), .Y(n_966) );
INVx1_ASAP7_75t_L g469 ( .A(n_327), .Y(n_469) );
INVxp67_ASAP7_75t_SL g1186 ( .A(n_328), .Y(n_1186) );
INVx1_ASAP7_75t_L g859 ( .A(n_329), .Y(n_859) );
INVxp67_ASAP7_75t_SL g1052 ( .A(n_330), .Y(n_1052) );
OAI211xp5_ASAP7_75t_L g1070 ( .A1(n_330), .A2(n_449), .B(n_1071), .C(n_1075), .Y(n_1070) );
INVx1_ASAP7_75t_L g1660 ( .A(n_331), .Y(n_1660) );
CKINVDCx16_ASAP7_75t_R g1442 ( .A(n_332), .Y(n_1442) );
CKINVDCx5p33_ASAP7_75t_R g610 ( .A(n_337), .Y(n_610) );
OAI21xp33_ASAP7_75t_L g1554 ( .A1(n_339), .A2(n_743), .B(n_1555), .Y(n_1554) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_344), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g937 ( .A(n_346), .Y(n_937) );
OAI211xp5_ASAP7_75t_L g715 ( .A1(n_347), .A2(n_716), .B(n_717), .C(n_724), .Y(n_715) );
INVx1_ASAP7_75t_L g777 ( .A(n_347), .Y(n_777) );
AOI221xp5_ASAP7_75t_L g728 ( .A1(n_348), .A2(n_367), .B1(n_457), .B2(n_729), .C(n_731), .Y(n_728) );
INVx1_ASAP7_75t_L g747 ( .A(n_348), .Y(n_747) );
CKINVDCx5p33_ASAP7_75t_R g1202 ( .A(n_349), .Y(n_1202) );
INVxp67_ASAP7_75t_SL g1013 ( .A(n_350), .Y(n_1013) );
AOI22xp33_ASAP7_75t_SL g1027 ( .A1(n_350), .A2(n_359), .B1(n_542), .B2(n_1028), .Y(n_1027) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_352), .Y(n_397) );
INVx1_ASAP7_75t_L g1344 ( .A(n_353), .Y(n_1344) );
INVxp67_ASAP7_75t_SL g793 ( .A(n_354), .Y(n_793) );
NOR2xp33_ASAP7_75t_R g1465 ( .A(n_355), .B(n_1466), .Y(n_1465) );
INVx1_ASAP7_75t_L g1409 ( .A(n_356), .Y(n_1409) );
INVx1_ASAP7_75t_L g1245 ( .A(n_357), .Y(n_1245) );
OAI221xp5_ASAP7_75t_SL g1270 ( .A1(n_357), .A2(n_374), .B1(n_413), .B2(n_1010), .C(n_1271), .Y(n_1270) );
INVx1_ASAP7_75t_L g1349 ( .A(n_361), .Y(n_1349) );
INVx2_ASAP7_75t_L g476 ( .A(n_364), .Y(n_476) );
INVx1_ASAP7_75t_L g489 ( .A(n_364), .Y(n_489) );
INVx1_ASAP7_75t_L g494 ( .A(n_364), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g1141 ( .A(n_366), .Y(n_1141) );
INVxp67_ASAP7_75t_SL g760 ( .A(n_367), .Y(n_760) );
INVxp67_ASAP7_75t_SL g985 ( .A(n_368), .Y(n_985) );
OAI22xp33_ASAP7_75t_SL g1303 ( .A1(n_369), .A2(n_372), .B1(n_776), .B2(n_1304), .Y(n_1303) );
OAI221xp5_ASAP7_75t_L g1313 ( .A1(n_369), .A2(n_372), .B1(n_413), .B2(n_1011), .C(n_1314), .Y(n_1313) );
INVx1_ASAP7_75t_L g1077 ( .A(n_370), .Y(n_1077) );
XNOR2xp5_ASAP7_75t_L g1282 ( .A(n_371), .B(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1246 ( .A(n_374), .Y(n_1246) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_402), .B(n_1582), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx4f_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_387), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g1846 ( .A(n_381), .B(n_390), .Y(n_1846) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g1843 ( .A(n_383), .B(n_386), .Y(n_1843) );
INVx1_ASAP7_75t_L g1911 ( .A(n_383), .Y(n_1911) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g1913 ( .A(n_386), .B(n_1911), .Y(n_1913) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_392), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g673 ( .A(n_390), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g438 ( .A(n_391), .B(n_400), .Y(n_438) );
AND2x4_ASAP7_75t_L g459 ( .A(n_391), .B(n_401), .Y(n_459) );
INVx1_ASAP7_75t_L g669 ( .A(n_392), .Y(n_669) );
AND2x4_ASAP7_75t_SL g1845 ( .A(n_392), .B(n_1846), .Y(n_1845) );
INVx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x6_ASAP7_75t_L g393 ( .A(n_394), .B(n_399), .Y(n_393) );
OR2x6_ASAP7_75t_L g661 ( .A(n_394), .B(n_662), .Y(n_661) );
BUFx4f_ASAP7_75t_L g1879 ( .A(n_394), .Y(n_1879) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx4f_ASAP7_75t_L g621 ( .A(n_395), .Y(n_621) );
INVx3_ASAP7_75t_L g638 ( .A(n_395), .Y(n_638) );
INVx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
AND2x2_ASAP7_75t_L g420 ( .A(n_397), .B(n_398), .Y(n_420) );
NAND2x1_ASAP7_75t_L g431 ( .A(n_397), .B(n_398), .Y(n_431) );
AND2x2_ASAP7_75t_L g435 ( .A(n_397), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g443 ( .A(n_397), .Y(n_443) );
INVx2_ASAP7_75t_L g447 ( .A(n_397), .Y(n_447) );
INVx1_ASAP7_75t_L g507 ( .A(n_397), .Y(n_507) );
BUFx2_ASAP7_75t_L g424 ( .A(n_398), .Y(n_424) );
INVx2_ASAP7_75t_L g436 ( .A(n_398), .Y(n_436) );
INVx1_ASAP7_75t_L g444 ( .A(n_398), .Y(n_444) );
AND2x2_ASAP7_75t_L g446 ( .A(n_398), .B(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_398), .B(n_447), .Y(n_627) );
OR2x2_ASAP7_75t_L g630 ( .A(n_398), .B(n_443), .Y(n_630) );
OR2x6_ASAP7_75t_L g1891 ( .A(n_399), .B(n_638), .Y(n_1891) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g649 ( .A(n_400), .Y(n_649) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g653 ( .A(n_401), .Y(n_653) );
AND2x4_ASAP7_75t_L g657 ( .A(n_401), .B(n_506), .Y(n_657) );
OAI22xp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B1(n_1193), .B2(n_1194), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_990), .B1(n_991), .B2(n_1192), .Y(n_404) );
INVx1_ASAP7_75t_L g1192 ( .A(n_405), .Y(n_1192) );
XNOR2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_829), .Y(n_405) );
AO22x2_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_709), .B1(n_827), .B2(n_828), .Y(n_406) );
INVx1_ASAP7_75t_L g827 ( .A(n_407), .Y(n_827) );
XNOR2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_573), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND3xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_477), .C(n_521), .Y(n_410) );
OAI21xp5_ASAP7_75t_SL g411 ( .A1(n_412), .A2(n_448), .B(n_472), .Y(n_411) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g716 ( .A(n_414), .Y(n_716) );
INVx2_ASAP7_75t_L g1079 ( .A(n_414), .Y(n_1079) );
INVx4_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx3_ASAP7_75t_L g841 ( .A(n_416), .Y(n_841) );
AND2x4_ASAP7_75t_SL g416 ( .A(n_417), .B(n_419), .Y(n_416) );
AND2x4_ASAP7_75t_L g450 ( .A(n_417), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g468 ( .A(n_417), .B(n_442), .Y(n_468) );
AND2x4_ASAP7_75t_L g471 ( .A(n_417), .B(n_434), .Y(n_471) );
AND2x2_ASAP7_75t_L g736 ( .A(n_417), .B(n_737), .Y(n_736) );
BUFx2_ASAP7_75t_L g1375 ( .A(n_417), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_417), .B(n_434), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_417), .B(n_494), .Y(n_1467) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_418), .Y(n_662) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_419), .Y(n_457) );
AND2x6_ASAP7_75t_L g464 ( .A(n_419), .B(n_425), .Y(n_464) );
AND2x2_ASAP7_75t_L g648 ( .A(n_419), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g720 ( .A(n_419), .Y(n_720) );
BUFx3_ASAP7_75t_L g852 ( .A(n_419), .Y(n_852) );
BUFx3_ASAP7_75t_L g971 ( .A(n_419), .Y(n_971) );
BUFx3_ASAP7_75t_L g989 ( .A(n_419), .Y(n_989) );
BUFx3_ASAP7_75t_L g1123 ( .A(n_419), .Y(n_1123) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g846 ( .A(n_420), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_426), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_422), .A2(n_727), .B1(n_728), .B2(n_732), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_422), .B(n_791), .Y(n_790) );
AOI222xp33_ASAP7_75t_L g839 ( .A1(n_422), .A2(n_840), .B1(n_841), .B2(n_842), .C1(n_843), .C2(n_847), .Y(n_839) );
INVx1_ASAP7_75t_L g932 ( .A(n_422), .Y(n_932) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_425), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g1369 ( .A1(n_423), .A2(n_1370), .B1(n_1371), .B2(n_1373), .Y(n_1369) );
AOI22xp33_ASAP7_75t_L g1501 ( .A1(n_423), .A2(n_1371), .B1(n_1502), .B2(n_1503), .Y(n_1501) );
BUFx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g652 ( .A(n_424), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g978 ( .A(n_424), .Y(n_978) );
INVx1_ASAP7_75t_L g1464 ( .A(n_424), .Y(n_1464) );
AND2x2_ASAP7_75t_L g1884 ( .A(n_424), .B(n_653), .Y(n_1884) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_425), .B(n_442), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_425), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g979 ( .A(n_425), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g1462 ( .A(n_425), .B(n_476), .Y(n_1462) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_426), .A2(n_524), .B1(n_528), .B2(n_529), .Y(n_523) );
OAI211xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_429), .B(n_432), .C(n_439), .Y(n_427) );
OAI211xp5_ASAP7_75t_L g792 ( .A1(n_429), .A2(n_793), .B(n_794), .C(n_796), .Y(n_792) );
BUFx4f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx4_ASAP7_75t_L g1083 ( .A(n_430), .Y(n_1083) );
OR2x6_ASAP7_75t_L g1476 ( .A(n_430), .B(n_1477), .Y(n_1476) );
BUFx4f_ASAP7_75t_L g1567 ( .A(n_430), .Y(n_1567) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx3_ASAP7_75t_L g633 ( .A(n_431), .Y(n_633) );
BUFx3_ASAP7_75t_L g1279 ( .A(n_433), .Y(n_1279) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g730 ( .A(n_434), .Y(n_730) );
INVx2_ASAP7_75t_L g854 ( .A(n_434), .Y(n_854) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx3_ASAP7_75t_L g456 ( .A(n_435), .Y(n_456) );
AND2x4_ASAP7_75t_L g671 ( .A(n_435), .B(n_662), .Y(n_671) );
INVx2_ASAP7_75t_L g917 ( .A(n_435), .Y(n_917) );
INVx3_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g731 ( .A(n_438), .Y(n_731) );
INVx1_ASAP7_75t_L g795 ( .A(n_438), .Y(n_795) );
INVx2_ASAP7_75t_L g929 ( .A(n_438), .Y(n_929) );
OAI221xp5_ASAP7_75t_L g1566 ( .A1(n_438), .A2(n_1567), .B1(n_1568), .B2(n_1569), .C(n_1572), .Y(n_1566) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g722 ( .A(n_441), .Y(n_722) );
INVx2_ASAP7_75t_SL g848 ( .A(n_441), .Y(n_848) );
INVx2_ASAP7_75t_L g969 ( .A(n_441), .Y(n_969) );
INVx2_ASAP7_75t_L g1008 ( .A(n_441), .Y(n_1008) );
INVx1_ASAP7_75t_L g1508 ( .A(n_441), .Y(n_1508) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_442), .Y(n_463) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
HB1xp67_ASAP7_75t_L g1372 ( .A(n_443), .Y(n_1372) );
INVx1_ASAP7_75t_SL g1131 ( .A(n_445), .Y(n_1131) );
BUFx3_ASAP7_75t_L g1227 ( .A(n_445), .Y(n_1227) );
BUFx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_446), .Y(n_451) );
INVx2_ASAP7_75t_L g738 ( .A(n_446), .Y(n_738) );
BUFx3_ASAP7_75t_L g857 ( .A(n_446), .Y(n_857) );
INVx2_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
INVx3_ASAP7_75t_L g798 ( .A(n_450), .Y(n_798) );
AOI221xp5_ASAP7_75t_SL g912 ( .A1(n_450), .A2(n_464), .B1(n_902), .B2(n_913), .C(n_919), .Y(n_912) );
AOI221xp5_ASAP7_75t_L g1223 ( .A1(n_450), .A2(n_464), .B1(n_1201), .B2(n_1224), .C(n_1226), .Y(n_1223) );
NAND2xp5_ASAP7_75t_R g1564 ( .A(n_450), .B(n_1546), .Y(n_1564) );
BUFx2_ASAP7_75t_L g723 ( .A(n_451), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_460), .B(n_464), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g1085 ( .A(n_455), .Y(n_1085) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_456), .Y(n_801) );
BUFx2_ASAP7_75t_L g1225 ( .A(n_456), .Y(n_1225) );
INVx1_ASAP7_75t_L g1263 ( .A(n_457), .Y(n_1263) );
INVx1_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_459), .B(n_643), .Y(n_642) );
INVx4_ASAP7_75t_L g802 ( .A(n_459), .Y(n_802) );
INVx4_ASAP7_75t_L g855 ( .A(n_459), .Y(n_855) );
AND2x2_ASAP7_75t_SL g1470 ( .A(n_459), .B(n_487), .Y(n_1470) );
NAND4xp25_ASAP7_75t_L g1505 ( .A(n_459), .B(n_1506), .C(n_1507), .D(n_1509), .Y(n_1505) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_SL g925 ( .A(n_462), .Y(n_925) );
INVx1_ASAP7_75t_L g1827 ( .A(n_462), .Y(n_1827) );
INVx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx6f_ASAP7_75t_L g1074 ( .A(n_463), .Y(n_1074) );
INVx1_ASAP7_75t_L g724 ( .A(n_464), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g799 ( .A1(n_464), .A2(n_800), .B(n_803), .Y(n_799) );
AOI221xp5_ASAP7_75t_L g849 ( .A1(n_464), .A2(n_736), .B1(n_850), .B2(n_851), .C(n_856), .Y(n_849) );
AOI21xp5_ASAP7_75t_L g967 ( .A1(n_464), .A2(n_968), .B(n_970), .Y(n_967) );
AOI21xp5_ASAP7_75t_L g1005 ( .A1(n_464), .A2(n_1006), .B(n_1007), .Y(n_1005) );
AOI21xp5_ASAP7_75t_L g1071 ( .A1(n_464), .A2(n_1072), .B(n_1073), .Y(n_1071) );
AOI21xp5_ASAP7_75t_L g1125 ( .A1(n_464), .A2(n_1126), .B(n_1129), .Y(n_1125) );
AOI21xp5_ASAP7_75t_L g1260 ( .A1(n_464), .A2(n_1261), .B(n_1264), .Y(n_1260) );
AOI21xp5_ASAP7_75t_L g1307 ( .A1(n_464), .A2(n_1308), .B(n_1309), .Y(n_1307) );
AOI21xp5_ASAP7_75t_L g1324 ( .A1(n_464), .A2(n_1325), .B(n_1326), .Y(n_1324) );
AOI21xp5_ASAP7_75t_L g1561 ( .A1(n_464), .A2(n_1562), .B(n_1563), .Y(n_1561) );
AOI221xp5_ASAP7_75t_L g1824 ( .A1(n_464), .A2(n_736), .B1(n_1807), .B2(n_1825), .C(n_1826), .Y(n_1824) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B1(n_469), .B2(n_470), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_467), .B(n_740), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_467), .A2(n_471), .B1(n_859), .B2(n_860), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_467), .A2(n_471), .B1(n_910), .B2(n_911), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_467), .A2(n_470), .B1(n_1003), .B2(n_1004), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_467), .A2(n_471), .B1(n_1076), .B2(n_1077), .Y(n_1075) );
INVx1_ASAP7_75t_L g1173 ( .A(n_467), .Y(n_1173) );
HB1xp67_ASAP7_75t_L g1221 ( .A(n_467), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g1310 ( .A1(n_467), .A2(n_471), .B1(n_1311), .B2(n_1312), .Y(n_1310) );
AOI22xp5_ASAP7_75t_L g1828 ( .A1(n_467), .A2(n_471), .B1(n_1829), .B2(n_1830), .Y(n_1828) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g807 ( .A(n_468), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g1327 ( .A1(n_468), .A2(n_471), .B1(n_1328), .B2(n_1329), .Y(n_1327) );
AND2x4_ASAP7_75t_L g1414 ( .A(n_468), .B(n_1392), .Y(n_1414) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_470), .A2(n_805), .B1(n_806), .B2(n_808), .Y(n_804) );
AOI22xp5_ASAP7_75t_L g972 ( .A1(n_470), .A2(n_806), .B1(n_973), .B2(n_974), .Y(n_972) );
INVxp67_ASAP7_75t_SL g1166 ( .A(n_470), .Y(n_1166) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_470), .A2(n_1220), .B1(n_1221), .B2(n_1222), .Y(n_1219) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_471), .A2(n_734), .B1(n_735), .B2(n_736), .Y(n_733) );
HB1xp67_ASAP7_75t_L g1135 ( .A(n_471), .Y(n_1135) );
INVx1_ASAP7_75t_L g1269 ( .A(n_471), .Y(n_1269) );
AOI22xp33_ASAP7_75t_L g1560 ( .A1(n_471), .A2(n_806), .B1(n_1556), .B2(n_1557), .Y(n_1560) );
OAI21xp5_ASAP7_75t_L g714 ( .A1(n_472), .A2(n_715), .B(n_725), .Y(n_714) );
OAI21xp5_ASAP7_75t_SL g788 ( .A1(n_472), .A2(n_789), .B(n_797), .Y(n_788) );
OAI21xp5_ASAP7_75t_L g1069 ( .A1(n_472), .A2(n_1070), .B(n_1078), .Y(n_1069) );
AOI21xp5_ASAP7_75t_L g1217 ( .A1(n_472), .A2(n_1218), .B(n_1237), .Y(n_1217) );
OAI21xp5_ASAP7_75t_L g1305 ( .A1(n_472), .A2(n_1306), .B(n_1313), .Y(n_1305) );
OAI21xp5_ASAP7_75t_L g1558 ( .A1(n_472), .A2(n_1559), .B(n_1565), .Y(n_1558) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g837 ( .A(n_473), .Y(n_837) );
BUFx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g1020 ( .A(n_474), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1487 ( .A(n_474), .B(n_1488), .Y(n_1487) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OR2x6_ASAP7_75t_L g555 ( .A(n_475), .B(n_556), .Y(n_555) );
AND2x4_ASAP7_75t_L g615 ( .A(n_475), .B(n_616), .Y(n_615) );
BUFx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g538 ( .A(n_476), .Y(n_538) );
AOI21xp33_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_496), .B(n_497), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_478), .A2(n_810), .B(n_811), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_478), .B(n_835), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_478), .B(n_937), .Y(n_936) );
AOI21xp33_ASAP7_75t_SL g961 ( .A1(n_478), .A2(n_962), .B(n_963), .Y(n_961) );
AOI21xp33_ASAP7_75t_L g997 ( .A1(n_478), .A2(n_998), .B(n_999), .Y(n_997) );
NAND2xp33_ASAP7_75t_L g1061 ( .A(n_478), .B(n_1062), .Y(n_1061) );
AOI21xp33_ASAP7_75t_L g1140 ( .A1(n_478), .A2(n_1141), .B(n_1142), .Y(n_1140) );
AOI221xp5_ASAP7_75t_L g1200 ( .A1(n_478), .A2(n_866), .B1(n_1201), .B2(n_1202), .C(n_1203), .Y(n_1200) );
AOI21xp5_ASAP7_75t_L g1255 ( .A1(n_478), .A2(n_1256), .B(n_1257), .Y(n_1255) );
AOI21xp5_ASAP7_75t_L g1284 ( .A1(n_478), .A2(n_1285), .B(n_1286), .Y(n_1284) );
AOI21xp5_ASAP7_75t_L g1348 ( .A1(n_478), .A2(n_1349), .B(n_1350), .Y(n_1348) );
AOI211x1_ASAP7_75t_L g1537 ( .A1(n_478), .A2(n_1538), .B(n_1539), .C(n_1554), .Y(n_1537) );
INVx8_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_492), .Y(n_479) );
INVx1_ASAP7_75t_L g1399 ( .A(n_480), .Y(n_1399) );
OR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_486), .Y(n_480) );
INVx1_ASAP7_75t_L g751 ( .A(n_481), .Y(n_751) );
BUFx3_ASAP7_75t_L g764 ( .A(n_481), .Y(n_764) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_482), .Y(n_594) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx2_ASAP7_75t_L g703 ( .A(n_483), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_484), .Y(n_503) );
INVx2_ASAP7_75t_L g512 ( .A(n_484), .Y(n_512) );
AND2x4_ASAP7_75t_L g544 ( .A(n_484), .B(n_534), .Y(n_544) );
OR2x2_ASAP7_75t_L g566 ( .A(n_484), .B(n_514), .Y(n_566) );
INVx1_ASAP7_75t_L g502 ( .A(n_485), .Y(n_502) );
INVx2_ASAP7_75t_L g534 ( .A(n_485), .Y(n_534) );
OR2x2_ASAP7_75t_L g499 ( .A(n_486), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g568 ( .A(n_486), .Y(n_568) );
INVx1_ASAP7_75t_L g783 ( .A(n_486), .Y(n_783) );
OR2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_490), .Y(n_486) );
OR2x2_ASAP7_75t_L g579 ( .A(n_487), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g644 ( .A(n_487), .Y(n_644) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_487), .Y(n_708) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g508 ( .A(n_488), .Y(n_508) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g1420 ( .A(n_490), .Y(n_1420) );
INVx3_ASAP7_75t_L g517 ( .A(n_491), .Y(n_517) );
BUFx3_ASAP7_75t_L g537 ( .A(n_491), .Y(n_537) );
NAND2xp33_ASAP7_75t_SL g580 ( .A(n_491), .B(n_519), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g1486 ( .A(n_492), .B(n_1487), .Y(n_1486) );
OR2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_495), .Y(n_492) );
AND2x4_ASAP7_75t_L g525 ( .A(n_493), .B(n_516), .Y(n_525) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g608 ( .A(n_494), .Y(n_608) );
INVx1_ASAP7_75t_SL g1806 ( .A(n_498), .Y(n_1806) );
AND2x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_504), .Y(n_498) );
AND2x4_ASAP7_75t_L g743 ( .A(n_499), .B(n_504), .Y(n_743) );
INVx2_ASAP7_75t_L g1396 ( .A(n_499), .Y(n_1396) );
INVx3_ASAP7_75t_L g587 ( .A(n_500), .Y(n_587) );
INVx4_ASAP7_75t_L g758 ( .A(n_500), .Y(n_758) );
BUFx6f_ASAP7_75t_L g1868 ( .A(n_500), .Y(n_1868) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx3_ASAP7_75t_L g602 ( .A(n_501), .Y(n_602) );
BUFx2_ASAP7_75t_L g770 ( .A(n_501), .Y(n_770) );
NAND2x1p5_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
BUFx2_ASAP7_75t_L g695 ( .A(n_502), .Y(n_695) );
INVx2_ASAP7_75t_L g527 ( .A(n_503), .Y(n_527) );
AND2x4_ASAP7_75t_L g551 ( .A(n_503), .B(n_533), .Y(n_551) );
BUFx2_ASAP7_75t_L g692 ( .A(n_503), .Y(n_692) );
OR2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_508), .Y(n_504) );
OR2x2_ASAP7_75t_L g1457 ( .A(n_505), .B(n_508), .Y(n_1457) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVxp67_ASAP7_75t_L g520 ( .A(n_508), .Y(n_520) );
INVx1_ASAP7_75t_L g674 ( .A(n_508), .Y(n_674) );
INVx1_ASAP7_75t_L g1392 ( .A(n_508), .Y(n_1392) );
INVx5_ASAP7_75t_L g780 ( .A(n_509), .Y(n_780) );
INVx3_ASAP7_75t_L g866 ( .A(n_509), .Y(n_866) );
OR2x6_ASAP7_75t_L g509 ( .A(n_510), .B(n_520), .Y(n_509) );
OR2x2_ASAP7_75t_L g964 ( .A(n_510), .B(n_520), .Y(n_964) );
NAND2x1p5_ASAP7_75t_L g510 ( .A(n_511), .B(n_516), .Y(n_510) );
BUFx3_ASAP7_75t_L g542 ( .A(n_511), .Y(n_542) );
INVx8_ASAP7_75t_L g560 ( .A(n_511), .Y(n_560) );
BUFx3_ASAP7_75t_L g1035 ( .A(n_511), .Y(n_1035) );
HB1xp67_ASAP7_75t_L g1528 ( .A(n_511), .Y(n_1528) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
AND2x4_ASAP7_75t_L g548 ( .A(n_512), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVxp67_ASAP7_75t_L g549 ( .A(n_515), .Y(n_549) );
INVx1_ASAP7_75t_L g1439 ( .A(n_516), .Y(n_1439) );
AND2x6_ASAP7_75t_L g1446 ( .A(n_516), .B(n_526), .Y(n_1446) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_516), .B(n_532), .Y(n_1448) );
AND2x4_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g556 ( .A(n_517), .B(n_557), .Y(n_556) );
NAND3x1_ASAP7_75t_L g607 ( .A(n_517), .B(n_557), .C(n_608), .Y(n_607) );
OR2x4_ASAP7_75t_L g679 ( .A(n_517), .B(n_566), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_517), .Y(n_682) );
AND2x4_ASAP7_75t_L g687 ( .A(n_517), .B(n_544), .Y(n_687) );
OR2x6_ASAP7_75t_L g702 ( .A(n_517), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND3x4_ASAP7_75t_L g536 ( .A(n_519), .B(n_537), .C(n_538), .Y(n_536) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_519), .Y(n_706) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_519), .B(n_537), .Y(n_1429) );
NOR3xp33_ASAP7_75t_L g521 ( .A(n_522), .B(n_562), .C(n_571), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_535), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_524), .A2(n_529), .B1(n_791), .B2(n_815), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_524), .A2(n_529), .B1(n_840), .B2(n_842), .Y(n_868) );
AOI221xp5_ASAP7_75t_L g1386 ( .A1(n_524), .A2(n_529), .B1(n_572), .B2(n_1370), .C(n_1387), .Y(n_1386) );
AND2x4_ASAP7_75t_SL g524 ( .A(n_525), .B(n_526), .Y(n_524) );
AND2x4_ASAP7_75t_SL g529 ( .A(n_525), .B(n_530), .Y(n_529) );
AND2x4_ASAP7_75t_L g572 ( .A(n_525), .B(n_543), .Y(n_572) );
NAND2x1_ASAP7_75t_L g776 ( .A(n_525), .B(n_526), .Y(n_776) );
AND2x4_ASAP7_75t_L g778 ( .A(n_525), .B(n_530), .Y(n_778) );
AND2x2_ASAP7_75t_L g905 ( .A(n_525), .B(n_526), .Y(n_905) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_525), .B(n_526), .Y(n_1039) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g1304 ( .A(n_529), .Y(n_1304) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AOI33xp33_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_539), .A3(n_545), .B1(n_552), .B2(n_554), .B3(n_558), .Y(n_535) );
AOI33xp33_ASAP7_75t_L g816 ( .A1(n_536), .A2(n_554), .A3(n_817), .B1(n_819), .B2(n_820), .B3(n_821), .Y(n_816) );
AOI33xp33_ASAP7_75t_L g869 ( .A1(n_536), .A2(n_554), .A3(n_870), .B1(n_872), .B2(n_873), .B3(n_876), .Y(n_869) );
BUFx3_ASAP7_75t_L g890 ( .A(n_536), .Y(n_890) );
AOI33xp33_ASAP7_75t_L g946 ( .A1(n_536), .A2(n_947), .A3(n_949), .B1(n_954), .B2(n_955), .B3(n_957), .Y(n_946) );
AOI33xp33_ASAP7_75t_L g1026 ( .A1(n_536), .A2(n_894), .A3(n_1027), .B1(n_1029), .B2(n_1032), .B3(n_1033), .Y(n_1026) );
AOI33xp33_ASAP7_75t_L g1053 ( .A1(n_536), .A2(n_605), .A3(n_1054), .B1(n_1055), .B2(n_1059), .B3(n_1060), .Y(n_1053) );
AOI33xp33_ASAP7_75t_L g1379 ( .A1(n_536), .A2(n_1380), .A3(n_1381), .B1(n_1382), .B2(n_1384), .B3(n_1385), .Y(n_1379) );
INVx3_ASAP7_75t_L g691 ( .A(n_537), .Y(n_691) );
INVx2_ASAP7_75t_SL g933 ( .A(n_538), .Y(n_933) );
INVx1_ASAP7_75t_L g1139 ( .A(n_538), .Y(n_1139) );
OAI31xp33_ASAP7_75t_L g1416 ( .A1(n_538), .A2(n_1417), .A3(n_1421), .B(n_1440), .Y(n_1416) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
BUFx3_ASAP7_75t_L g818 ( .A(n_542), .Y(n_818) );
BUFx2_ASAP7_75t_L g892 ( .A(n_543), .Y(n_892) );
BUFx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx2_ASAP7_75t_L g561 ( .A(n_544), .Y(n_561) );
INVx2_ASAP7_75t_L g878 ( .A(n_544), .Y(n_878) );
BUFx3_ASAP7_75t_L g948 ( .A(n_544), .Y(n_948) );
BUFx2_ASAP7_75t_L g956 ( .A(n_544), .Y(n_956) );
BUFx2_ASAP7_75t_L g1028 ( .A(n_544), .Y(n_1028) );
BUFx2_ASAP7_75t_L g1296 ( .A(n_544), .Y(n_1296) );
AND2x2_ASAP7_75t_L g570 ( .A(n_546), .B(n_568), .Y(n_570) );
INVx2_ASAP7_75t_L g1816 ( .A(n_546), .Y(n_1816) );
INVx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx2_ASAP7_75t_L g1251 ( .A(n_547), .Y(n_1251) );
OAI221xp5_ASAP7_75t_L g1289 ( .A1(n_547), .A2(n_1290), .B1(n_1291), .B2(n_1294), .C(n_1295), .Y(n_1289) );
OR2x6_ASAP7_75t_SL g1418 ( .A(n_547), .B(n_1419), .Y(n_1418) );
BUFx2_ASAP7_75t_L g1861 ( .A(n_547), .Y(n_1861) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx8_ASAP7_75t_L g553 ( .A(n_548), .Y(n_553) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_548), .Y(n_591) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_548), .Y(n_599) );
BUFx2_ASAP7_75t_L g899 ( .A(n_550), .Y(n_899) );
BUFx12f_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx3_ASAP7_75t_L g822 ( .A(n_551), .Y(n_822) );
INVx5_ASAP7_75t_L g953 ( .A(n_551), .Y(n_953) );
BUFx3_ASAP7_75t_L g1031 ( .A(n_551), .Y(n_1031) );
BUFx2_ASAP7_75t_L g1058 ( .A(n_551), .Y(n_1058) );
AND2x4_ASAP7_75t_L g1488 ( .A(n_551), .B(n_1420), .Y(n_1488) );
INVx3_ASAP7_75t_L g748 ( .A(n_553), .Y(n_748) );
AND2x4_ASAP7_75t_L g782 ( .A(n_553), .B(n_783), .Y(n_782) );
HB1xp67_ASAP7_75t_L g888 ( .A(n_553), .Y(n_888) );
INVx2_ASAP7_75t_SL g1111 ( .A(n_553), .Y(n_1111) );
INVx2_ASAP7_75t_SL g1339 ( .A(n_553), .Y(n_1339) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g1385 ( .A(n_555), .Y(n_1385) );
OAI33xp33_ASAP7_75t_L g1851 ( .A1(n_555), .A2(n_1180), .A3(n_1852), .B1(n_1859), .B2(n_1863), .B3(n_1866), .Y(n_1851) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g864 ( .A(n_560), .Y(n_864) );
INVx8_ASAP7_75t_L g871 ( .A(n_560), .Y(n_871) );
INVx2_ASAP7_75t_L g1189 ( .A(n_560), .Y(n_1189) );
INVx1_ASAP7_75t_L g897 ( .A(n_561), .Y(n_897) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_567), .Y(n_563) );
OR2x6_ASAP7_75t_L g772 ( .A(n_564), .B(n_567), .Y(n_772) );
INVx2_ASAP7_75t_SL g1106 ( .A(n_564), .Y(n_1106) );
INVx2_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
INVx3_ASAP7_75t_L g1855 ( .A(n_565), .Y(n_1855) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
BUFx4f_ASAP7_75t_L g584 ( .A(n_566), .Y(n_584) );
OR2x4_ASAP7_75t_L g700 ( .A(n_566), .B(n_682), .Y(n_700) );
BUFx3_ASAP7_75t_L g754 ( .A(n_566), .Y(n_754) );
BUFx3_ASAP7_75t_L g767 ( .A(n_566), .Y(n_767) );
INVxp67_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2x1_ASAP7_75t_L g1389 ( .A(n_569), .B(n_1390), .Y(n_1389) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_570), .A2(n_859), .B1(n_860), .B2(n_863), .Y(n_862) );
NOR3xp33_ASAP7_75t_L g1287 ( .A(n_571), .B(n_1288), .C(n_1303), .Y(n_1287) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx3_ASAP7_75t_L g784 ( .A(n_572), .Y(n_784) );
NOR3xp33_ASAP7_75t_L g812 ( .A(n_572), .B(n_813), .C(n_823), .Y(n_812) );
AOI211xp5_ASAP7_75t_L g865 ( .A1(n_572), .A2(n_850), .B(n_866), .C(n_867), .Y(n_865) );
INVx3_ASAP7_75t_L g1022 ( .A(n_572), .Y(n_1022) );
NOR3xp33_ASAP7_75t_L g1336 ( .A(n_572), .B(n_1337), .C(n_1347), .Y(n_1336) );
NOR3xp33_ASAP7_75t_SL g1808 ( .A(n_572), .B(n_1809), .C(n_1820), .Y(n_1808) );
NAND3xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_645), .C(n_675), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_613), .Y(n_575) );
OAI33xp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_581), .A3(n_588), .B1(n_595), .B2(n_604), .B3(n_609), .Y(n_576) );
BUFx3_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI22xp5_ASAP7_75t_SL g1288 ( .A1(n_578), .A2(n_1289), .B1(n_1297), .B2(n_1298), .Y(n_1288) );
BUFx4f_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx8_ASAP7_75t_L g752 ( .A(n_579), .Y(n_752) );
BUFx2_ASAP7_75t_L g1180 ( .A(n_579), .Y(n_1180) );
BUFx4f_ASAP7_75t_L g1810 ( .A(n_579), .Y(n_1810) );
OAI22xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_583), .B1(n_585), .B2(n_586), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_582), .A2(n_610), .B1(n_618), .B2(n_622), .Y(n_617) );
OAI22xp33_ASAP7_75t_L g609 ( .A1(n_583), .A2(n_610), .B1(n_611), .B2(n_612), .Y(n_609) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g1183 ( .A(n_584), .Y(n_1183) );
OAI22xp5_ASAP7_75t_L g1422 ( .A1(n_584), .A2(n_611), .B1(n_1423), .B2(n_1424), .Y(n_1422) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_585), .A2(n_612), .B1(n_622), .B2(n_629), .Y(n_634) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g1102 ( .A(n_587), .Y(n_1102) );
INVx3_ASAP7_75t_L g1435 ( .A(n_587), .Y(n_1435) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B1(n_592), .B2(n_593), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_589), .A2(n_600), .B1(n_629), .B2(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g1030 ( .A(n_590), .Y(n_1030) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x4_ASAP7_75t_L g681 ( .A(n_591), .B(n_682), .Y(n_681) );
BUFx6f_ASAP7_75t_L g762 ( .A(n_591), .Y(n_762) );
INVx2_ASAP7_75t_L g875 ( .A(n_591), .Y(n_875) );
INVx2_ASAP7_75t_L g951 ( .A(n_591), .Y(n_951) );
BUFx6f_ASAP7_75t_L g1383 ( .A(n_591), .Y(n_1383) );
OAI22xp33_ASAP7_75t_L g635 ( .A1(n_592), .A2(n_603), .B1(n_636), .B2(n_639), .Y(n_635) );
OAI22xp33_ASAP7_75t_L g1100 ( .A1(n_593), .A2(n_1101), .B1(n_1102), .B2(n_1103), .Y(n_1100) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_593), .A2(n_1111), .B1(n_1112), .B2(n_1113), .Y(n_1110) );
OAI22xp5_ASAP7_75t_L g1430 ( .A1(n_593), .A2(n_1431), .B1(n_1432), .B2(n_1433), .Y(n_1430) );
INVx3_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx3_ASAP7_75t_L g611 ( .A(n_594), .Y(n_611) );
INVx3_ASAP7_75t_L g1179 ( .A(n_594), .Y(n_1179) );
CKINVDCx8_ASAP7_75t_R g1300 ( .A(n_594), .Y(n_1300) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_600), .B1(n_601), .B2(n_603), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx8_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
BUFx3_ASAP7_75t_L g1108 ( .A(n_598), .Y(n_1108) );
OAI221xp5_ASAP7_75t_L g1525 ( .A1(n_598), .A2(n_764), .B1(n_1511), .B2(n_1526), .C(n_1527), .Y(n_1525) );
INVx5_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_SL g1057 ( .A(n_599), .Y(n_1057) );
INVx3_ASAP7_75t_L g1427 ( .A(n_599), .Y(n_1427) );
INVx2_ASAP7_75t_SL g1431 ( .A(n_599), .Y(n_1431) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g685 ( .A(n_602), .Y(n_685) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
BUFx2_ASAP7_75t_L g894 ( .A(n_606), .Y(n_894) );
BUFx2_ASAP7_75t_L g957 ( .A(n_606), .Y(n_957) );
BUFx2_ASAP7_75t_L g1552 ( .A(n_606), .Y(n_1552) );
INVx3_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx3_ASAP7_75t_L g1212 ( .A(n_607), .Y(n_1212) );
OAI33xp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_617), .A3(n_628), .B1(n_634), .B2(n_635), .B3(n_640), .Y(n_613) );
INVx2_ASAP7_75t_SL g1872 ( .A(n_614), .Y(n_1872) );
INVx4_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g1452 ( .A(n_615), .B(n_1453), .Y(n_1452) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
INVx3_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
BUFx6f_ASAP7_75t_L g1273 ( .A(n_621), .Y(n_1273) );
INVx4_ASAP7_75t_L g1499 ( .A(n_621), .Y(n_1499) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OAI22xp33_ASAP7_75t_L g1873 ( .A1(n_624), .A2(n_636), .B1(n_1853), .B2(n_1867), .Y(n_1873) );
INVx4_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_SL g984 ( .A(n_625), .Y(n_984) );
INVx2_ASAP7_75t_L g1016 ( .A(n_625), .Y(n_1016) );
INVx1_ASAP7_75t_L g1275 ( .A(n_625), .Y(n_1275) );
BUFx6f_ASAP7_75t_L g1577 ( .A(n_625), .Y(n_1577) );
INVx1_ASAP7_75t_L g1836 ( .A(n_625), .Y(n_1836) );
INVx8_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g667 ( .A(n_626), .B(n_653), .Y(n_667) );
BUFx2_ASAP7_75t_L g1169 ( .A(n_626), .Y(n_1169) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g1874 ( .A1(n_629), .A2(n_1860), .B1(n_1864), .B2(n_1875), .Y(n_1874) );
OAI22xp5_ASAP7_75t_L g1876 ( .A1(n_629), .A2(n_1856), .B1(n_1869), .B2(n_1875), .Y(n_1876) );
BUFx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g1473 ( .A(n_630), .Y(n_1473) );
BUFx2_ASAP7_75t_L g1571 ( .A(n_630), .Y(n_1571) );
OAI211xp5_ASAP7_75t_L g1331 ( .A1(n_631), .A2(n_1332), .B(n_1333), .C(n_1334), .Y(n_1331) );
OAI211xp5_ASAP7_75t_L g1510 ( .A1(n_631), .A2(n_1511), .B(n_1512), .C(n_1513), .Y(n_1510) );
INVx5_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx2_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
BUFx2_ASAP7_75t_SL g639 ( .A(n_633), .Y(n_639) );
OR2x2_ASAP7_75t_L g1466 ( .A(n_633), .B(n_1467), .Y(n_1466) );
BUFx3_ASAP7_75t_L g1875 ( .A(n_633), .Y(n_1875) );
OAI221xp5_ASAP7_75t_L g1012 ( .A1(n_636), .A2(n_1013), .B1(n_1014), .B2(n_1017), .C(n_1018), .Y(n_1012) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
BUFx6f_ASAP7_75t_L g981 ( .A(n_638), .Y(n_981) );
BUFx3_ASAP7_75t_L g1833 ( .A(n_638), .Y(n_1833) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI31xp33_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_658), .A3(n_668), .B(n_672), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx3_ASAP7_75t_L g1882 ( .A(n_648), .Y(n_1882) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_654), .B1(n_655), .B2(n_656), .Y(n_650) );
BUFx3_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_654), .A2(n_689), .B1(n_693), .B2(n_696), .Y(n_688) );
BUFx3_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g1887 ( .A(n_657), .Y(n_1887) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx3_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
INVx4_ASAP7_75t_L g1892 ( .A(n_671), .Y(n_1892) );
BUFx3_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI31xp33_ASAP7_75t_L g1880 ( .A1(n_673), .A2(n_1881), .A3(n_1889), .B(n_1890), .Y(n_1880) );
OAI31xp33_ASAP7_75t_SL g675 ( .A1(n_676), .A2(n_683), .A3(n_697), .B(n_704), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g1895 ( .A(n_681), .Y(n_1895) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
CKINVDCx8_ASAP7_75t_R g686 ( .A(n_687), .Y(n_686) );
CKINVDCx8_ASAP7_75t_R g1899 ( .A(n_687), .Y(n_1899) );
BUFx3_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
AND2x4_ASAP7_75t_L g694 ( .A(n_691), .B(n_695), .Y(n_694) );
AND2x4_ASAP7_75t_L g1901 ( .A(n_691), .B(n_692), .Y(n_1901) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g1900 ( .A1(n_694), .A2(n_1885), .B1(n_1901), .B2(n_1902), .Y(n_1900) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g1904 ( .A(n_699), .Y(n_1904) );
INVx2_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
BUFx3_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g1906 ( .A(n_702), .Y(n_1906) );
BUFx3_ASAP7_75t_L g1187 ( .A(n_703), .Y(n_1187) );
INVx1_ASAP7_75t_L g1293 ( .A(n_703), .Y(n_1293) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_707), .Y(n_704) );
AND2x2_ASAP7_75t_L g1907 ( .A(n_705), .B(n_707), .Y(n_1907) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g828 ( .A(n_709), .Y(n_828) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_711), .B1(n_786), .B2(n_826), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NOR3xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_773), .C(n_785), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_741), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_721), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g928 ( .A(n_720), .Y(n_928) );
NAND3xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_733), .C(n_739), .Y(n_725) );
INVx2_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_732), .A2(n_775), .B1(n_777), .B2(n_778), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_734), .B(n_782), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_735), .B(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g1361 ( .A(n_736), .Y(n_1361) );
AND2x4_ASAP7_75t_L g1482 ( .A(n_737), .B(n_1483), .Y(n_1482) );
INVx3_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g926 ( .A(n_738), .Y(n_926) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_744), .B(n_745), .Y(n_741) );
AOI21xp5_ASAP7_75t_L g1066 ( .A1(n_742), .A2(n_1067), .B(n_1068), .Y(n_1066) );
AOI21xp5_ASAP7_75t_SL g1174 ( .A1(n_742), .A2(n_1175), .B(n_1176), .Y(n_1174) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
HB1xp67_ASAP7_75t_L g1143 ( .A(n_743), .Y(n_1143) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_748), .B1(n_749), .B2(n_750), .Y(n_746) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
OAI33xp33_ASAP7_75t_L g1099 ( .A1(n_752), .A2(n_1100), .A3(n_1104), .B1(n_1110), .B2(n_1114), .B3(n_1117), .Y(n_1099) );
OAI22xp5_ASAP7_75t_SL g1337 ( .A1(n_752), .A2(n_1211), .B1(n_1338), .B2(n_1343), .Y(n_1337) );
OAI22xp33_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_755), .B1(n_756), .B2(n_757), .Y(n_753) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g1898 ( .A(n_758), .Y(n_1898) );
OAI22xp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_761), .B1(n_763), .B2(n_764), .Y(n_759) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g1863 ( .A1(n_764), .A2(n_1861), .B1(n_1864), .B2(n_1865), .Y(n_1863) );
OAI22xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_767), .B1(n_768), .B2(n_771), .Y(n_765) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
OAI221xp5_ASAP7_75t_L g1425 ( .A1(n_770), .A2(n_1426), .B1(n_1427), .B2(n_1428), .C(n_1429), .Y(n_1425) );
OR2x6_ASAP7_75t_L g1438 ( .A(n_770), .B(n_1439), .Y(n_1438) );
INVx1_ASAP7_75t_L g1858 ( .A(n_770), .Y(n_1858) );
NAND2xp5_ASAP7_75t_L g1531 ( .A(n_772), .B(n_1532), .Y(n_1531) );
NAND4xp25_ASAP7_75t_L g773 ( .A(n_774), .B(n_779), .C(n_781), .D(n_784), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_775), .A2(n_778), .B1(n_944), .B2(n_945), .Y(n_943) );
AOI22xp5_ASAP7_75t_L g1048 ( .A1(n_775), .A2(n_778), .B1(n_1049), .B2(n_1050), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g1214 ( .A1(n_775), .A2(n_778), .B1(n_1215), .B2(n_1216), .Y(n_1214) );
AOI221x1_ASAP7_75t_L g1518 ( .A1(n_775), .A2(n_778), .B1(n_1496), .B2(n_1502), .C(n_1519), .Y(n_1518) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_778), .A2(n_904), .B1(n_905), .B2(n_906), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_778), .A2(n_1038), .B1(n_1039), .B2(n_1040), .Y(n_1037) );
HB1xp67_ASAP7_75t_L g1097 ( .A(n_778), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g1149 ( .A1(n_778), .A2(n_905), .B1(n_1150), .B2(n_1151), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_778), .A2(n_905), .B1(n_1245), .B2(n_1246), .Y(n_1244) );
AO22x1_ASAP7_75t_L g1541 ( .A1(n_778), .A2(n_905), .B1(n_1542), .B2(n_1543), .Y(n_1541) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_780), .B(n_1052), .Y(n_1051) );
NAND2xp5_ASAP7_75t_L g1533 ( .A(n_780), .B(n_1534), .Y(n_1533) );
NAND2xp5_ASAP7_75t_L g1545 ( .A(n_780), .B(n_1546), .Y(n_1545) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_782), .A2(n_863), .B1(n_910), .B2(n_911), .Y(n_935) );
INVx2_ASAP7_75t_L g959 ( .A(n_782), .Y(n_959) );
INVx2_ASAP7_75t_L g1025 ( .A(n_782), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g1238 ( .A1(n_782), .A2(n_863), .B1(n_1220), .B2(n_1222), .Y(n_1238) );
AOI22xp33_ASAP7_75t_L g1318 ( .A1(n_782), .A2(n_863), .B1(n_1311), .B2(n_1312), .Y(n_1318) );
AOI22xp33_ASAP7_75t_L g1351 ( .A1(n_782), .A2(n_863), .B1(n_1328), .B2(n_1329), .Y(n_1351) );
AOI22xp33_ASAP7_75t_L g1555 ( .A1(n_782), .A2(n_863), .B1(n_1556), .B2(n_1557), .Y(n_1555) );
AND2x4_ASAP7_75t_L g863 ( .A(n_783), .B(n_864), .Y(n_863) );
AND2x4_ASAP7_75t_L g1397 ( .A(n_783), .B(n_864), .Y(n_1397) );
NAND3xp33_ASAP7_75t_L g900 ( .A(n_784), .B(n_901), .C(n_903), .Y(n_900) );
INVx1_ASAP7_75t_L g960 ( .A(n_784), .Y(n_960) );
NAND4xp25_ASAP7_75t_SL g1047 ( .A(n_784), .B(n_1048), .C(n_1051), .D(n_1053), .Y(n_1047) );
NAND2xp5_ASAP7_75t_SL g1544 ( .A(n_784), .B(n_1545), .Y(n_1544) );
INVx1_ASAP7_75t_L g826 ( .A(n_786), .Y(n_826) );
INVx1_ASAP7_75t_L g825 ( .A(n_787), .Y(n_825) );
NAND3xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_809), .C(n_812), .Y(n_787) );
HB1xp67_ASAP7_75t_SL g1128 ( .A(n_802), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_806), .A2(n_1133), .B1(n_1134), .B2(n_1135), .Y(n_1132) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_814), .B(n_816), .Y(n_813) );
XNOR2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_880), .Y(n_829) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
NAND3xp33_ASAP7_75t_L g833 ( .A(n_834), .B(n_836), .C(n_865), .Y(n_833) );
AOI21xp5_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_838), .B(n_861), .Y(n_836) );
OAI21xp5_ASAP7_75t_L g1822 ( .A1(n_837), .A2(n_1823), .B(n_1831), .Y(n_1822) );
NAND3xp33_ASAP7_75t_L g838 ( .A(n_839), .B(n_849), .C(n_858), .Y(n_838) );
INVx1_ASAP7_75t_L g931 ( .A(n_841), .Y(n_931) );
AOI222xp33_ASAP7_75t_L g1228 ( .A1(n_841), .A2(n_1215), .B1(n_1216), .B2(n_1229), .C1(n_1230), .C2(n_1236), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1495 ( .A(n_841), .B(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx2_ASAP7_75t_L g918 ( .A(n_845), .Y(n_918) );
INVx1_ASAP7_75t_L g1278 ( .A(n_845), .Y(n_1278) );
BUFx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g1233 ( .A(n_846), .Y(n_1233) );
INVx1_ASAP7_75t_L g1235 ( .A(n_853), .Y(n_1235) );
INVx2_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx2_ASAP7_75t_L g923 ( .A(n_854), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_863), .B(n_1156), .Y(n_1155) );
AOI22xp5_ASAP7_75t_L g1839 ( .A1(n_863), .A2(n_1829), .B1(n_1830), .B2(n_1840), .Y(n_1839) );
AOI22xp5_ASAP7_75t_L g1441 ( .A1(n_864), .A2(n_877), .B1(n_1413), .B2(n_1442), .Y(n_1441) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_866), .B(n_902), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_866), .B(n_1153), .Y(n_1152) );
AOI22xp5_ASAP7_75t_L g1804 ( .A1(n_866), .A2(n_1805), .B1(n_1806), .B2(n_1807), .Y(n_1804) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_868), .B(n_869), .Y(n_867) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
OAI221xp5_ASAP7_75t_L g1298 ( .A1(n_875), .A2(n_1299), .B1(n_1300), .B2(n_1301), .C(n_1302), .Y(n_1298) );
INVx2_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g1036 ( .A(n_878), .Y(n_1036) );
INVx1_ASAP7_75t_L g1190 ( .A(n_878), .Y(n_1190) );
INVx2_ASAP7_75t_L g1346 ( .A(n_878), .Y(n_1346) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_881), .A2(n_882), .B1(n_938), .B2(n_939), .Y(n_880) );
INVx2_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
XNOR2x1_ASAP7_75t_L g882 ( .A(n_883), .B(n_884), .Y(n_882) );
AND3x2_ASAP7_75t_L g884 ( .A(n_885), .B(n_907), .C(n_936), .Y(n_884) );
NOR2xp33_ASAP7_75t_SL g885 ( .A(n_886), .B(n_900), .Y(n_885) );
OAI21xp5_ASAP7_75t_SL g886 ( .A1(n_887), .A2(n_889), .B(n_893), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_890), .B(n_891), .Y(n_889) );
AOI33xp33_ASAP7_75t_L g1204 ( .A1(n_890), .A2(n_1205), .A3(n_1206), .B1(n_1209), .B2(n_1210), .B3(n_1213), .Y(n_1204) );
AOI33xp33_ASAP7_75t_L g1247 ( .A1(n_890), .A2(n_1210), .A3(n_1248), .B1(n_1249), .B2(n_1252), .B3(n_1253), .Y(n_1247) );
AOI33xp33_ASAP7_75t_L g1547 ( .A1(n_890), .A2(n_1548), .A3(n_1549), .B1(n_1551), .B2(n_1552), .B3(n_1553), .Y(n_1547) );
NAND3xp33_ASAP7_75t_L g893 ( .A(n_894), .B(n_895), .C(n_898), .Y(n_893) );
INVx1_ASAP7_75t_L g1117 ( .A(n_894), .Y(n_1117) );
INVx1_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
AOI21xp5_ASAP7_75t_SL g907 ( .A1(n_908), .A2(n_933), .B(n_934), .Y(n_907) );
NAND3xp33_ASAP7_75t_L g908 ( .A(n_909), .B(n_912), .C(n_920), .Y(n_908) );
INVx2_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
INVx2_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g988 ( .A(n_916), .Y(n_988) );
HB1xp67_ASAP7_75t_L g1127 ( .A(n_916), .Y(n_1127) );
INVx2_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx2_ASAP7_75t_L g1019 ( .A(n_917), .Y(n_1019) );
AOI31xp33_ASAP7_75t_L g920 ( .A1(n_921), .A2(n_924), .A3(n_927), .B(n_930), .Y(n_920) );
BUFx2_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g1236 ( .A(n_932), .Y(n_1236) );
OAI21xp5_ASAP7_75t_L g965 ( .A1(n_933), .A2(n_966), .B(n_975), .Y(n_965) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
NAND3xp33_ASAP7_75t_L g940 ( .A(n_941), .B(n_961), .C(n_965), .Y(n_940) );
NOR3xp33_ASAP7_75t_L g941 ( .A(n_942), .B(n_958), .C(n_960), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_943), .B(n_946), .Y(n_942) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
OAI22xp5_ASAP7_75t_L g1177 ( .A1(n_951), .A2(n_1161), .B1(n_1178), .B2(n_1179), .Y(n_1177) );
INVx2_ASAP7_75t_R g952 ( .A(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g1208 ( .A(n_953), .Y(n_1208) );
INVx2_ASAP7_75t_L g1550 ( .A(n_953), .Y(n_1550) );
INVxp67_ASAP7_75t_L g1840 ( .A(n_959), .Y(n_1840) );
NAND2xp5_ASAP7_75t_L g1480 ( .A(n_964), .B(n_1481), .Y(n_1480) );
INVx2_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
INVx2_ASAP7_75t_L g1011 ( .A(n_977), .Y(n_1011) );
NOR2x1_ASAP7_75t_L g977 ( .A(n_978), .B(n_979), .Y(n_977) );
INVx1_ASAP7_75t_L g1374 ( .A(n_979), .Y(n_1374) );
OAI221xp5_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_982), .B1(n_983), .B2(n_985), .C(n_986), .Y(n_980) );
OAI221xp5_ASAP7_75t_SL g1121 ( .A1(n_981), .A2(n_1014), .B1(n_1107), .B2(n_1115), .C(n_1122), .Y(n_1121) );
OAI221xp5_ASAP7_75t_L g1160 ( .A1(n_981), .A2(n_1161), .B1(n_1162), .B2(n_1163), .C(n_1164), .Y(n_1160) );
OAI221xp5_ASAP7_75t_L g1167 ( .A1(n_981), .A2(n_1168), .B1(n_1169), .B2(n_1170), .C(n_1171), .Y(n_1167) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
HB1xp67_ASAP7_75t_L g1162 ( .A(n_984), .Y(n_1162) );
INVx1_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
XNOR2xp5_ASAP7_75t_L g991 ( .A(n_992), .B(n_1145), .Y(n_991) );
XNOR2x1_ASAP7_75t_L g992 ( .A(n_993), .B(n_1091), .Y(n_992) );
OAI22x1_ASAP7_75t_L g993 ( .A1(n_994), .A2(n_1042), .B1(n_1043), .B2(n_1090), .Y(n_993) );
INVx2_ASAP7_75t_L g1090 ( .A(n_994), .Y(n_1090) );
AO21x2_ASAP7_75t_L g994 ( .A1(n_995), .A2(n_996), .B(n_1041), .Y(n_994) );
NAND3xp33_ASAP7_75t_SL g996 ( .A(n_997), .B(n_1000), .C(n_1021), .Y(n_996) );
OAI21xp5_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1009), .B(n_1020), .Y(n_1000) );
BUFx2_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
BUFx2_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
BUFx6f_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
OAI31xp33_ASAP7_75t_L g1158 ( .A1(n_1020), .A2(n_1159), .A3(n_1165), .B(n_1172), .Y(n_1158) );
AND4x1_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1023), .C(n_1026), .D(n_1037), .Y(n_1021) );
INVx2_ASAP7_75t_SL g1118 ( .A(n_1022), .Y(n_1118) );
NAND5xp2_ASAP7_75t_L g1148 ( .A(n_1022), .B(n_1149), .C(n_1152), .D(n_1154), .E(n_1155), .Y(n_1148) );
NAND3xp33_ASAP7_75t_SL g1203 ( .A(n_1022), .B(n_1204), .C(n_1214), .Y(n_1203) );
AND5x1_ASAP7_75t_L g1492 ( .A(n_1022), .B(n_1493), .C(n_1518), .D(n_1529), .E(n_1533), .Y(n_1492) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
BUFx2_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
INVx1_ASAP7_75t_L g1821 ( .A(n_1039), .Y(n_1821) );
INVx2_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
NAND2x1p5_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1063), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1061), .Y(n_1045) );
INVxp67_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
NOR2xp33_ASAP7_75t_SL g1087 ( .A(n_1047), .B(n_1088), .Y(n_1087) );
INVx2_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_1061), .B(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1069), .Y(n_1065) );
OAI211xp5_ASAP7_75t_L g1080 ( .A1(n_1081), .A2(n_1082), .B(n_1084), .C(n_1086), .Y(n_1080) );
INVx2_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1083), .Y(n_1315) );
INVx2_ASAP7_75t_L g1500 ( .A(n_1083), .Y(n_1500) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
AND3x2_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1119), .C(n_1140), .Y(n_1093) );
NOR4xp25_ASAP7_75t_L g1094 ( .A(n_1095), .B(n_1098), .C(n_1099), .D(n_1118), .Y(n_1094) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
OAI22xp33_ASAP7_75t_L g1114 ( .A1(n_1102), .A2(n_1105), .B1(n_1115), .B2(n_1116), .Y(n_1114) );
OAI22xp33_ASAP7_75t_L g1181 ( .A1(n_1102), .A2(n_1168), .B1(n_1182), .B2(n_1184), .Y(n_1181) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_1105), .A2(n_1107), .B1(n_1108), .B2(n_1109), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
OAI221xp5_ASAP7_75t_L g1185 ( .A1(n_1108), .A2(n_1163), .B1(n_1186), .B2(n_1187), .C(n_1188), .Y(n_1185) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1111), .Y(n_1207) );
NOR3xp33_ASAP7_75t_L g1242 ( .A(n_1118), .B(n_1243), .C(n_1254), .Y(n_1242) );
OAI21xp5_ASAP7_75t_L g1119 ( .A1(n_1120), .A2(n_1124), .B(n_1136), .Y(n_1119) );
INVx1_ASAP7_75t_SL g1130 ( .A(n_1131), .Y(n_1130) );
OAI21xp5_ASAP7_75t_L g1258 ( .A1(n_1136), .A2(n_1259), .B(n_1270), .Y(n_1258) );
INVx2_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
HB1xp67_ASAP7_75t_L g1514 ( .A(n_1138), .Y(n_1514) );
BUFx2_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
BUFx2_ASAP7_75t_L g1335 ( .A(n_1139), .Y(n_1335) );
AOI21x1_ASAP7_75t_L g1359 ( .A1(n_1139), .A2(n_1360), .B(n_1377), .Y(n_1359) );
INVx2_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
XNOR2x1_ASAP7_75t_L g1146 ( .A(n_1147), .B(n_1191), .Y(n_1146) );
NOR2x1_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1157), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1174), .Y(n_1157) );
OAI22xp5_ASAP7_75t_L g1878 ( .A1(n_1169), .A2(n_1862), .B1(n_1865), .B2(n_1879), .Y(n_1878) );
OAI221xp5_ASAP7_75t_L g1520 ( .A1(n_1179), .A2(n_1431), .B1(n_1521), .B2(n_1522), .C(n_1523), .Y(n_1520) );
OAI22xp5_ASAP7_75t_L g1859 ( .A1(n_1179), .A2(n_1860), .B1(n_1861), .B2(n_1862), .Y(n_1859) );
OAI22xp5_ASAP7_75t_SL g1519 ( .A1(n_1180), .A2(n_1520), .B1(n_1524), .B2(n_1525), .Y(n_1519) );
INVx2_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
OAI221xp5_ASAP7_75t_L g1815 ( .A1(n_1187), .A2(n_1816), .B1(n_1817), .B2(n_1818), .C(n_1819), .Y(n_1815) );
INVxp67_ASAP7_75t_SL g1193 ( .A(n_1194), .Y(n_1193) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
AO22x2_ASAP7_75t_L g1195 ( .A1(n_1196), .A2(n_1353), .B1(n_1354), .B2(n_1581), .Y(n_1195) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1196), .Y(n_1581) );
XNOR2xp5_ASAP7_75t_L g1196 ( .A(n_1197), .B(n_1280), .Y(n_1196) );
XOR2xp5_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1240), .Y(n_1197) );
XNOR2xp5_ASAP7_75t_L g1198 ( .A(n_1199), .B(n_1239), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1200), .B(n_1217), .Y(n_1199) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
CKINVDCx5p33_ASAP7_75t_R g1211 ( .A(n_1212), .Y(n_1211) );
INVx2_ASAP7_75t_L g1297 ( .A(n_1212), .Y(n_1297) );
INVx2_ASAP7_75t_L g1524 ( .A(n_1212), .Y(n_1524) );
NAND3xp33_ASAP7_75t_L g1218 ( .A(n_1219), .B(n_1223), .C(n_1228), .Y(n_1218) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_1221), .A2(n_1266), .B1(n_1267), .B2(n_1268), .Y(n_1265) );
INVx2_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
NAND3xp33_ASAP7_75t_L g1241 ( .A(n_1242), .B(n_1255), .C(n_1258), .Y(n_1241) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1247), .Y(n_1243) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
OAI221xp5_ASAP7_75t_L g1271 ( .A1(n_1272), .A2(n_1274), .B1(n_1275), .B2(n_1276), .C(n_1277), .Y(n_1271) );
OAI22xp5_ASAP7_75t_L g1573 ( .A1(n_1272), .A2(n_1574), .B1(n_1575), .B2(n_1576), .Y(n_1573) );
INVx2_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
BUFx3_ASAP7_75t_L g1280 ( .A(n_1281), .Y(n_1280) );
AO22x2_ASAP7_75t_L g1281 ( .A1(n_1282), .A2(n_1319), .B1(n_1320), .B2(n_1352), .Y(n_1281) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1282), .Y(n_1352) );
AND4x1_ASAP7_75t_L g1283 ( .A(n_1284), .B(n_1287), .C(n_1305), .D(n_1318), .Y(n_1283) );
OAI221xp5_ASAP7_75t_L g1338 ( .A1(n_1291), .A2(n_1339), .B1(n_1340), .B2(n_1341), .C(n_1342), .Y(n_1338) );
INVx3_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
BUFx2_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
OAI211xp5_ASAP7_75t_L g1314 ( .A1(n_1299), .A2(n_1315), .B(n_1316), .C(n_1317), .Y(n_1314) );
OAI221xp5_ASAP7_75t_L g1343 ( .A1(n_1300), .A2(n_1332), .B1(n_1339), .B2(n_1344), .C(n_1345), .Y(n_1343) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
AND4x1_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1336), .C(n_1348), .D(n_1351), .Y(n_1321) );
OAI21xp5_ASAP7_75t_L g1322 ( .A1(n_1323), .A2(n_1330), .B(n_1335), .Y(n_1322) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1354), .Y(n_1353) );
AO22x2_ASAP7_75t_L g1354 ( .A1(n_1355), .A2(n_1535), .B1(n_1579), .B2(n_1580), .Y(n_1354) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1355), .Y(n_1579) );
XNOR2xp5_ASAP7_75t_L g1355 ( .A(n_1356), .B(n_1491), .Y(n_1355) );
OAI22xp5_ASAP7_75t_L g1356 ( .A1(n_1357), .A2(n_1408), .B1(n_1489), .B2(n_1490), .Y(n_1356) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1357), .Y(n_1490) );
NAND3xp33_ASAP7_75t_L g1357 ( .A(n_1358), .B(n_1401), .C(n_1405), .Y(n_1357) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1359), .Y(n_1402) );
AOI22xp5_ASAP7_75t_L g1362 ( .A1(n_1363), .A2(n_1364), .B1(n_1365), .B2(n_1366), .Y(n_1362) );
AOI22xp5_ASAP7_75t_L g1367 ( .A1(n_1368), .A2(n_1374), .B1(n_1375), .B2(n_1376), .Y(n_1367) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
AOI222xp33_ASAP7_75t_L g1395 ( .A1(n_1373), .A2(n_1396), .B1(n_1397), .B2(n_1398), .C1(n_1399), .C2(n_1400), .Y(n_1395) );
AOI22xp5_ASAP7_75t_L g1497 ( .A1(n_1374), .A2(n_1375), .B1(n_1498), .B2(n_1504), .Y(n_1497) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1378), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1379), .B(n_1386), .Y(n_1378) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1388), .Y(n_1407) );
NAND2xp5_ASAP7_75t_L g1388 ( .A(n_1389), .B(n_1394), .Y(n_1388) );
INVx2_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
AOI22xp33_ASAP7_75t_L g1412 ( .A1(n_1391), .A2(n_1413), .B1(n_1414), .B2(n_1415), .Y(n_1412) );
AND2x4_ASAP7_75t_L g1391 ( .A(n_1392), .B(n_1393), .Y(n_1391) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1395), .Y(n_1406) );
AOI22xp5_ASAP7_75t_L g1516 ( .A1(n_1396), .A2(n_1399), .B1(n_1503), .B2(n_1517), .Y(n_1516) );
OAI21xp5_ASAP7_75t_L g1401 ( .A1(n_1402), .A2(n_1403), .B(n_1404), .Y(n_1401) );
OAI21xp33_ASAP7_75t_L g1405 ( .A1(n_1404), .A2(n_1406), .B(n_1407), .Y(n_1405) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1408), .Y(n_1489) );
XNOR2xp5_ASAP7_75t_L g1408 ( .A(n_1409), .B(n_1410), .Y(n_1408) );
NOR2x1_ASAP7_75t_L g1410 ( .A(n_1411), .B(n_1449), .Y(n_1410) );
NAND2xp5_ASAP7_75t_L g1411 ( .A(n_1412), .B(n_1416), .Y(n_1411) );
INVx3_ASAP7_75t_L g1532 ( .A(n_1414), .Y(n_1532) );
INVx2_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
HB1xp67_ASAP7_75t_L g1444 ( .A(n_1420), .Y(n_1444) );
OAI221xp5_ASAP7_75t_L g1421 ( .A1(n_1422), .A2(n_1425), .B1(n_1430), .B2(n_1434), .C(n_1438), .Y(n_1421) );
OAI211xp5_ASAP7_75t_L g1471 ( .A1(n_1426), .A2(n_1472), .B(n_1474), .C(n_1475), .Y(n_1471) );
OAI211xp5_ASAP7_75t_L g1811 ( .A1(n_1431), .A2(n_1812), .B(n_1813), .C(n_1814), .Y(n_1811) );
OAI21xp5_ASAP7_75t_SL g1434 ( .A1(n_1435), .A2(n_1436), .B(n_1437), .Y(n_1434) );
AOI22xp5_ASAP7_75t_L g1455 ( .A1(n_1442), .A2(n_1456), .B1(n_1458), .B2(n_1459), .Y(n_1455) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
INVx4_ASAP7_75t_L g1445 ( .A(n_1446), .Y(n_1445) );
INVx2_ASAP7_75t_L g1447 ( .A(n_1448), .Y(n_1447) );
NAND3xp33_ASAP7_75t_L g1449 ( .A(n_1450), .B(n_1478), .C(n_1484), .Y(n_1449) );
NOR3xp33_ASAP7_75t_SL g1450 ( .A(n_1451), .B(n_1465), .C(n_1468), .Y(n_1450) );
OAI21xp5_ASAP7_75t_SL g1451 ( .A1(n_1452), .A2(n_1454), .B(n_1455), .Y(n_1451) );
INVx1_ASAP7_75t_SL g1456 ( .A(n_1457), .Y(n_1456) );
INVx2_ASAP7_75t_SL g1459 ( .A(n_1460), .Y(n_1459) );
NAND2x2_ASAP7_75t_L g1460 ( .A(n_1461), .B(n_1463), .Y(n_1460) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1461), .Y(n_1477) );
INVx2_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
INVx2_ASAP7_75t_SL g1463 ( .A(n_1464), .Y(n_1463) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1467), .Y(n_1483) );
OAI21xp5_ASAP7_75t_L g1468 ( .A1(n_1469), .A2(n_1471), .B(n_1476), .Y(n_1468) );
INVx2_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
INVx2_ASAP7_75t_L g1877 ( .A(n_1470), .Y(n_1877) );
INVx2_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
NAND2xp5_ASAP7_75t_L g1478 ( .A(n_1479), .B(n_1480), .Y(n_1478) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
NAND2xp5_ASAP7_75t_L g1484 ( .A(n_1485), .B(n_1486), .Y(n_1484) );
AOI21xp5_ASAP7_75t_L g1493 ( .A1(n_1494), .A2(n_1514), .B(n_1515), .Y(n_1493) );
NAND4xp25_ASAP7_75t_L g1494 ( .A(n_1495), .B(n_1497), .C(n_1505), .D(n_1510), .Y(n_1494) );
OAI22xp5_ASAP7_75t_L g1809 ( .A1(n_1524), .A2(n_1810), .B1(n_1811), .B2(n_1815), .Y(n_1809) );
NAND2xp5_ASAP7_75t_L g1529 ( .A(n_1530), .B(n_1531), .Y(n_1529) );
INVx2_ASAP7_75t_L g1580 ( .A(n_1535), .Y(n_1580) );
XOR2x2_ASAP7_75t_L g1535 ( .A(n_1536), .B(n_1578), .Y(n_1535) );
NAND2xp5_ASAP7_75t_SL g1536 ( .A(n_1537), .B(n_1558), .Y(n_1536) );
NAND2xp5_ASAP7_75t_L g1539 ( .A(n_1540), .B(n_1547), .Y(n_1539) );
NOR2xp33_ASAP7_75t_L g1540 ( .A(n_1541), .B(n_1544), .Y(n_1540) );
NAND3xp33_ASAP7_75t_SL g1559 ( .A(n_1560), .B(n_1561), .C(n_1564), .Y(n_1559) );
INVx2_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
INVx4_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
INVx5_ASAP7_75t_L g1576 ( .A(n_1577), .Y(n_1576) );
OAI221xp5_ASAP7_75t_SL g1582 ( .A1(n_1583), .A2(n_1798), .B1(n_1800), .B2(n_1841), .C(n_1844), .Y(n_1582) );
NOR3xp33_ASAP7_75t_L g1583 ( .A(n_1584), .B(n_1778), .C(n_1792), .Y(n_1583) );
OAI221xp5_ASAP7_75t_L g1584 ( .A1(n_1585), .A2(n_1677), .B1(n_1699), .B2(n_1735), .C(n_1736), .Y(n_1584) );
OAI21xp5_ASAP7_75t_SL g1585 ( .A1(n_1586), .A2(n_1623), .B(n_1671), .Y(n_1585) );
OAI22xp5_ASAP7_75t_L g1794 ( .A1(n_1586), .A2(n_1650), .B1(n_1723), .B2(n_1795), .Y(n_1794) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
NAND2xp5_ASAP7_75t_SL g1587 ( .A(n_1588), .B(n_1618), .Y(n_1587) );
AOI211xp5_ASAP7_75t_L g1786 ( .A1(n_1588), .A2(n_1664), .B(n_1787), .C(n_1788), .Y(n_1786) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
OR2x2_ASAP7_75t_L g1589 ( .A(n_1590), .B(n_1605), .Y(n_1589) );
NAND2xp5_ASAP7_75t_L g1652 ( .A(n_1590), .B(n_1643), .Y(n_1652) );
AND2x2_ASAP7_75t_L g1682 ( .A(n_1590), .B(n_1666), .Y(n_1682) );
CKINVDCx5p33_ASAP7_75t_R g1690 ( .A(n_1590), .Y(n_1690) );
NAND2xp5_ASAP7_75t_L g1701 ( .A(n_1590), .B(n_1702), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1721 ( .A(n_1590), .B(n_1722), .Y(n_1721) );
OAI21xp5_ASAP7_75t_SL g1791 ( .A1(n_1590), .A2(n_1722), .B(n_1788), .Y(n_1791) );
INVx4_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
OR2x2_ASAP7_75t_L g1670 ( .A(n_1591), .B(n_1634), .Y(n_1670) );
AND2x2_ASAP7_75t_L g1678 ( .A(n_1591), .B(n_1679), .Y(n_1678) );
INVx4_ASAP7_75t_L g1687 ( .A(n_1591), .Y(n_1687) );
NOR2xp33_ASAP7_75t_L g1693 ( .A(n_1591), .B(n_1636), .Y(n_1693) );
NOR2xp33_ASAP7_75t_L g1697 ( .A(n_1591), .B(n_1698), .Y(n_1697) );
AOI322xp5_ASAP7_75t_L g1703 ( .A1(n_1591), .A2(n_1704), .A3(n_1706), .B1(n_1708), .B2(n_1710), .C1(n_1711), .C2(n_1713), .Y(n_1703) );
AND2x2_ASAP7_75t_L g1710 ( .A(n_1591), .B(n_1639), .Y(n_1710) );
NAND2xp5_ASAP7_75t_SL g1730 ( .A(n_1591), .B(n_1634), .Y(n_1730) );
NAND2xp5_ASAP7_75t_L g1777 ( .A(n_1591), .B(n_1618), .Y(n_1777) );
AND2x4_ASAP7_75t_SL g1591 ( .A(n_1592), .B(n_1600), .Y(n_1591) );
AND2x4_ASAP7_75t_L g1593 ( .A(n_1594), .B(n_1595), .Y(n_1593) );
AND2x6_ASAP7_75t_L g1598 ( .A(n_1594), .B(n_1599), .Y(n_1598) );
AND2x6_ASAP7_75t_L g1601 ( .A(n_1594), .B(n_1602), .Y(n_1601) );
AND2x2_ASAP7_75t_L g1603 ( .A(n_1594), .B(n_1604), .Y(n_1603) );
AND2x2_ASAP7_75t_L g1609 ( .A(n_1594), .B(n_1604), .Y(n_1609) );
NAND2xp5_ASAP7_75t_L g1657 ( .A(n_1594), .B(n_1595), .Y(n_1657) );
AND2x2_ASAP7_75t_L g1662 ( .A(n_1594), .B(n_1604), .Y(n_1662) );
AND2x2_ASAP7_75t_L g1595 ( .A(n_1596), .B(n_1597), .Y(n_1595) );
INVx2_ASAP7_75t_L g1659 ( .A(n_1598), .Y(n_1659) );
OAI21xp5_ASAP7_75t_L g1910 ( .A1(n_1604), .A2(n_1911), .B(n_1912), .Y(n_1910) );
INVx1_ASAP7_75t_L g1787 ( .A(n_1605), .Y(n_1787) );
OR2x2_ASAP7_75t_L g1605 ( .A(n_1606), .B(n_1610), .Y(n_1605) );
AND2x2_ASAP7_75t_L g1638 ( .A(n_1606), .B(n_1639), .Y(n_1638) );
OR2x2_ASAP7_75t_L g1647 ( .A(n_1606), .B(n_1648), .Y(n_1647) );
OR2x2_ASAP7_75t_L g1747 ( .A(n_1606), .B(n_1612), .Y(n_1747) );
NAND2xp5_ASAP7_75t_L g1781 ( .A(n_1606), .B(n_1693), .Y(n_1781) );
AND2x2_ASAP7_75t_L g1606 ( .A(n_1607), .B(n_1608), .Y(n_1606) );
AND2x2_ASAP7_75t_L g1634 ( .A(n_1607), .B(n_1608), .Y(n_1634) );
OR2x2_ASAP7_75t_L g1683 ( .A(n_1610), .B(n_1633), .Y(n_1683) );
INVx1_ASAP7_75t_L g1715 ( .A(n_1610), .Y(n_1715) );
OR2x2_ASAP7_75t_L g1729 ( .A(n_1610), .B(n_1730), .Y(n_1729) );
NAND2xp5_ASAP7_75t_L g1763 ( .A(n_1610), .B(n_1764), .Y(n_1763) );
NAND2xp5_ASAP7_75t_L g1610 ( .A(n_1611), .B(n_1615), .Y(n_1610) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1612), .Y(n_1611) );
OR2x2_ASAP7_75t_L g1636 ( .A(n_1612), .B(n_1615), .Y(n_1636) );
AND2x2_ASAP7_75t_L g1639 ( .A(n_1612), .B(n_1640), .Y(n_1639) );
AND2x2_ASAP7_75t_L g1643 ( .A(n_1612), .B(n_1615), .Y(n_1643) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1612), .Y(n_1707) );
NAND2xp5_ASAP7_75t_L g1734 ( .A(n_1612), .B(n_1634), .Y(n_1734) );
NAND3xp33_ASAP7_75t_L g1738 ( .A(n_1612), .B(n_1654), .C(n_1674), .Y(n_1738) );
AND2x2_ASAP7_75t_L g1612 ( .A(n_1613), .B(n_1614), .Y(n_1612) );
INVx2_ASAP7_75t_L g1640 ( .A(n_1615), .Y(n_1640) );
OR2x2_ASAP7_75t_L g1774 ( .A(n_1615), .B(n_1634), .Y(n_1774) );
NAND2x1p5_ASAP7_75t_L g1615 ( .A(n_1616), .B(n_1617), .Y(n_1615) );
AOI221xp5_ASAP7_75t_L g1677 ( .A1(n_1618), .A2(n_1650), .B1(n_1678), .B2(n_1680), .C(n_1691), .Y(n_1677) );
NAND2xp5_ASAP7_75t_L g1796 ( .A(n_1618), .B(n_1689), .Y(n_1796) );
INVx2_ASAP7_75t_L g1618 ( .A(n_1619), .Y(n_1618) );
AND2x2_ASAP7_75t_L g1625 ( .A(n_1619), .B(n_1626), .Y(n_1625) );
AND2x2_ASAP7_75t_L g1733 ( .A(n_1619), .B(n_1687), .Y(n_1733) );
OAI322xp33_ASAP7_75t_L g1748 ( .A1(n_1619), .A2(n_1631), .A3(n_1671), .B1(n_1749), .B2(n_1752), .C1(n_1753), .C2(n_1756), .Y(n_1748) );
OR2x2_ASAP7_75t_L g1760 ( .A(n_1619), .B(n_1673), .Y(n_1760) );
INVx1_ASAP7_75t_L g1619 ( .A(n_1620), .Y(n_1619) );
OR2x2_ASAP7_75t_L g1645 ( .A(n_1620), .B(n_1626), .Y(n_1645) );
INVx1_ASAP7_75t_L g1667 ( .A(n_1620), .Y(n_1667) );
NAND2xp5_ASAP7_75t_L g1620 ( .A(n_1621), .B(n_1622), .Y(n_1620) );
OAI211xp5_ASAP7_75t_L g1623 ( .A1(n_1624), .A2(n_1630), .B(n_1641), .C(n_1663), .Y(n_1623) );
NOR2xp33_ASAP7_75t_L g1728 ( .A(n_1624), .B(n_1729), .Y(n_1728) );
OAI21xp5_ASAP7_75t_L g1797 ( .A1(n_1624), .A2(n_1645), .B(n_1711), .Y(n_1797) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
AOI21xp5_ASAP7_75t_L g1696 ( .A1(n_1625), .A2(n_1653), .B(n_1697), .Y(n_1696) );
NAND2xp5_ASAP7_75t_L g1727 ( .A(n_1625), .B(n_1668), .Y(n_1727) );
AND2x2_ASAP7_75t_L g1740 ( .A(n_1625), .B(n_1741), .Y(n_1740) );
INVx2_ASAP7_75t_L g1650 ( .A(n_1626), .Y(n_1650) );
OAI21xp33_ASAP7_75t_L g1651 ( .A1(n_1626), .A2(n_1652), .B(n_1653), .Y(n_1651) );
AND2x2_ASAP7_75t_L g1713 ( .A(n_1626), .B(n_1674), .Y(n_1713) );
OR2x2_ASAP7_75t_L g1723 ( .A(n_1626), .B(n_1667), .Y(n_1723) );
OR2x2_ASAP7_75t_L g1752 ( .A(n_1626), .B(n_1674), .Y(n_1752) );
INVx1_ASAP7_75t_L g1755 ( .A(n_1626), .Y(n_1755) );
AND2x2_ASAP7_75t_L g1790 ( .A(n_1626), .B(n_1673), .Y(n_1790) );
INVx2_ASAP7_75t_L g1626 ( .A(n_1627), .Y(n_1626) );
OR2x2_ASAP7_75t_L g1695 ( .A(n_1627), .B(n_1667), .Y(n_1695) );
NAND2xp5_ASAP7_75t_L g1627 ( .A(n_1628), .B(n_1629), .Y(n_1627) );
AND2x2_ASAP7_75t_L g1630 ( .A(n_1631), .B(n_1637), .Y(n_1630) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
AND2x2_ASAP7_75t_L g1689 ( .A(n_1632), .B(n_1690), .Y(n_1689) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1633), .B(n_1635), .Y(n_1632) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_1633), .B(n_1639), .Y(n_1679) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1633), .B(n_1686), .Y(n_1685) );
INVx1_ASAP7_75t_L g1633 ( .A(n_1634), .Y(n_1633) );
AND2x2_ASAP7_75t_L g1642 ( .A(n_1634), .B(n_1643), .Y(n_1642) );
OR2x2_ASAP7_75t_L g1698 ( .A(n_1634), .B(n_1640), .Y(n_1698) );
AND2x2_ASAP7_75t_L g1706 ( .A(n_1634), .B(n_1707), .Y(n_1706) );
AND2x2_ASAP7_75t_L g1769 ( .A(n_1634), .B(n_1640), .Y(n_1769) );
NAND2xp5_ASAP7_75t_L g1720 ( .A(n_1635), .B(n_1721), .Y(n_1720) );
AND2x2_ASAP7_75t_L g1750 ( .A(n_1635), .B(n_1751), .Y(n_1750) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1636), .Y(n_1635) );
OR2x2_ASAP7_75t_L g1669 ( .A(n_1636), .B(n_1670), .Y(n_1669) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
NAND2xp5_ASAP7_75t_L g1756 ( .A(n_1639), .B(n_1757), .Y(n_1756) );
INVx1_ASAP7_75t_L g1764 ( .A(n_1639), .Y(n_1764) );
OAI211xp5_ASAP7_75t_L g1772 ( .A1(n_1639), .A2(n_1773), .B(n_1775), .C(n_1776), .Y(n_1772) );
NAND3xp33_ASAP7_75t_L g1785 ( .A(n_1639), .B(n_1672), .C(n_1682), .Y(n_1785) );
AOI221xp5_ASAP7_75t_L g1641 ( .A1(n_1642), .A2(n_1644), .B1(n_1646), .B2(n_1649), .C(n_1651), .Y(n_1641) );
NAND2x1_ASAP7_75t_L g1712 ( .A(n_1642), .B(n_1687), .Y(n_1712) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1643), .Y(n_1648) );
INVx1_ASAP7_75t_L g1644 ( .A(n_1645), .Y(n_1644) );
OR2x2_ASAP7_75t_L g1717 ( .A(n_1645), .B(n_1718), .Y(n_1717) );
OAI21xp33_ASAP7_75t_L g1745 ( .A1(n_1646), .A2(n_1716), .B(n_1746), .Y(n_1745) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
NOR2x1_ASAP7_75t_L g1686 ( .A(n_1648), .B(n_1687), .Y(n_1686) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1650), .Y(n_1649) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1653), .Y(n_1735) );
OAI321xp33_ASAP7_75t_L g1766 ( .A1(n_1653), .A2(n_1752), .A3(n_1767), .B1(n_1768), .B2(n_1771), .C(n_1772), .Y(n_1766) );
OAI221xp5_ASAP7_75t_L g1778 ( .A1(n_1653), .A2(n_1779), .B1(n_1786), .B2(n_1789), .C(n_1791), .Y(n_1778) );
INVx2_ASAP7_75t_L g1653 ( .A(n_1654), .Y(n_1653) );
INVx1_ASAP7_75t_L g1654 ( .A(n_1655), .Y(n_1654) );
NAND2xp5_ASAP7_75t_L g1671 ( .A(n_1655), .B(n_1672), .Y(n_1671) );
NOR2xp33_ASAP7_75t_SL g1775 ( .A(n_1655), .B(n_1674), .Y(n_1775) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
OAI221xp5_ASAP7_75t_L g1656 ( .A1(n_1657), .A2(n_1658), .B1(n_1659), .B2(n_1660), .C(n_1661), .Y(n_1656) );
HB1xp67_ASAP7_75t_L g1799 ( .A(n_1662), .Y(n_1799) );
INVxp67_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
AND2x2_ASAP7_75t_L g1664 ( .A(n_1665), .B(n_1668), .Y(n_1664) );
NAND2xp5_ASAP7_75t_L g1684 ( .A(n_1665), .B(n_1685), .Y(n_1684) );
NAND2xp5_ASAP7_75t_L g1749 ( .A(n_1665), .B(n_1750), .Y(n_1749) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1666), .Y(n_1665) );
OR2x2_ASAP7_75t_L g1705 ( .A(n_1666), .B(n_1673), .Y(n_1705) );
NOR3xp33_ASAP7_75t_L g1743 ( .A(n_1666), .B(n_1729), .C(n_1744), .Y(n_1743) );
INVx1_ASAP7_75t_L g1666 ( .A(n_1667), .Y(n_1666) );
INVx1_ASAP7_75t_L g1668 ( .A(n_1669), .Y(n_1668) );
AOI221xp5_ASAP7_75t_L g1758 ( .A1(n_1669), .A2(n_1704), .B1(n_1756), .B2(n_1759), .C(n_1761), .Y(n_1758) );
INVx1_ASAP7_75t_L g1757 ( .A(n_1670), .Y(n_1757) );
AOI31xp33_ASAP7_75t_L g1761 ( .A1(n_1672), .A2(n_1751), .A3(n_1762), .B(n_1765), .Y(n_1761) );
NOR2xp33_ASAP7_75t_L g1788 ( .A(n_1672), .B(n_1683), .Y(n_1788) );
CKINVDCx14_ASAP7_75t_R g1672 ( .A(n_1673), .Y(n_1672) );
OR2x2_ASAP7_75t_L g1709 ( .A(n_1673), .B(n_1695), .Y(n_1709) );
OR2x2_ASAP7_75t_L g1726 ( .A(n_1673), .B(n_1723), .Y(n_1726) );
OAI21xp5_ASAP7_75t_L g1768 ( .A1(n_1673), .A2(n_1769), .B(n_1770), .Y(n_1768) );
INVx3_ASAP7_75t_L g1673 ( .A(n_1674), .Y(n_1673) );
INVx1_ASAP7_75t_L g1718 ( .A(n_1674), .Y(n_1718) );
AND2x2_ASAP7_75t_L g1754 ( .A(n_1674), .B(n_1755), .Y(n_1754) );
AND2x2_ASAP7_75t_L g1674 ( .A(n_1675), .B(n_1676), .Y(n_1674) );
INVx1_ASAP7_75t_L g1694 ( .A(n_1679), .Y(n_1694) );
OAI211xp5_ASAP7_75t_L g1680 ( .A1(n_1681), .A2(n_1683), .B(n_1684), .C(n_1688), .Y(n_1680) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
INVx1_ASAP7_75t_L g1702 ( .A(n_1683), .Y(n_1702) );
O2A1O1Ixp33_ASAP7_75t_SL g1792 ( .A1(n_1683), .A2(n_1793), .B(n_1794), .C(n_1797), .Y(n_1792) );
INVx1_ASAP7_75t_L g1725 ( .A(n_1686), .Y(n_1725) );
O2A1O1Ixp33_ASAP7_75t_L g1779 ( .A1(n_1686), .A2(n_1704), .B(n_1780), .C(n_1782), .Y(n_1779) );
CKINVDCx5p33_ASAP7_75t_R g1741 ( .A(n_1687), .Y(n_1741) );
NOR2xp33_ASAP7_75t_L g1746 ( .A(n_1687), .B(n_1747), .Y(n_1746) );
INVx1_ASAP7_75t_L g1688 ( .A(n_1689), .Y(n_1688) );
OR2x2_ASAP7_75t_L g1783 ( .A(n_1690), .B(n_1734), .Y(n_1783) );
A2O1A1Ixp33_ASAP7_75t_L g1691 ( .A1(n_1692), .A2(n_1694), .B(n_1695), .C(n_1696), .Y(n_1691) );
INVx1_ASAP7_75t_L g1692 ( .A(n_1693), .Y(n_1692) );
OAI211xp5_ASAP7_75t_SL g1700 ( .A1(n_1695), .A2(n_1701), .B(n_1703), .C(n_1714), .Y(n_1700) );
CKINVDCx5p33_ASAP7_75t_R g1765 ( .A(n_1695), .Y(n_1765) );
NAND2xp5_ASAP7_75t_L g1784 ( .A(n_1697), .B(n_1713), .Y(n_1784) );
INVx1_ASAP7_75t_L g1770 ( .A(n_1698), .Y(n_1770) );
NOR5xp2_ASAP7_75t_L g1699 ( .A(n_1700), .B(n_1719), .C(n_1724), .D(n_1728), .E(n_1731), .Y(n_1699) );
INVx1_ASAP7_75t_L g1704 ( .A(n_1705), .Y(n_1704) );
INVx1_ASAP7_75t_L g1708 ( .A(n_1709), .Y(n_1708) );
INVx1_ASAP7_75t_L g1767 ( .A(n_1710), .Y(n_1767) );
INVx1_ASAP7_75t_L g1711 ( .A(n_1712), .Y(n_1711) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1713), .Y(n_1744) );
NAND2xp5_ASAP7_75t_L g1714 ( .A(n_1715), .B(n_1716), .Y(n_1714) );
INVx1_ASAP7_75t_L g1716 ( .A(n_1717), .Y(n_1716) );
INVx1_ASAP7_75t_L g1719 ( .A(n_1720), .Y(n_1719) );
INVx1_ASAP7_75t_L g1771 ( .A(n_1721), .Y(n_1771) );
CKINVDCx5p33_ASAP7_75t_R g1722 ( .A(n_1723), .Y(n_1722) );
OAI21xp33_ASAP7_75t_L g1724 ( .A1(n_1725), .A2(n_1726), .B(n_1727), .Y(n_1724) );
INVx1_ASAP7_75t_L g1751 ( .A(n_1730), .Y(n_1751) );
NOR2xp33_ASAP7_75t_L g1731 ( .A(n_1732), .B(n_1734), .Y(n_1731) );
INVx1_ASAP7_75t_L g1732 ( .A(n_1733), .Y(n_1732) );
NOR4xp25_ASAP7_75t_L g1736 ( .A(n_1737), .B(n_1748), .C(n_1758), .D(n_1766), .Y(n_1736) );
OAI211xp5_ASAP7_75t_SL g1737 ( .A1(n_1738), .A2(n_1739), .B(n_1742), .C(n_1745), .Y(n_1737) );
INVxp67_ASAP7_75t_L g1739 ( .A(n_1740), .Y(n_1739) );
INVxp67_ASAP7_75t_SL g1742 ( .A(n_1743), .Y(n_1742) );
OAI211xp5_ASAP7_75t_L g1782 ( .A1(n_1753), .A2(n_1783), .B(n_1784), .C(n_1785), .Y(n_1782) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1754), .Y(n_1753) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1760), .Y(n_1759) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1763), .Y(n_1762) );
INVx1_ASAP7_75t_L g1773 ( .A(n_1774), .Y(n_1773) );
INVx1_ASAP7_75t_L g1793 ( .A(n_1775), .Y(n_1793) );
INVx1_ASAP7_75t_L g1776 ( .A(n_1777), .Y(n_1776) );
INVx1_ASAP7_75t_L g1780 ( .A(n_1781), .Y(n_1780) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1790), .Y(n_1789) );
INVxp67_ASAP7_75t_L g1795 ( .A(n_1796), .Y(n_1795) );
INVx4_ASAP7_75t_L g1798 ( .A(n_1799), .Y(n_1798) );
HB1xp67_ASAP7_75t_L g1801 ( .A(n_1802), .Y(n_1801) );
NAND4xp75_ASAP7_75t_L g1802 ( .A(n_1803), .B(n_1808), .C(n_1822), .D(n_1839), .Y(n_1802) );
NAND2xp5_ASAP7_75t_L g1823 ( .A(n_1824), .B(n_1828), .Y(n_1823) );
OAI221xp5_ASAP7_75t_L g1832 ( .A1(n_1833), .A2(n_1834), .B1(n_1835), .B2(n_1837), .C(n_1838), .Y(n_1832) );
BUFx3_ASAP7_75t_L g1835 ( .A(n_1836), .Y(n_1835) );
INVxp67_ASAP7_75t_L g1841 ( .A(n_1842), .Y(n_1841) );
BUFx3_ASAP7_75t_L g1842 ( .A(n_1843), .Y(n_1842) );
HB1xp67_ASAP7_75t_L g1847 ( .A(n_1848), .Y(n_1847) );
NAND3xp33_ASAP7_75t_L g1849 ( .A(n_1850), .B(n_1880), .C(n_1893), .Y(n_1849) );
NOR2xp33_ASAP7_75t_L g1850 ( .A(n_1851), .B(n_1870), .Y(n_1850) );
OAI22xp33_ASAP7_75t_L g1852 ( .A1(n_1853), .A2(n_1854), .B1(n_1856), .B2(n_1857), .Y(n_1852) );
BUFx4f_ASAP7_75t_SL g1854 ( .A(n_1855), .Y(n_1854) );
OAI22xp33_ASAP7_75t_L g1866 ( .A1(n_1855), .A2(n_1867), .B1(n_1868), .B2(n_1869), .Y(n_1866) );
INVx1_ASAP7_75t_L g1857 ( .A(n_1858), .Y(n_1857) );
OAI33xp33_ASAP7_75t_L g1870 ( .A1(n_1871), .A2(n_1873), .A3(n_1874), .B1(n_1876), .B2(n_1877), .B3(n_1878), .Y(n_1870) );
INVx1_ASAP7_75t_L g1871 ( .A(n_1872), .Y(n_1871) );
AOI22xp33_ASAP7_75t_L g1883 ( .A1(n_1884), .A2(n_1885), .B1(n_1886), .B2(n_1888), .Y(n_1883) );
INVx2_ASAP7_75t_L g1886 ( .A(n_1887), .Y(n_1886) );
OAI31xp33_ASAP7_75t_L g1893 ( .A1(n_1894), .A2(n_1896), .A3(n_1903), .B(n_1907), .Y(n_1893) );
HB1xp67_ASAP7_75t_L g1897 ( .A(n_1898), .Y(n_1897) );
INVx2_ASAP7_75t_L g1905 ( .A(n_1906), .Y(n_1905) );
INVx1_ASAP7_75t_L g1908 ( .A(n_1909), .Y(n_1908) );
INVx1_ASAP7_75t_L g1909 ( .A(n_1910), .Y(n_1909) );
INVx1_ASAP7_75t_L g1912 ( .A(n_1913), .Y(n_1912) );
endmodule