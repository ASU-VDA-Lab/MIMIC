module real_jpeg_31142_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_0),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_0),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_1),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_1),
.B(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_1),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_1),
.B(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_2),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_2),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_2),
.B(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

NAND2x1_ASAP7_75t_SL g66 ( 
.A(n_3),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g145 ( 
.A(n_3),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_3),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_4),
.Y(n_76)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_5),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_6),
.B(n_127),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_7),
.Y(n_123)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_7),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_8),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_8),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_8),
.B(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_9),
.Y(n_98)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_11),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_11),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_11),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_11),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_11),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_11),
.B(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_12),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_12),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_13),
.B(n_103),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_135),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_133),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_83),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_17),
.B(n_83),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_44),
.C(n_63),
.Y(n_17)
);

INVxp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_19),
.B(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_28),
.B2(n_29),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_21),
.B(n_29),
.C(n_36),
.Y(n_105)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_27),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_27),
.Y(n_164)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

XOR2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_32),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_32),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_34),
.Y(n_178)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_41),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_37),
.A2(n_41),
.B1(n_42),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_37),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_42),
.B(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_44),
.A2(n_45),
.B1(n_64),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.C(n_57),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_46),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_140)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_57),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_58),
.B(n_111),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_61),
.Y(n_183)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_64),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_77),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_72),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_66),
.B(n_72),
.C(n_77),
.Y(n_132)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_106),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_105),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_100),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_93),
.B1(n_94),
.B2(n_99),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_88),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_102),
.A2(n_126),
.B1(n_130),
.B2(n_131),
.Y(n_125)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_124),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_119),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_114),
.B2(n_118),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_132),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21x1_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_155),
.B(n_199),
.Y(n_135)
);

NOR2xp67_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_152),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_137),
.B(n_152),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.C(n_144),
.Y(n_137)
);

XNOR2x2_ASAP7_75t_L g195 ( 
.A(n_138),
.B(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_141),
.A2(n_142),
.B1(n_144),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_144),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_149),
.Y(n_159)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI21x1_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_193),
.B(n_198),
.Y(n_155)
);

OAI21x1_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_179),
.B(n_192),
.Y(n_156)
);

NOR2x1_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_172),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_158),
.B(n_172),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_162),
.C(n_165),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_165),
.B2(n_166),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_177),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_173),
.B(n_186),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_185),
.B(n_191),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_184),
.Y(n_191)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp67_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_195),
.Y(n_198)
);


endmodule