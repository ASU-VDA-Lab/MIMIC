module fake_jpeg_3640_n_534 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_534);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx4f_ASAP7_75t_SL g165 ( 
.A(n_62),
.Y(n_165)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_66),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_25),
.B(n_15),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_67),
.B(n_92),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_71),
.Y(n_167)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_74),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_17),
.B(n_8),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_77),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_23),
.B(n_8),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_79),
.Y(n_161)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx6_ASAP7_75t_SL g168 ( 
.A(n_83),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_84),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_85),
.Y(n_172)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_90),
.B(n_93),
.Y(n_143)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_36),
.B(n_15),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_35),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_54),
.B(n_8),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_94),
.B(n_95),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_38),
.B(n_6),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_14),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_96),
.B(n_102),
.Y(n_166)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_20),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

BUFx2_ASAP7_75t_SL g111 ( 
.A(n_104),
.Y(n_111)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_105),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_37),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_106),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_37),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_110),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

CKINVDCx12_ASAP7_75t_R g199 ( 
.A(n_113),
.Y(n_199)
);

AO22x2_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_33),
.B1(n_52),
.B2(n_24),
.Y(n_120)
);

NOR2x1_ASAP7_75t_L g208 ( 
.A(n_120),
.B(n_104),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_55),
.A2(n_33),
.B1(n_39),
.B2(n_44),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_125),
.A2(n_18),
.B1(n_80),
.B2(n_72),
.Y(n_180)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_57),
.A2(n_53),
.B1(n_45),
.B2(n_24),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_135),
.A2(n_142),
.B1(n_149),
.B2(n_42),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_59),
.A2(n_22),
.B1(n_47),
.B2(n_26),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_138),
.A2(n_41),
.B1(n_40),
.B2(n_26),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_86),
.A2(n_103),
.B1(n_91),
.B2(n_79),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_56),
.A2(n_53),
.B1(n_45),
.B2(n_52),
.Y(n_149)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_70),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_156),
.Y(n_186)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_97),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_98),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_81),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_62),
.A2(n_30),
.B(n_46),
.Y(n_169)
);

OR2x2_ASAP7_75t_SL g181 ( 
.A(n_169),
.B(n_48),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_107),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_173),
.Y(n_229)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_69),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_174),
.Y(n_223)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_65),
.Y(n_175)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_30),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_176),
.B(n_190),
.Y(n_232)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_177),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_166),
.A2(n_71),
.B1(n_85),
.B2(n_46),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_178),
.B(n_208),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_131),
.B(n_114),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_179),
.B(n_204),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_180),
.A2(n_205),
.B1(n_211),
.B2(n_124),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_181),
.Y(n_257)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_182),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_120),
.B(n_108),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_183),
.B(n_222),
.Y(n_262)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_185),
.Y(n_249)
);

INVxp33_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_187),
.Y(n_252)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_145),
.B(n_114),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_191),
.A2(n_203),
.B1(n_219),
.B2(n_220),
.Y(n_241)
);

OA22x2_ASAP7_75t_L g259 ( 
.A1(n_192),
.A2(n_153),
.B1(n_159),
.B2(n_129),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_145),
.B(n_101),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_193),
.B(n_207),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_194),
.Y(n_265)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_196),
.Y(n_230)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_126),
.Y(n_197)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_197),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_201),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_137),
.B(n_41),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_202),
.B(n_218),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_112),
.A2(n_40),
.B1(n_47),
.B2(n_43),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_147),
.B(n_22),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_L g205 ( 
.A1(n_149),
.A2(n_75),
.B1(n_63),
.B2(n_82),
.Y(n_205)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_206),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_116),
.B(n_43),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_143),
.A2(n_58),
.B1(n_60),
.B2(n_68),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_124),
.B1(n_160),
.B2(n_130),
.Y(n_238)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_148),
.Y(n_210)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_210),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_120),
.A2(n_88),
.B1(n_84),
.B2(n_66),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_118),
.Y(n_212)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_212),
.Y(n_267)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_213),
.Y(n_269)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_143),
.Y(n_214)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

CKINVDCx12_ASAP7_75t_R g215 ( 
.A(n_165),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_215),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_117),
.Y(n_216)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_161),
.Y(n_217)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_165),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_112),
.A2(n_42),
.B1(n_18),
.B2(n_19),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_163),
.A2(n_49),
.B1(n_9),
.B2(n_10),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_127),
.Y(n_221)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_221),
.Y(n_270)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_122),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_127),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_225),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_132),
.B(n_9),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_172),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_226),
.B(n_227),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_136),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_139),
.B(n_9),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_228),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_183),
.A2(n_135),
.B(n_121),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_234),
.A2(n_258),
.B(n_229),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_235),
.A2(n_250),
.B1(n_254),
.B2(n_214),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_238),
.A2(n_245),
.B1(n_268),
.B2(n_217),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_178),
.A2(n_171),
.B1(n_157),
.B2(n_158),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_183),
.A2(n_208),
.B1(n_193),
.B2(n_187),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_176),
.A2(n_180),
.B1(n_211),
.B2(n_181),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_205),
.A2(n_115),
.B(n_154),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_259),
.B(n_177),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_191),
.A2(n_134),
.B1(n_130),
.B2(n_160),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_271),
.B(n_273),
.Y(n_319)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_272),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_262),
.Y(n_273)
);

AND2x6_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_190),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_274),
.B(n_292),
.Y(n_306)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_275),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_260),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_276),
.B(n_280),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_277),
.A2(n_197),
.B1(n_185),
.B2(n_182),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_242),
.B(n_228),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_278),
.B(n_287),
.Y(n_304)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_279),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_262),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_281),
.Y(n_318)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_282),
.Y(n_329)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_233),
.Y(n_283)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_283),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_222),
.C(n_195),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_240),
.C(n_231),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_247),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_285),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_286),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_242),
.B(n_186),
.Y(n_287)
);

AOI32xp33_ASAP7_75t_L g288 ( 
.A1(n_230),
.A2(n_227),
.A3(n_224),
.B1(n_221),
.B2(n_213),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_288),
.A2(n_291),
.B(n_290),
.Y(n_321)
);

NAND2xp33_ASAP7_75t_SL g328 ( 
.A(n_289),
.B(n_259),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_252),
.A2(n_188),
.B(n_217),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_290),
.A2(n_231),
.B(n_258),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_255),
.A2(n_200),
.B(n_184),
.Y(n_291)
);

A2O1A1Ixp33_ASAP7_75t_L g292 ( 
.A1(n_250),
.A2(n_133),
.B(n_119),
.C(n_144),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_230),
.B(n_232),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_300),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_244),
.B(n_201),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_294),
.B(n_295),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_232),
.B(n_244),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_237),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_298),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_297),
.Y(n_311)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_237),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_251),
.B(n_266),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_299),
.B(n_303),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_263),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_270),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_301),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_246),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_302),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_240),
.B(n_184),
.Y(n_303)
);

OAI32xp33_ASAP7_75t_L g305 ( 
.A1(n_293),
.A2(n_262),
.A3(n_255),
.B1(n_254),
.B2(n_252),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_305),
.B(n_287),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_313),
.C(n_315),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_273),
.B(n_255),
.C(n_234),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_295),
.B(n_241),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_321),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_323),
.A2(n_328),
.B(n_291),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_289),
.A2(n_235),
.B(n_259),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_325),
.A2(n_303),
.B(n_279),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_277),
.A2(n_251),
.B1(n_259),
.B2(n_164),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_326),
.A2(n_330),
.B1(n_292),
.B2(n_275),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_301),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_276),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_328),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_334),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_319),
.Y(n_335)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_335),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_324),
.B(n_278),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_336),
.B(n_337),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_324),
.B(n_299),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_307),
.Y(n_338)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_338),
.Y(n_371)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_339),
.Y(n_383)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_314),
.Y(n_340)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_340),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_342),
.A2(n_327),
.B1(n_322),
.B2(n_329),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_312),
.B(n_294),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_343),
.B(n_309),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_344),
.A2(n_353),
.B(n_334),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_304),
.B(n_302),
.Y(n_345)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_345),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_304),
.B(n_300),
.Y(n_346)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_346),
.Y(n_392)
);

AO21x1_ASAP7_75t_L g347 ( 
.A1(n_306),
.A2(n_297),
.B(n_274),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_347),
.B(n_352),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_325),
.A2(n_297),
.B1(n_292),
.B2(n_280),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_348),
.A2(n_331),
.B1(n_330),
.B2(n_305),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_308),
.B(n_284),
.C(n_274),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_349),
.B(n_341),
.C(n_313),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_319),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_350),
.B(n_314),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_351),
.A2(n_360),
.B(n_361),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g352 ( 
.A(n_317),
.B(n_288),
.Y(n_352)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_352),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_323),
.B(n_298),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_307),
.Y(n_354)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_354),
.Y(n_384)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_307),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g388 ( 
.A1(n_355),
.A2(n_356),
.B1(n_358),
.B2(n_362),
.Y(n_388)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_307),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_320),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_359),
.A2(n_310),
.B1(n_316),
.B2(n_333),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_321),
.A2(n_311),
.B(n_325),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_311),
.A2(n_296),
.B(n_283),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_312),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_363),
.B(n_387),
.C(n_338),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_364),
.A2(n_334),
.B(n_353),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_351),
.A2(n_326),
.B1(n_317),
.B2(n_306),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_365),
.A2(n_366),
.B1(n_372),
.B2(n_379),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_308),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_370),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_313),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_351),
.A2(n_309),
.B1(n_318),
.B2(n_331),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_373),
.B(n_374),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_341),
.B(n_315),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_375),
.B(n_347),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_376),
.A2(n_385),
.B1(n_389),
.B2(n_285),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_356),
.A2(n_330),
.B1(n_305),
.B2(n_316),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_380),
.Y(n_421)
);

BUFx12_ASAP7_75t_L g381 ( 
.A(n_360),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_381),
.B(n_382),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_337),
.B(n_233),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_336),
.B(n_315),
.Y(n_386)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_386),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_341),
.B(n_327),
.C(n_322),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_352),
.A2(n_310),
.B1(n_320),
.B2(n_329),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_388),
.A2(n_362),
.B1(n_357),
.B2(n_344),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_394),
.A2(n_400),
.B1(n_405),
.B2(n_415),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_397),
.B(n_399),
.Y(n_437)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_390),
.Y(n_398)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_398),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_368),
.B(n_347),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_365),
.A2(n_357),
.B1(n_348),
.B2(n_342),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_387),
.B(n_347),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_402),
.B(n_407),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_364),
.A2(n_346),
.B(n_345),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_403),
.A2(n_409),
.B(n_413),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_379),
.A2(n_348),
.B1(n_342),
.B2(n_353),
.Y(n_405)
);

AOI21xp33_ASAP7_75t_L g406 ( 
.A1(n_369),
.A2(n_343),
.B(n_361),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_406),
.B(n_414),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_375),
.B(n_334),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_410),
.B(n_412),
.C(n_416),
.Y(n_429)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_392),
.Y(n_411)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_411),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_363),
.B(n_358),
.C(n_355),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_391),
.A2(n_353),
.B(n_339),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_370),
.B(n_354),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_372),
.A2(n_340),
.B1(n_359),
.B2(n_332),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_384),
.B(n_332),
.C(n_236),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_378),
.A2(n_340),
.B1(n_359),
.B2(n_282),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_417),
.A2(n_422),
.B1(n_377),
.B2(n_367),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_383),
.B(n_359),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_391),
.C(n_389),
.Y(n_434)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_384),
.Y(n_419)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_419),
.Y(n_446)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_371),
.Y(n_420)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_420),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_423),
.A2(n_399),
.B1(n_414),
.B2(n_397),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_418),
.B(n_377),
.Y(n_424)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_424),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_401),
.A2(n_376),
.B1(n_393),
.B2(n_378),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_427),
.A2(n_445),
.B1(n_409),
.B2(n_415),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_396),
.Y(n_430)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_430),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_367),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_431),
.B(n_434),
.Y(n_458)
);

BUFx5_ASAP7_75t_L g433 ( 
.A(n_404),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_433),
.Y(n_462)
);

CKINVDCx14_ASAP7_75t_R g436 ( 
.A(n_408),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_436),
.B(n_442),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_410),
.B(n_393),
.C(n_380),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_438),
.B(n_444),
.C(n_395),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_413),
.A2(n_381),
.B(n_285),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_439),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_421),
.B(n_272),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_441),
.Y(n_455)
);

CKINVDCx14_ASAP7_75t_R g442 ( 
.A(n_416),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_395),
.B(n_381),
.C(n_236),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_422),
.A2(n_247),
.B1(n_265),
.B2(n_216),
.Y(n_445)
);

NOR2x1_ASAP7_75t_L g448 ( 
.A(n_438),
.B(n_402),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_448),
.B(n_437),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_449),
.A2(n_452),
.B1(n_427),
.B2(n_426),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_429),
.B(n_412),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_450),
.B(n_456),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_440),
.B(n_407),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_L g477 ( 
.A(n_451),
.B(n_440),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_443),
.A2(n_405),
.B1(n_394),
.B2(n_400),
.Y(n_452)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_454),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_443),
.A2(n_265),
.B1(n_194),
.B2(n_243),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_457),
.A2(n_445),
.B1(n_428),
.B2(n_463),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_L g459 ( 
.A(n_429),
.B(n_269),
.Y(n_459)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_459),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_267),
.C(n_256),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_461),
.B(n_465),
.Y(n_471)
);

AOI221xp5_ASAP7_75t_L g464 ( 
.A1(n_432),
.A2(n_267),
.B1(n_272),
.B2(n_256),
.C(n_261),
.Y(n_464)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_464),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_430),
.B(n_261),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_SL g466 ( 
.A1(n_447),
.A2(n_430),
.B1(n_431),
.B2(n_441),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_466),
.A2(n_467),
.B1(n_189),
.B2(n_198),
.Y(n_497)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_468),
.Y(n_488)
);

FAx1_ASAP7_75t_SL g473 ( 
.A(n_452),
.B(n_434),
.CI(n_426),
.CON(n_473),
.SN(n_473)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_473),
.B(n_474),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_462),
.B(n_458),
.Y(n_474)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_453),
.Y(n_476)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_476),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_433),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_478),
.A2(n_451),
.B1(n_461),
.B2(n_425),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_425),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_480),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_456),
.B(n_424),
.C(n_437),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_447),
.A2(n_439),
.B(n_428),
.Y(n_481)
);

XOR2x2_ASAP7_75t_L g491 ( 
.A(n_481),
.B(n_446),
.Y(n_491)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_455),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_482),
.B(n_446),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_470),
.B(n_435),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_483),
.A2(n_486),
.B1(n_490),
.B2(n_493),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_448),
.C(n_449),
.Y(n_485)
);

NOR2xp67_ASAP7_75t_SL g502 ( 
.A(n_485),
.B(n_494),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_472),
.B(n_435),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_469),
.A2(n_455),
.B1(n_460),
.B2(n_454),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_487),
.A2(n_226),
.B1(n_206),
.B2(n_223),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_467),
.A2(n_457),
.B(n_428),
.Y(n_489)
);

OAI21xp33_ASAP7_75t_L g506 ( 
.A1(n_489),
.A2(n_188),
.B(n_212),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_491),
.B(n_496),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_471),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_495),
.A2(n_497),
.B1(n_475),
.B2(n_468),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_480),
.B(n_249),
.C(n_239),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_498),
.B(n_492),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_499),
.A2(n_500),
.B(n_504),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_485),
.B(n_478),
.C(n_481),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_503),
.A2(n_506),
.B1(n_146),
.B2(n_170),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_484),
.B(n_466),
.C(n_473),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_473),
.C(n_199),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_505),
.B(n_508),
.C(n_500),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_496),
.B(n_249),
.C(n_239),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_488),
.B(n_264),
.C(n_134),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_509),
.B(n_510),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_489),
.B(n_264),
.C(n_210),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_511),
.B(n_170),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_512),
.B(n_516),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_502),
.B(n_491),
.C(n_487),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_514),
.B(n_519),
.Y(n_525)
);

NAND3xp33_ASAP7_75t_L g515 ( 
.A(n_507),
.B(n_497),
.C(n_223),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_515),
.A2(n_510),
.B(n_509),
.Y(n_521)
);

AOI322xp5_ASAP7_75t_L g516 ( 
.A1(n_506),
.A2(n_146),
.A3(n_170),
.B1(n_164),
.B2(n_136),
.C1(n_113),
.C2(n_111),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_517),
.B(n_518),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_501),
.B(n_9),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_521),
.B(n_524),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_520),
.B(n_111),
.C(n_49),
.Y(n_524)
);

AOI322xp5_ASAP7_75t_L g526 ( 
.A1(n_522),
.A2(n_513),
.A3(n_516),
.B1(n_10),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_526),
.A2(n_527),
.B(n_11),
.Y(n_530)
);

AOI322xp5_ASAP7_75t_L g527 ( 
.A1(n_525),
.A2(n_6),
.A3(n_13),
.B1(n_11),
.B2(n_5),
.C1(n_14),
.C2(n_2),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_528),
.A2(n_523),
.B(n_11),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_529),
.A2(n_530),
.B(n_13),
.Y(n_531)
);

O2A1O1Ixp33_ASAP7_75t_SL g532 ( 
.A1(n_531),
.A2(n_14),
.B(n_1),
.C(n_2),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_0),
.C(n_1),
.Y(n_533)
);

O2A1O1Ixp33_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_0),
.B(n_1),
.C(n_514),
.Y(n_534)
);


endmodule