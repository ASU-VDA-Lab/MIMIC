module fake_jpeg_20220_n_209 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_209);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_209;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_34),
.Y(n_47)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_22),
.B1(n_14),
.B2(n_15),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_20),
.B1(n_23),
.B2(n_21),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_20),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_36),
.A2(n_18),
.B1(n_22),
.B2(n_14),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_38),
.B1(n_39),
.B2(n_36),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_18),
.B1(n_22),
.B2(n_15),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_28),
.A2(n_36),
.B1(n_35),
.B2(n_23),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_26),
.B1(n_21),
.B2(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_27),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_13),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_13),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_49),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_25),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_26),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_55),
.A2(n_62),
.B1(n_50),
.B2(n_40),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_17),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_61),
.Y(n_71)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_29),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_9),
.C(n_10),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_31),
.B1(n_19),
.B2(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_67),
.Y(n_78)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_69),
.Y(n_86)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

AND2x6_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_38),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_79),
.B(n_58),
.C(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_83),
.Y(n_103)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

AND2x6_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_37),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_85),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_52),
.B(n_29),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_55),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_87),
.A2(n_64),
.B1(n_63),
.B2(n_50),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_40),
.B(n_45),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_105),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_102),
.B1(n_107),
.B2(n_41),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_54),
.B1(n_50),
.B2(n_51),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_92),
.A2(n_94),
.B1(n_106),
.B2(n_77),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_60),
.B1(n_69),
.B2(n_31),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_45),
.B(n_66),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_95),
.A2(n_41),
.B(n_25),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_81),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_76),
.A2(n_72),
.B1(n_79),
.B2(n_75),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_45),
.B1(n_67),
.B2(n_42),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_56),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_75),
.A2(n_31),
.B1(n_42),
.B2(n_33),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_42),
.B1(n_29),
.B2(n_16),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_88),
.B(n_70),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_108),
.A2(n_117),
.B(n_126),
.Y(n_132)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_83),
.C(n_70),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_108),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_86),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_90),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_86),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_118),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_116),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_71),
.B(n_74),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_71),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_84),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_119),
.B(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_84),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_29),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_81),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_106),
.B1(n_94),
.B2(n_107),
.Y(n_128)
);

BUFx4f_ASAP7_75t_SL g124 ( 
.A(n_96),
.Y(n_124)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_129),
.B1(n_116),
.B2(n_125),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_123),
.A2(n_100),
.B1(n_89),
.B2(n_91),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_139),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_120),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_133),
.B(n_138),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_90),
.Y(n_135)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_117),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_103),
.C(n_105),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_143),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_97),
.B(n_96),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_109),
.A2(n_81),
.B(n_16),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_110),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_16),
.B1(n_7),
.B2(n_8),
.Y(n_142)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_121),
.C(n_126),
.Y(n_143)
);

NAND2x1_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_112),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_SL g169 ( 
.A(n_146),
.B(n_122),
.C(n_127),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_149),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_143),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_152),
.B1(n_158),
.B2(n_159),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_125),
.B1(n_122),
.B2(n_110),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_141),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_154),
.Y(n_164)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_132),
.Y(n_160)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_166),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_137),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_144),
.Y(n_181)
);

AOI31xp67_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_149),
.A3(n_135),
.B(n_168),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_118),
.C(n_129),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_140),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_138),
.C(n_135),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_152),
.C(n_156),
.Y(n_179)
);

OAI21x1_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_166),
.B(n_163),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_179),
.C(n_150),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_177),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_167),
.A2(n_158),
.B(n_157),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_161),
.A2(n_151),
.B1(n_159),
.B2(n_157),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_181),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_179),
.B(n_164),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_183),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_162),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_174),
.B(n_177),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_187),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_180),
.A2(n_163),
.B1(n_124),
.B2(n_7),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_174),
.B(n_6),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_5),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_124),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_195),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_191),
.A2(n_192),
.B(n_9),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_186),
.A2(n_124),
.B(n_6),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_194),
.A2(n_190),
.B(n_9),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_8),
.B1(n_11),
.B2(n_10),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_4),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_193),
.A2(n_8),
.B(n_11),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_198),
.A2(n_200),
.B(n_3),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_202),
.A2(n_12),
.B(n_1),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_204),
.A2(n_199),
.B(n_10),
.Y(n_205)
);

AOI321xp33_ASAP7_75t_L g207 ( 
.A1(n_205),
.A2(n_206),
.A3(n_203),
.B1(n_1),
.B2(n_2),
.C(n_0),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_207),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_2),
.Y(n_209)
);


endmodule