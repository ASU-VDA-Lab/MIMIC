module real_jpeg_18577_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_205;
wire n_110;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_202;
wire n_216;
wire n_167;
wire n_179;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_0),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_1),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_1),
.B(n_116),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_2),
.Y(n_116)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_2),
.Y(n_160)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_3),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_3),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_4),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_4),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_4),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_4),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_4),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_4),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_4),
.B(n_208),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_5),
.Y(n_120)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_5),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_6),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_6),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_6),
.B(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_6),
.A2(n_9),
.B1(n_102),
.B2(n_104),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_6),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_6),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_6),
.B(n_187),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_7),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_7),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_7),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_7),
.B(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_7),
.B(n_169),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g23 ( 
.A(n_8),
.B(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_8),
.B(n_138),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_9),
.Y(n_97)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_12),
.Y(n_141)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_12),
.Y(n_167)
);

BUFx4f_ASAP7_75t_L g210 ( 
.A(n_12),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_13),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_13),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_13),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_13),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_13),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_13),
.B(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_13),
.Y(n_136)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_14),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_146),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_144),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_89),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_18),
.B(n_89),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_56),
.C(n_74),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_19),
.A2(n_20),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_44),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_32),
.Y(n_21)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_22),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_28),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_23),
.B(n_28),
.Y(n_129)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_32),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_37),
.C(n_39),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_33),
.A2(n_39),
.B1(n_40),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_33),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

XOR2x1_ASAP7_75t_L g176 ( 
.A(n_37),
.B(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_42),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_44),
.B(n_124),
.C(n_125),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_45),
.B(n_49),
.C(n_52),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_51),
.B1(n_52),
.B2(n_55),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_49),
.A2(n_55),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_49),
.B(n_190),
.C(n_194),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_56),
.A2(n_74),
.B1(n_75),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_56),
.Y(n_224)
);

MAJx2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_65),
.C(n_67),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_57),
.B(n_65),
.Y(n_180)
);

XNOR2x1_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_62),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_62),
.Y(n_76)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_62),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_62),
.A2(n_185),
.B1(n_186),
.B2(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_67),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_72),
.Y(n_67)
);

AO22x1_ASAP7_75t_SL g171 ( 
.A1(n_68),
.A2(n_69),
.B1(n_72),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_72),
.Y(n_172)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_82),
.C(n_87),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_82),
.B1(n_87),
.B2(n_88),
.Y(n_77)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_80),
.B(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_82),
.Y(n_88)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_122),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_109),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_96),
.B(n_101),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.Y(n_109)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_117),
.B1(n_118),
.B2(n_121),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_115),
.Y(n_121)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_116),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_117),
.B(n_153),
.C(n_157),
.Y(n_175)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

XNOR2x1_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_137),
.B1(n_142),
.B2(n_143),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_135),
.Y(n_143)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

BUFx2_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_220),
.B(n_226),
.Y(n_147)
);

OAI21x1_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_181),
.B(n_219),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_173),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_150),
.B(n_173),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_161),
.C(n_171),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_151),
.B(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_161),
.A2(n_162),
.B1(n_171),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_168),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_163),
.B(n_168),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_179),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_175),
.B(n_176),
.C(n_179),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_213),
.B(n_218),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_199),
.B(n_212),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_189),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_189),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_206),
.B(n_211),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_204),
.Y(n_211)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_217),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_225),
.Y(n_220)
);

NOR2xp67_ASAP7_75t_SL g226 ( 
.A(n_221),
.B(n_225),
.Y(n_226)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);


endmodule