module real_jpeg_4090_n_31 (n_17, n_8, n_0, n_21, n_2, n_188, n_185, n_29, n_180, n_10, n_186, n_9, n_12, n_24, n_189, n_187, n_6, n_28, n_183, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_5, n_4, n_181, n_1, n_26, n_27, n_20, n_19, n_182, n_184, n_30, n_16, n_15, n_13, n_31);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_188;
input n_185;
input n_29;
input n_180;
input n_10;
input n_186;
input n_9;
input n_12;
input n_24;
input n_189;
input n_187;
input n_6;
input n_28;
input n_183;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_181;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_182;
input n_184;
input n_30;
input n_16;
input n_15;
input n_13;

output n_31;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_174;
wire n_87;
wire n_173;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_150;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_0),
.B(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_0),
.B(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_0),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_0),
.B(n_159),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_0),
.B(n_51),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_0),
.A2(n_48),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_1),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_2),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_3),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_4),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_4),
.B(n_145),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_5),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_5),
.B(n_67),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_6),
.Y(n_160)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_7),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_8),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_9),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_9),
.B(n_70),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_10),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_10),
.B(n_108),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_12),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_12),
.B(n_63),
.Y(n_131)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_13),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_14),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_16),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_17),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_18),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_19),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_19),
.B(n_81),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_20),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_21),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_21),
.B(n_84),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_22),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_23),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_23),
.B(n_162),
.Y(n_170)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_24),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_25),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_25),
.B(n_119),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_26),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_26),
.B(n_133),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_28),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_28),
.B(n_58),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_29),
.B(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_30),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_175),
.Y(n_31)
);

AO21x1_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_41),
.B(n_173),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_35),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_68),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_37),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_37),
.B(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_37),
.B(n_160),
.Y(n_159)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_39),
.B(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx11_ASAP7_75t_L g167 ( 
.A(n_40),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_49),
.B(n_172),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_48),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_43),
.B(n_48),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_45),
.B(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_45),
.B(n_146),
.Y(n_145)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_48),
.B(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_53),
.B(n_171),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_157),
.B(n_168),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_135),
.B(n_151),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_75),
.B(n_123),
.C(n_132),
.Y(n_55)
);

NOR4xp25_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.C(n_66),
.D(n_69),
.Y(n_56)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_60),
.B(n_134),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_66),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_82),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_104),
.Y(n_103)
);

OAI21x1_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_118),
.B(n_122),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_113),
.B(n_117),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_87),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_83),
.B(n_86),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_97),
.B(n_112),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_96),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_96),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_107),
.B(n_111),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_102),
.B(n_106),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_105),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_116),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B(n_129),
.C(n_130),
.D(n_131),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_143),
.C(n_147),
.Y(n_135)
);

A2O1A1O1Ixp25_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_147),
.B(n_152),
.C(n_155),
.D(n_156),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_138),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_153),
.B(n_154),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_150),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_180),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_181),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_182),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_183),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_184),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_185),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_186),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_187),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_188),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_189),
.Y(n_120)
);


endmodule