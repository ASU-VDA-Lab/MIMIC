module fake_jpeg_9995_n_314 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_5),
.B(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_10),
.B(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_41),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_36),
.Y(n_52)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_49),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_51),
.A2(n_24),
.B1(n_26),
.B2(n_32),
.Y(n_88)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_17),
.Y(n_70)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_34),
.A2(n_29),
.B1(n_30),
.B2(n_23),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_32),
.B1(n_22),
.B2(n_23),
.Y(n_67)
);

AND2x4_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_28),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_36),
.Y(n_87)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_34),
.A2(n_29),
.B1(n_24),
.B2(n_33),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_62),
.B1(n_26),
.B2(n_22),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_29),
.B1(n_24),
.B2(n_30),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_33),
.B1(n_19),
.B2(n_53),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_75),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_SL g72 ( 
.A1(n_57),
.A2(n_31),
.B(n_19),
.Y(n_72)
);

NOR2x1_ASAP7_75t_R g92 ( 
.A(n_72),
.B(n_31),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_46),
.B1(n_59),
.B2(n_52),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_37),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_40),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_84),
.Y(n_99)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_83),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_57),
.B(n_37),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_78),
.C(n_71),
.Y(n_102)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_39),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_61),
.B(n_37),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_17),
.Y(n_100)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_36),
.B(n_60),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_60),
.B1(n_18),
.B2(n_21),
.Y(n_108)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_92),
.A2(n_100),
.B(n_77),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_93),
.B(n_109),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_50),
.C(n_54),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_102),
.C(n_81),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_53),
.B1(n_46),
.B2(n_51),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_96),
.A2(n_103),
.B1(n_101),
.B2(n_100),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_108),
.B1(n_82),
.B2(n_65),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_48),
.B1(n_17),
.B2(n_36),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_27),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_25),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_117),
.Y(n_120)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_111),
.B(n_112),
.Y(n_140)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_91),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_25),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_119),
.A2(n_136),
.B1(n_138),
.B2(n_118),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_81),
.B1(n_87),
.B2(n_75),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_121),
.A2(n_128),
.B1(n_131),
.B2(n_137),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_122),
.B(n_124),
.C(n_133),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_75),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_135),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_87),
.C(n_69),
.Y(n_124)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_147),
.Y(n_151)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_127),
.B(n_130),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_67),
.B1(n_77),
.B2(n_69),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_123),
.B(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_90),
.B1(n_65),
.B2(n_79),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_58),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_134),
.B(n_144),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_68),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_97),
.A2(n_65),
.B1(n_80),
.B2(n_86),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_97),
.A2(n_80),
.B1(n_68),
.B2(n_82),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_141),
.B1(n_144),
.B2(n_112),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_98),
.A2(n_60),
.B1(n_18),
.B2(n_58),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_27),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_146),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_103),
.Y(n_167)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_21),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_145),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_27),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_150),
.B(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_154),
.B(n_155),
.Y(n_193)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_SL g184 ( 
.A(n_156),
.B(n_158),
.C(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_157),
.B(n_173),
.Y(n_205)
);

AO21x2_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_108),
.B(n_105),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_21),
.B1(n_27),
.B2(n_9),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_111),
.Y(n_160)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

OA21x2_ASAP7_75t_L g161 ( 
.A1(n_127),
.A2(n_130),
.B(n_129),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_164),
.B(n_21),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_118),
.Y(n_162)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_121),
.A2(n_95),
.B(n_92),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_169),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_104),
.C(n_18),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_118),
.Y(n_168)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_178),
.Y(n_203)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_125),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_120),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_174),
.Y(n_206)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_139),
.A2(n_92),
.B1(n_116),
.B2(n_93),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_177),
.A2(n_107),
.B1(n_124),
.B2(n_122),
.Y(n_180)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_180),
.B(n_186),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_172),
.A2(n_143),
.B1(n_94),
.B2(n_104),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_182),
.A2(n_192),
.B1(n_196),
.B2(n_197),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_176),
.C(n_178),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_190),
.B(n_159),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_158),
.A2(n_27),
.B1(n_21),
.B2(n_2),
.Y(n_191)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_192)
);

OAI22x1_ASAP7_75t_SL g195 ( 
.A1(n_158),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_201),
.B1(n_202),
.B2(n_179),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_158),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_158),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_199),
.Y(n_207)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_6),
.B(n_7),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_222),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_205),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_212),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_176),
.C(n_156),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_211),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_164),
.C(n_153),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_188),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_153),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_217),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_196),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_216),
.B(n_221),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_167),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_220),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_197),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_183),
.B(n_150),
.C(n_166),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_199),
.B(n_155),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_228),
.Y(n_241)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_181),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_224),
.B(n_200),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_195),
.A2(n_154),
.B1(n_152),
.B2(n_171),
.Y(n_225)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_226),
.B(n_191),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_201),
.Y(n_228)
);

INVx3_ASAP7_75t_SL g230 ( 
.A(n_184),
.Y(n_230)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_230),
.Y(n_246)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_194),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_230),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_247),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_236),
.B(n_202),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_213),
.A2(n_189),
.B1(n_182),
.B2(n_206),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_237),
.A2(n_229),
.B1(n_226),
.B2(n_220),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_239),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_166),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_244),
.C(n_222),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_193),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_245),
.Y(n_256)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_207),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_207),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_250),
.Y(n_265)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_254),
.Y(n_277)
);

INVx13_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_210),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_246),
.A2(n_219),
.B(n_213),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_266),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_240),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_185),
.Y(n_271)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_261),
.A2(n_262),
.B1(n_236),
.B2(n_237),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_240),
.A2(n_231),
.B1(n_215),
.B2(n_185),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_232),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_204),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_241),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_264),
.B(n_267),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_218),
.Y(n_266)
);

AOI221xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_229),
.B1(n_161),
.B2(n_194),
.C(n_177),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_266),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_271),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_275),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_280),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_257),
.B(n_187),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_227),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_276),
.B(n_279),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_165),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_262),
.A2(n_248),
.B1(n_238),
.B2(n_169),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_285),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_258),
.C(n_252),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_288),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_278),
.A2(n_256),
.B1(n_238),
.B2(n_260),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_290),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_265),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_234),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_254),
.C(n_234),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_208),
.C(n_280),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_235),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_293),
.C(n_298),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_235),
.C(n_265),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_291),
.A2(n_274),
.B(n_255),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_281),
.B(n_287),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_274),
.B(n_192),
.Y(n_297)
);

AO21x1_ASAP7_75t_L g304 ( 
.A1(n_297),
.A2(n_11),
.B(n_12),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_243),
.C(n_261),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_7),
.C(n_8),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_11),
.Y(n_303)
);

MAJx2_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_302),
.C(n_304),
.Y(n_308)
);

OAI21x1_ASAP7_75t_L g302 ( 
.A1(n_294),
.A2(n_9),
.B(n_11),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_303),
.A2(n_305),
.B(n_295),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_12),
.Y(n_305)
);

AO21x1_ASAP7_75t_L g310 ( 
.A1(n_307),
.A2(n_309),
.B(n_308),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_306),
.A2(n_299),
.B(n_13),
.Y(n_309)
);

NAND3xp33_ASAP7_75t_SL g311 ( 
.A(n_310),
.B(n_12),
.C(n_13),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_14),
.Y(n_312)
);

A2O1A1Ixp33_ASAP7_75t_SL g313 ( 
.A1(n_312),
.A2(n_14),
.B(n_15),
.C(n_302),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_14),
.Y(n_314)
);


endmodule