module fake_jpeg_27349_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_37),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_16),
.B(n_34),
.C(n_26),
.Y(n_54)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_43),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_31),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_60),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_54),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_58),
.B(n_63),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_31),
.B1(n_25),
.B2(n_20),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_61),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_38),
.B(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_31),
.B1(n_28),
.B2(n_17),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_65),
.A2(n_43),
.B1(n_26),
.B2(n_22),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_38),
.B(n_34),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_68),
.Y(n_98)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_69),
.B(n_71),
.Y(n_106)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_21),
.Y(n_71)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_77),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_80),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_82),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_57),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_85),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_23),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_86),
.A2(n_25),
.B1(n_22),
.B2(n_16),
.Y(n_127)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_87),
.A2(n_104),
.B1(n_108),
.B2(n_55),
.Y(n_120)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_89),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_23),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_92),
.B(n_95),
.Y(n_131)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_93),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_71),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_94),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_49),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_99),
.Y(n_124)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_102),
.B(n_105),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_55),
.A2(n_43),
.B1(n_17),
.B2(n_19),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_107),
.B(n_110),
.Y(n_111)
);

BUFx16f_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_63),
.B(n_34),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_53),
.B1(n_66),
.B2(n_69),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_112),
.A2(n_117),
.B1(n_118),
.B2(n_87),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_19),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_128),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_44),
.B1(n_56),
.B2(n_68),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_56),
.B1(n_40),
.B2(n_25),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_76),
.A2(n_26),
.B1(n_22),
.B2(n_40),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_132),
.B1(n_84),
.B2(n_82),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_18),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_84),
.A2(n_18),
.B1(n_47),
.B2(n_48),
.Y(n_132)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_141),
.B(n_143),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_106),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_142),
.B(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_144),
.A2(n_147),
.B1(n_42),
.B2(n_37),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_103),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_154),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_79),
.B1(n_109),
.B2(n_99),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_104),
.B(n_78),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_148),
.A2(n_169),
.B(n_116),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_109),
.Y(n_150)
);

AND2x6_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_9),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_165),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_133),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_152),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_158),
.B1(n_167),
.B2(n_119),
.Y(n_174)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_112),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_162),
.Y(n_185)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_111),
.B(n_131),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_157),
.B(n_161),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_73),
.B1(n_91),
.B2(n_77),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_140),
.Y(n_159)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_127),
.A2(n_30),
.B(n_33),
.C(n_3),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_126),
.B(n_123),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_30),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_124),
.Y(n_163)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_75),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_173),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_116),
.A2(n_96),
.B1(n_48),
.B2(n_47),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_134),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_168),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_48),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_135),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_171),
.Y(n_196)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_123),
.B(n_75),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_174),
.A2(n_143),
.B1(n_158),
.B2(n_160),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_178),
.A2(n_186),
.B(n_190),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_180),
.A2(n_159),
.B(n_156),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_27),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_181),
.B(n_167),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_135),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_182),
.B(n_37),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_139),
.B1(n_119),
.B2(n_136),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_183),
.A2(n_189),
.B1(n_191),
.B2(n_199),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_46),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_164),
.A2(n_119),
.B1(n_136),
.B2(n_114),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_149),
.B(n_148),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_114),
.B1(n_108),
.B2(n_46),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_201),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_198),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_149),
.A2(n_36),
.B1(n_33),
.B2(n_37),
.Y(n_199)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_202),
.B(n_206),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_141),
.B(n_27),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_207),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_152),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_204),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_144),
.A2(n_36),
.B1(n_37),
.B2(n_33),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_27),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_208),
.A2(n_219),
.B(n_186),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_217),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_145),
.Y(n_212)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_174),
.A2(n_146),
.B1(n_145),
.B2(n_151),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_215),
.A2(n_202),
.B1(n_186),
.B2(n_205),
.Y(n_248)
);

INVx13_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_175),
.B(n_154),
.Y(n_218)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_190),
.A2(n_165),
.B(n_171),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_225),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_193),
.C(n_178),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_181),
.C(n_200),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_224),
.A2(n_180),
.B(n_206),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_187),
.B(n_30),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_1),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_227),
.Y(n_238)
);

NOR3xp33_ASAP7_75t_SL g227 ( 
.A(n_195),
.B(n_159),
.C(n_37),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_229),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_185),
.B(n_1),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_183),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_232),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_188),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_184),
.B(n_9),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_234),
.Y(n_249)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_235),
.B(n_189),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_203),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_236),
.B(n_246),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_242),
.A2(n_250),
.B(n_219),
.Y(n_268)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_257),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_230),
.A2(n_216),
.B1(n_234),
.B2(n_220),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_247),
.A2(n_208),
.B1(n_210),
.B2(n_213),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_248),
.A2(n_224),
.B1(n_222),
.B2(n_221),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_176),
.Y(n_251)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_251),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_229),
.Y(n_252)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_252),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_256),
.C(n_235),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_201),
.Y(n_254)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_214),
.B(n_197),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_255),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_196),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_177),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_209),
.B(n_179),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_259),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_179),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_218),
.Y(n_261)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_261),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_231),
.Y(n_262)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_244),
.A2(n_241),
.B1(n_248),
.B2(n_216),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_263),
.A2(n_264),
.B1(n_240),
.B2(n_227),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_231),
.Y(n_267)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_268),
.A2(n_274),
.B(n_249),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_237),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_236),
.B(n_228),
.C(n_221),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_278),
.C(n_253),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_271),
.A2(n_279),
.B1(n_238),
.B2(n_237),
.Y(n_287)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_244),
.Y(n_272)
);

OAI21xp33_ASAP7_75t_SL g292 ( 
.A1(n_272),
.A2(n_252),
.B(n_240),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_250),
.A2(n_211),
.B(n_225),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_211),
.C(n_210),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_249),
.A2(n_217),
.B1(n_227),
.B2(n_194),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_260),
.C(n_265),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_247),
.B1(n_239),
.B2(n_241),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_281),
.A2(n_295),
.B1(n_265),
.B2(n_260),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_269),
.C(n_277),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_284),
.C(n_278),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_256),
.C(n_242),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_262),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_290),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_289),
.A2(n_293),
.B(n_261),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_294),
.Y(n_298)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_268),
.A2(n_238),
.B(n_194),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_272),
.A2(n_217),
.B1(n_199),
.B2(n_2),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_289),
.A2(n_266),
.B(n_274),
.Y(n_296)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_303),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_300),
.A2(n_307),
.B1(n_288),
.B2(n_286),
.Y(n_310)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_281),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_305),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_273),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_291),
.C(n_280),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_295),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_271),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_306),
.A2(n_283),
.B1(n_276),
.B2(n_275),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_293),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_313),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_312),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_302),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_318),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_3),
.C(n_4),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_308),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_323),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_300),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_319),
.B(n_299),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_325),
.A2(n_309),
.B(n_312),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_314),
.A2(n_306),
.B(n_307),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_317),
.Y(n_330)
);

AOI322xp5_ASAP7_75t_L g332 ( 
.A1(n_327),
.A2(n_323),
.A3(n_321),
.B1(n_324),
.B2(n_12),
.C1(n_7),
.C2(n_15),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_319),
.C(n_301),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_329),
.B(n_330),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_328),
.C(n_329),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_331),
.B(n_10),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_7),
.C(n_10),
.Y(n_335)
);

OAI221xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.C(n_15),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_15),
.B(n_11),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_11),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_14),
.B(n_336),
.Y(n_339)
);


endmodule