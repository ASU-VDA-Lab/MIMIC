module fake_jpeg_14628_n_63 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

AND2x2_ASAP7_75t_SL g26 ( 
.A(n_4),
.B(n_21),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

OR2x2_ASAP7_75t_SL g29 ( 
.A(n_3),
.B(n_13),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_0),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_30),
.A2(n_33),
.B1(n_27),
.B2(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_34),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_27),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_38),
.B(n_23),
.Y(n_44)
);

AOI22x1_ASAP7_75t_SL g38 ( 
.A1(n_30),
.A2(n_29),
.B1(n_16),
.B2(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_7),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_23),
.B1(n_24),
.B2(n_14),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_47)
);

AO22x1_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_28),
.B1(n_5),
.B2(n_6),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_7),
.B(n_8),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_49),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_35),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_50),
.C(n_51),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_9),
.B1(n_43),
.B2(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_48),
.B(n_45),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_37),
.C(n_36),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_50),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_58),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_59),
.A2(n_56),
.B(n_53),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_60),
.A2(n_52),
.B1(n_43),
.B2(n_19),
.Y(n_61)
);

OAI31xp33_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_10),
.A3(n_15),
.B(n_20),
.Y(n_62)
);

XOR2x2_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_22),
.Y(n_63)
);


endmodule