module fake_jpeg_450_n_107 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_107);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_43),
.Y(n_53)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_44),
.B(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_40),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_37),
.B1(n_34),
.B2(n_32),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_50),
.A2(n_52),
.B1(n_30),
.B2(n_31),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_37),
.B1(n_34),
.B2(n_32),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_60),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_57),
.B(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_53),
.B(n_1),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_2),
.Y(n_59)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_60),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_51),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_11),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_48),
.B(n_47),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_64),
.B(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_71),
.A2(n_40),
.B(n_43),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_4),
.C(n_5),
.Y(n_85)
);

CKINVDCx10_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_77),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_78),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_43),
.B1(n_3),
.B2(n_4),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_5),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_72),
.A2(n_2),
.B(n_3),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_6),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

NOR3xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_89),
.C(n_91),
.Y(n_94)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_6),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_7),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_92),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_96)
);

AO221x1_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_80),
.B1(n_76),
.B2(n_83),
.C(n_10),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

OA21x2_ASAP7_75t_SL g99 ( 
.A1(n_96),
.A2(n_86),
.B(n_88),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_93),
.C(n_88),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_98),
.C(n_84),
.Y(n_101)
);

OAI221xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_98),
.B1(n_97),
.B2(n_94),
.C(n_87),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_8),
.B(n_10),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_12),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_13),
.A3(n_15),
.B1(n_17),
.B2(n_20),
.C1(n_21),
.C2(n_23),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_24),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_26),
.Y(n_107)
);


endmodule