module real_jpeg_15901_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B(n_549),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_0),
.B(n_550),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_1),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_1),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_1),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_1),
.B(n_310),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_1),
.B(n_348),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_1),
.B(n_458),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_1),
.B(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_1),
.B(n_478),
.Y(n_477)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_2),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_2),
.Y(n_247)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_2),
.Y(n_281)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_2),
.Y(n_401)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_3),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_4),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_4),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_4),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_5),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_5),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_5),
.B(n_82),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_5),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_5),
.B(n_233),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_5),
.B(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_5),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_5),
.B(n_96),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_6),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_6),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_6),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_6),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_6),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_6),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_6),
.B(n_254),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_6),
.A2(n_15),
.B1(n_279),
.B2(n_282),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_6),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_7),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_7),
.B(n_54),
.Y(n_53)
);

INVxp33_ASAP7_75t_L g114 ( 
.A(n_7),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_7),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_7),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_7),
.B(n_290),
.Y(n_289)
);

AND2x4_ASAP7_75t_SL g307 ( 
.A(n_7),
.B(n_308),
.Y(n_307)
);

AND2x2_ASAP7_75t_SL g345 ( 
.A(n_7),
.B(n_96),
.Y(n_345)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_8),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_8),
.Y(n_297)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_8),
.Y(n_354)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_9),
.Y(n_191)
);

BUFx4f_ASAP7_75t_L g251 ( 
.A(n_9),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_9),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_10),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_10),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_10),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_10),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_10),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_11),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_11),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_11),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_11),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_11),
.B(n_60),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_11),
.B(n_189),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_11),
.B(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_12),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_12),
.Y(n_90)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_12),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_13),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_13),
.Y(n_203)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_13),
.Y(n_305)
);

BUFx5_ASAP7_75t_L g492 ( 
.A(n_13),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_14),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_14),
.B(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_14),
.B(n_237),
.Y(n_236)
);

AND2x2_ASAP7_75t_SL g259 ( 
.A(n_14),
.B(n_260),
.Y(n_259)
);

AND2x4_ASAP7_75t_SL g302 ( 
.A(n_14),
.B(n_303),
.Y(n_302)
);

AND2x4_ASAP7_75t_L g351 ( 
.A(n_14),
.B(n_352),
.Y(n_351)
);

AND2x4_ASAP7_75t_SL g404 ( 
.A(n_14),
.B(n_405),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_14),
.B(n_464),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_15),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_15),
.B(n_229),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_15),
.B(n_356),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_15),
.B(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_15),
.B(n_432),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_15),
.B(n_254),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_15),
.B(n_454),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_15),
.B(n_498),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_16),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_16),
.B(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_16),
.B(n_429),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_16),
.B(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_16),
.B(n_491),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_16),
.B(n_506),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_16),
.B(n_513),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_17),
.Y(n_143)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_18),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_18),
.Y(n_186)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_18),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_166),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_164),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_145),
.Y(n_22)
);

NOR2xp67_ASAP7_75t_R g165 ( 
.A(n_23),
.B(n_145),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_105),
.C(n_120),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_24),
.B(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_73),
.C(n_92),
.Y(n_24)
);

INVxp33_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_26),
.B(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_44),
.C(n_58),
.Y(n_26)
);

XNOR2x2_ASAP7_75t_SL g220 ( 
.A(n_27),
.B(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_39),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_29),
.A2(n_30),
.B1(n_108),
.B2(n_112),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_30),
.B(n_34),
.C(n_39),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_SL g123 ( 
.A(n_30),
.B(n_108),
.C(n_113),
.Y(n_123)
);

OR2x2_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_34),
.A2(n_35),
.B1(n_95),
.B2(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_35),
.B(n_95),
.C(n_97),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_38),
.Y(n_406)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_42),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_43),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_44),
.B(n_58),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.C(n_53),
.Y(n_44)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_45),
.B(n_53),
.Y(n_182)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_47),
.Y(n_350)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_48),
.Y(n_433)
);

XNOR2x1_ASAP7_75t_L g181 ( 
.A(n_49),
.B(n_182),
.Y(n_181)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_51),
.Y(n_308)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_59),
.B(n_64),
.C(n_70),
.Y(n_119)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_62),
.Y(n_206)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_62),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_70),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_69),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_74),
.B(n_92),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_75),
.B(n_85),
.C(n_91),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_85),
.B1(n_86),
.B2(n_91),
.Y(n_78)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_84),
.Y(n_313)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g288 ( 
.A(n_90),
.Y(n_288)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_102),
.C(n_104),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_93),
.A2(n_94),
.B1(n_211),
.B2(n_213),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_95),
.B(n_184),
.C(n_187),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_95),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_95),
.A2(n_188),
.B1(n_196),
.B2(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_97),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_97),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_97),
.A2(n_193),
.B1(n_289),
.B2(n_340),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_102),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_102),
.B(n_244),
.C(n_248),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_102),
.B(n_276),
.Y(n_275)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_104),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_104),
.B(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_104),
.A2(n_207),
.B1(n_209),
.B2(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_105),
.B(n_121),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_118),
.C(n_119),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_106),
.B(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_113),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_108),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_112),
.B1(n_129),
.B2(n_132),
.Y(n_128)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_112),
.B(n_125),
.C(n_129),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_118),
.B(n_119),
.Y(n_177)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_133),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_133),
.C(n_163),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_129),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_132),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_144),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_139),
.C(n_144),
.Y(n_147)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_143),
.Y(n_261)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_143),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_162),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_156),
.B2(n_157),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_214),
.B(n_545),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_168),
.A2(n_547),
.B(n_548),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_169),
.B(n_171),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.C(n_178),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_176),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_178),
.B(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_197),
.C(n_210),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_219),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.C(n_192),
.Y(n_180)
);

XNOR2x1_ASAP7_75t_L g323 ( 
.A(n_181),
.B(n_183),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_225),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_191),
.Y(n_290)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_191),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_192),
.Y(n_322)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_193),
.B(n_287),
.C(n_289),
.Y(n_286)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_210),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_207),
.C(n_209),
.Y(n_197)
);

XNOR2x1_ASAP7_75t_L g262 ( 
.A(n_198),
.B(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.C(n_204),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_199),
.B(n_204),
.Y(n_241)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_241),
.Y(n_240)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_207),
.Y(n_264)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_211),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_268),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_265),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g547 ( 
.A(n_217),
.B(n_265),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.C(n_222),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_218),
.B(n_220),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_222),
.B(n_367),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_242),
.C(n_262),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_223),
.B(n_320),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.C(n_240),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_224),
.B(n_227),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_232),
.C(n_235),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_228),
.A2(n_235),
.B1(n_236),
.B2(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_228),
.Y(n_364)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_232),
.B(n_363),
.Y(n_362)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_235),
.B(n_428),
.C(n_431),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_235),
.A2(n_236),
.B1(n_428),
.B2(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_238),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_239),
.Y(n_357)
);

XNOR2x2_ASAP7_75t_L g332 ( 
.A(n_240),
.B(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_242),
.B(n_262),
.Y(n_320)
);

MAJx2_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_252),
.C(n_258),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_243),
.B(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_248),
.Y(n_276)
);

INVx6_ASAP7_75t_L g499 ( 
.A(n_245),
.Y(n_499)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_251),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_253),
.B(n_259),
.Y(n_317)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_258),
.A2(n_259),
.B1(n_408),
.B2(n_409),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_259),
.B(n_403),
.C(n_408),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_261),
.Y(n_260)
);

AO21x2_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_372),
.B(n_542),
.Y(n_268)
);

NOR2xp67_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_365),
.Y(n_269)
);

AND2x2_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_326),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_271),
.B(n_326),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_318),
.Y(n_271)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_272),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_291),
.C(n_314),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_274),
.B(n_330),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.C(n_286),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_275),
.B(n_413),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_277),
.A2(n_278),
.B1(n_286),
.B2(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_278),
.A2(n_388),
.B(n_395),
.Y(n_387)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_281),
.Y(n_458)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_285),
.Y(n_430)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_286),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_287),
.B(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_289),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_292),
.A2(n_315),
.B1(n_316),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_292),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_306),
.C(n_309),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_293),
.B(n_360),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_298),
.C(n_302),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_294),
.A2(n_302),
.B1(n_385),
.B2(n_386),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_294),
.Y(n_386)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_298),
.B(n_384),
.Y(n_383)
);

INVx6_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_302),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_302),
.B(n_445),
.Y(n_444)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_306),
.A2(n_307),
.B1(n_309),
.B2(n_361),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_309),
.Y(n_361)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_319),
.A2(n_321),
.B1(n_324),
.B2(n_325),
.Y(n_318)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_319),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_321),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_321),
.Y(n_371)
);

XOR2x2_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_324),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_332),
.C(n_334),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_328),
.A2(n_329),
.B1(n_332),
.B2(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_332),
.Y(n_377)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_335),
.B(n_376),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_358),
.C(n_362),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_336),
.B(n_381),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_341),
.C(n_346),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XNOR2x1_ASAP7_75t_L g436 ( 
.A(n_338),
.B(n_437),
.Y(n_436)
);

XNOR2x1_ASAP7_75t_L g437 ( 
.A(n_341),
.B(n_346),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_345),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_342),
.B(n_345),
.Y(n_435)
);

NOR2x1_ASAP7_75t_R g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_351),
.C(n_355),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_347),
.B(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_351),
.A2(n_355),
.B1(n_424),
.B2(n_425),
.Y(n_423)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_351),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_351),
.B(n_487),
.C(n_489),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_351),
.A2(n_425),
.B1(n_489),
.B2(n_490),
.Y(n_502)
);

INVx8_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_353),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_354),
.Y(n_508)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_355),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_359),
.B(n_362),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_365),
.A2(n_543),
.B(n_544),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_368),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_366),
.B(n_368),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.C(n_371),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_438),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_378),
.C(n_415),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_375),
.B(n_379),
.Y(n_541)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_382),
.C(n_412),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_380),
.B(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_382),
.B(n_412),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_387),
.C(n_402),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_383),
.B(n_387),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_385),
.B(n_446),
.C(n_450),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_401),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_402),
.B(n_420),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g528 ( 
.A(n_403),
.B(n_529),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_407),
.Y(n_403)
);

XNOR2x1_ASAP7_75t_L g476 ( 
.A(n_404),
.B(n_407),
.Y(n_476)
);

CKINVDCx14_ASAP7_75t_R g496 ( 
.A(n_404),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_404),
.A2(n_496),
.B1(n_497),
.B2(n_510),
.Y(n_509)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_418),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_416),
.B(n_418),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_421),
.C(n_436),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_419),
.B(n_538),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_421),
.B(n_436),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_426),
.C(n_434),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_422),
.B(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_427),
.B(n_435),
.Y(n_524)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_428),
.Y(n_472)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_431),
.B(n_471),
.Y(n_470)
);

INVx5_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

NAND3xp33_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_540),
.C(n_541),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_440),
.A2(n_535),
.B(n_539),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_441),
.A2(n_520),
.B(n_534),
.Y(n_440)
);

OAI21x1_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_481),
.B(n_519),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_467),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_443),
.B(n_467),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_451),
.C(n_459),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_444),
.B(n_484),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_450),
.Y(n_445)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_451),
.A2(n_452),
.B1(n_459),
.B2(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_457),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_453),
.B(n_457),
.Y(n_488)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_456),
.Y(n_515)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_459),
.Y(n_485)
);

AO22x1_ASAP7_75t_SL g459 ( 
.A1(n_460),
.A2(n_463),
.B1(n_465),
.B2(n_466),
.Y(n_459)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_460),
.Y(n_465)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_463),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_465),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_466),
.B(n_512),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_473),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_470),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_469),
.B(n_473),
.C(n_533),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_470),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_475),
.Y(n_473)
);

MAJx2_ASAP7_75t_L g531 ( 
.A(n_474),
.B(n_476),
.C(n_477),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

AOI21x1_ASAP7_75t_L g481 ( 
.A1(n_482),
.A2(n_493),
.B(n_518),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_483),
.B(n_486),
.Y(n_482)
);

NOR2xp67_ASAP7_75t_SL g518 ( 
.A(n_483),
.B(n_486),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_487),
.A2(n_488),
.B1(n_501),
.B2(n_502),
.Y(n_500)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_494),
.A2(n_503),
.B(n_517),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_500),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_495),
.B(n_500),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_496),
.B(n_497),
.Y(n_495)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_497),
.Y(n_510)
);

INVx5_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_504),
.A2(n_511),
.B(n_516),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_509),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_505),
.B(n_509),
.Y(n_516)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_521),
.B(n_532),
.Y(n_520)
);

NOR2xp67_ASAP7_75t_SL g534 ( 
.A(n_521),
.B(n_532),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_522),
.A2(n_523),
.B1(n_525),
.B2(n_526),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_522),
.B(n_527),
.C(n_531),
.Y(n_536)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_527),
.A2(n_528),
.B1(n_530),
.B2(n_531),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

NOR2xp67_ASAP7_75t_L g535 ( 
.A(n_536),
.B(n_537),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_536),
.B(n_537),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);


endmodule