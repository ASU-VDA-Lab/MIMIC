module fake_ariane_524_n_1732 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1732);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1732;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1252;
wire n_1129;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_11),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_38),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_54),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_161),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_135),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_79),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_10),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_143),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_128),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_9),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_13),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_95),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_35),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_60),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_110),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_162),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_115),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_100),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_124),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_104),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_16),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_154),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_27),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_26),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_12),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_99),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_61),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_6),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_132),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_118),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_23),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_37),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_106),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_34),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_12),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_178),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_182),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_141),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_150),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_9),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_164),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_108),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_65),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_136),
.Y(n_229)
);

HB1xp67_ASAP7_75t_SL g230 ( 
.A(n_69),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_121),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_54),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_7),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_153),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_30),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_165),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_55),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_72),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_47),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_53),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_123),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_68),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_64),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_92),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_17),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_31),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_91),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_183),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_14),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_179),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_168),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_166),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_35),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_170),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_98),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_4),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_56),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_163),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_139),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_169),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_111),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_127),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_23),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_160),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_105),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_28),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_51),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_53),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_45),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_52),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_101),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_24),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_17),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_119),
.Y(n_274)
);

BUFx2_ASAP7_75t_SL g275 ( 
.A(n_48),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_1),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_3),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_85),
.Y(n_278)
);

BUFx2_ASAP7_75t_SL g279 ( 
.A(n_75),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_67),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_39),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_151),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_172),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_44),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_122),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_90),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_45),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_138),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_88),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_140),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_20),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_8),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_120),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_152),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_103),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_8),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_137),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_13),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_18),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_158),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_27),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_84),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_102),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_55),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_130),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_29),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_82),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_89),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_83),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_2),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_147),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_6),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_71),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_56),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_21),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_74),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_46),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_38),
.Y(n_318)
);

BUFx10_ASAP7_75t_L g319 ( 
.A(n_180),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_5),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_58),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_37),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_134),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_97),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_30),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_173),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_48),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_155),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_107),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_22),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_181),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_24),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_142),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_39),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_86),
.Y(n_335)
);

BUFx10_ASAP7_75t_L g336 ( 
.A(n_52),
.Y(n_336)
);

BUFx5_ASAP7_75t_L g337 ( 
.A(n_51),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_31),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_109),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_33),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_177),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_11),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_1),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_145),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_19),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_44),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_174),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_80),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_96),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_87),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_5),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_63),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_171),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_125),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_66),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_167),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_116),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_40),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_49),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_14),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_59),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_43),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_148),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_29),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_15),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_133),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_131),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_337),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_204),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_209),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_291),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_275),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_231),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_240),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_242),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_208),
.Y(n_376)
);

INVxp33_ASAP7_75t_SL g377 ( 
.A(n_191),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_187),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_191),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_204),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_327),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_221),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_221),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_187),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_266),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_266),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_258),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_258),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_339),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_339),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_338),
.B(n_0),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_208),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_281),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_281),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_341),
.Y(n_395)
);

NOR2xp67_ASAP7_75t_L g396 ( 
.A(n_239),
.B(n_217),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_347),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_347),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_337),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_240),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_239),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_350),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_337),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_337),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_350),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_354),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_354),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_366),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_337),
.B(n_0),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_366),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_337),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_337),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_194),
.Y(n_413)
);

NOR2xp67_ASAP7_75t_L g414 ( 
.A(n_217),
.B(n_2),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_194),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_213),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_319),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_220),
.Y(n_418)
);

INVxp33_ASAP7_75t_SL g419 ( 
.A(n_195),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_195),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_319),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_235),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_197),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_245),
.Y(n_424)
);

BUFx6f_ASAP7_75t_SL g425 ( 
.A(n_319),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_246),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_348),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_240),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_193),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_348),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_193),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_198),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_198),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_257),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_336),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_336),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_263),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_272),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_273),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_336),
.Y(n_440)
);

INVxp33_ASAP7_75t_L g441 ( 
.A(n_276),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_287),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_367),
.B(n_4),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_292),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_199),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_301),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_199),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_306),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_197),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_201),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_312),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_315),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_240),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_317),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_201),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_184),
.B(n_7),
.Y(n_456)
);

BUFx2_ASAP7_75t_SL g457 ( 
.A(n_189),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_205),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_325),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_206),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_330),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_205),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_206),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_210),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_249),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_369),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_368),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_399),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_389),
.B(n_230),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_390),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_380),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_189),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_406),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_368),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_410),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_413),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_400),
.B(n_249),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_417),
.B(n_421),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_403),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_404),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_458),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_378),
.B(n_320),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_411),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_464),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_412),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_453),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_453),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_374),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_374),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_374),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_415),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_396),
.B(n_320),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_428),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_429),
.B(n_192),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_417),
.B(n_421),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_371),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_429),
.B(n_295),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_380),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_428),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_382),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_382),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_409),
.A2(n_202),
.B(n_196),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_428),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_384),
.B(n_320),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_416),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_418),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_422),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_431),
.B(n_203),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_424),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_385),
.B(n_320),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_426),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_383),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_434),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_381),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_437),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_383),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_438),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_439),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_442),
.Y(n_519)
);

AND2x6_ASAP7_75t_L g520 ( 
.A(n_443),
.B(n_190),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_387),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_444),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_386),
.B(n_393),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_446),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_448),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_388),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_451),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_452),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_454),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_431),
.B(n_222),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_388),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_459),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_394),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_376),
.B(n_392),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_414),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_456),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_427),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_432),
.B(n_223),
.Y(n_538)
);

NAND3xp33_ASAP7_75t_L g539 ( 
.A(n_391),
.B(n_340),
.C(n_332),
.Y(n_539)
);

OR2x6_ASAP7_75t_L g540 ( 
.A(n_496),
.B(n_435),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_472),
.B(n_432),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_474),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_506),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_467),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_508),
.B(n_538),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_536),
.B(n_433),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_506),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_515),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_467),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_494),
.B(n_425),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_474),
.Y(n_551)
);

AND2x6_ASAP7_75t_L g552 ( 
.A(n_467),
.B(n_465),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_479),
.Y(n_553)
);

INVx5_ASAP7_75t_L g554 ( 
.A(n_474),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_506),
.Y(n_555)
);

NOR3xp33_ASAP7_75t_L g556 ( 
.A(n_539),
.B(n_346),
.C(n_232),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_515),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_536),
.B(n_433),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_474),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_530),
.B(n_445),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_468),
.B(n_445),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_490),
.Y(n_562)
);

INVx8_ASAP7_75t_L g563 ( 
.A(n_520),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_L g564 ( 
.A(n_478),
.B(n_447),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_474),
.Y(n_565)
);

INVxp33_ASAP7_75t_L g566 ( 
.A(n_469),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_490),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_509),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_490),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_SL g570 ( 
.A(n_514),
.B(n_373),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_488),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_479),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_468),
.B(n_447),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_534),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_483),
.B(n_450),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_488),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_484),
.B(n_423),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_509),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_509),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_517),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_465),
.B(n_372),
.Y(n_581)
);

AND2x6_ASAP7_75t_L g582 ( 
.A(n_515),
.B(n_190),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_474),
.Y(n_583)
);

AO21x2_ASAP7_75t_L g584 ( 
.A1(n_502),
.A2(n_228),
.B(n_226),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_481),
.B(n_370),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_517),
.Y(n_586)
);

BUFx8_ASAP7_75t_SL g587 ( 
.A(n_466),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_483),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_517),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_SL g590 ( 
.A1(n_539),
.A2(n_395),
.B1(n_398),
.B2(n_397),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_524),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_477),
.B(n_430),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_537),
.B(n_423),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_524),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_515),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_485),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_524),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_470),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_485),
.B(n_450),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_479),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_484),
.B(n_395),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_529),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_488),
.Y(n_603)
);

BUFx10_ASAP7_75t_L g604 ( 
.A(n_471),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_495),
.B(n_455),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_497),
.B(n_425),
.Y(n_606)
);

BUFx10_ASAP7_75t_L g607 ( 
.A(n_498),
.Y(n_607)
);

AND2x6_ASAP7_75t_L g608 ( 
.A(n_529),
.B(n_227),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_476),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_480),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_520),
.A2(n_365),
.B1(n_345),
.B2(n_461),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_491),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_529),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_520),
.A2(n_507),
.B1(n_511),
.B2(n_505),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_529),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_480),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_520),
.B(n_455),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_533),
.Y(n_618)
);

OR2x6_ASAP7_75t_L g619 ( 
.A(n_535),
.B(n_401),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_477),
.B(n_420),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_477),
.B(n_449),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_500),
.B(n_397),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_520),
.B(n_460),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_533),
.B(n_425),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_532),
.B(n_460),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_511),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_533),
.B(n_463),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_513),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_533),
.B(n_463),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_532),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_513),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_532),
.B(n_373),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_486),
.Y(n_633)
);

BUFx10_ASAP7_75t_L g634 ( 
.A(n_501),
.Y(n_634)
);

INVxp67_ASAP7_75t_SL g635 ( 
.A(n_532),
.Y(n_635)
);

INVx8_ASAP7_75t_L g636 ( 
.A(n_520),
.Y(n_636)
);

OR2x6_ASAP7_75t_L g637 ( 
.A(n_535),
.B(n_462),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_518),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_520),
.A2(n_377),
.B1(n_419),
.B2(n_379),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_518),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_519),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_523),
.B(n_375),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_477),
.B(n_247),
.Y(n_643)
);

BUFx10_ASAP7_75t_L g644 ( 
.A(n_512),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_473),
.Y(n_645)
);

AO22x2_ASAP7_75t_L g646 ( 
.A1(n_522),
.A2(n_186),
.B1(n_233),
.B2(n_267),
.Y(n_646)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_510),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_522),
.B(n_375),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_516),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_525),
.B(n_250),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_489),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_486),
.Y(n_652)
);

NAND2xp33_ASAP7_75t_L g653 ( 
.A(n_527),
.B(n_295),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_528),
.B(n_260),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_510),
.Y(n_655)
);

INVx5_ASAP7_75t_L g656 ( 
.A(n_482),
.Y(n_656)
);

AND2x6_ASAP7_75t_L g657 ( 
.A(n_482),
.B(n_227),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_504),
.B(n_324),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_502),
.B(n_264),
.Y(n_659)
);

BUFx10_ASAP7_75t_L g660 ( 
.A(n_521),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_504),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_493),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_510),
.B(n_278),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_493),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_510),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_492),
.A2(n_313),
.B1(n_329),
.B2(n_279),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_499),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_503),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_503),
.Y(n_669)
);

INVxp33_ASAP7_75t_L g670 ( 
.A(n_469),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_492),
.B(n_288),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_492),
.B(n_303),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_487),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_487),
.B(n_305),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_545),
.B(n_627),
.Y(n_675)
);

NOR3xp33_ASAP7_75t_L g676 ( 
.A(n_649),
.B(n_531),
.C(n_526),
.Y(n_676)
);

A2O1A1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_545),
.A2(n_358),
.B(n_210),
.C(n_296),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_667),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_627),
.B(n_356),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_593),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_585),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_560),
.B(n_185),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_614),
.B(n_356),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_629),
.B(n_357),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_629),
.B(n_357),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_620),
.B(n_436),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_673),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_614),
.B(n_361),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_550),
.B(n_361),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_546),
.B(n_216),
.Y(n_690)
);

O2A1O1Ixp5_ASAP7_75t_L g691 ( 
.A1(n_617),
.A2(n_333),
.B(n_309),
.C(n_363),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_552),
.A2(n_407),
.B1(n_402),
.B2(n_405),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_550),
.B(n_402),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_581),
.B(n_405),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_667),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_635),
.B(n_408),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_635),
.B(n_408),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_548),
.B(n_307),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_558),
.B(n_219),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_639),
.A2(n_541),
.B1(n_623),
.B2(n_575),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_673),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_641),
.B(n_225),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_641),
.B(n_237),
.Y(n_703)
);

O2A1O1Ixp5_ASAP7_75t_L g704 ( 
.A1(n_659),
.A2(n_625),
.B(n_557),
.C(n_595),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_573),
.A2(n_557),
.B(n_548),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_605),
.B(n_253),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_648),
.B(n_256),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_648),
.B(n_268),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_630),
.B(n_269),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_544),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_595),
.B(n_326),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_561),
.B(n_270),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_592),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_611),
.A2(n_329),
.B1(n_313),
.B2(n_358),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_588),
.Y(n_715)
);

O2A1O1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_561),
.A2(n_328),
.B(n_355),
.C(n_296),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_552),
.A2(n_234),
.B1(n_262),
.B2(n_261),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_596),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_552),
.B(n_277),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_655),
.B(n_284),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_602),
.A2(n_224),
.B(n_316),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_587),
.Y(n_722)
);

NOR2x1p5_ASAP7_75t_L g723 ( 
.A(n_622),
.B(n_601),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_549),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_596),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_645),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_655),
.B(n_298),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_602),
.B(n_200),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_613),
.B(n_200),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_669),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_665),
.B(n_299),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_665),
.B(n_304),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_615),
.B(n_200),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_599),
.B(n_310),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_615),
.B(n_200),
.Y(n_735)
);

OR2x6_ASAP7_75t_L g736 ( 
.A(n_577),
.B(n_475),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_563),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_549),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_639),
.A2(n_211),
.B1(n_215),
.B2(n_214),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_611),
.A2(n_359),
.B1(n_360),
.B2(n_440),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_626),
.B(n_628),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_598),
.Y(n_742)
);

NOR3xp33_ASAP7_75t_L g743 ( 
.A(n_632),
.B(n_359),
.C(n_360),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_631),
.B(n_314),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_599),
.B(n_318),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_556),
.A2(n_666),
.B1(n_646),
.B2(n_636),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_638),
.B(n_322),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_609),
.B(n_334),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_669),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_625),
.B(n_342),
.Y(n_750)
);

NAND3xp33_ASAP7_75t_L g751 ( 
.A(n_570),
.B(n_364),
.C(n_362),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_553),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_642),
.B(n_343),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_604),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_640),
.B(n_351),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_563),
.B(n_207),
.Y(n_756)
);

AND2x6_ASAP7_75t_L g757 ( 
.A(n_624),
.B(n_229),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_563),
.B(n_636),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_636),
.B(n_207),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_664),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_604),
.Y(n_761)
);

AOI221xp5_ASAP7_75t_L g762 ( 
.A1(n_556),
.A2(n_353),
.B1(n_352),
.B2(n_349),
.C(n_344),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_L g763 ( 
.A1(n_574),
.A2(n_271),
.B1(n_331),
.B2(n_323),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_540),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_661),
.B(n_188),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_651),
.B(n_207),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_672),
.B(n_212),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_542),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_662),
.B(n_207),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_662),
.B(n_207),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_672),
.B(n_218),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_574),
.B(n_16),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_632),
.B(n_18),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_624),
.B(n_236),
.Y(n_774)
);

NOR3xp33_ASAP7_75t_L g775 ( 
.A(n_564),
.B(n_297),
.C(n_238),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_647),
.B(n_19),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_621),
.B(n_20),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_606),
.A2(n_280),
.B1(n_321),
.B2(n_311),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_650),
.A2(n_274),
.B(n_308),
.C(n_302),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_572),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_658),
.B(n_606),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_618),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_600),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_666),
.B(n_259),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_668),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_619),
.B(n_647),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_619),
.B(n_25),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_633),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_600),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_571),
.B(n_265),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_571),
.B(n_255),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_540),
.B(n_28),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_653),
.A2(n_32),
.B(n_33),
.C(n_36),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_540),
.B(n_36),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_576),
.B(n_282),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_576),
.B(n_254),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_612),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_603),
.B(n_283),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_657),
.A2(n_252),
.B1(n_300),
.B2(n_294),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_657),
.A2(n_251),
.B1(n_293),
.B2(n_290),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_656),
.B(n_618),
.Y(n_801)
);

INVx8_ASAP7_75t_L g802 ( 
.A(n_657),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_603),
.B(n_244),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_542),
.B(n_207),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_650),
.B(n_248),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_542),
.B(n_207),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_657),
.A2(n_289),
.B1(n_286),
.B2(n_285),
.Y(n_807)
);

AO21x1_ASAP7_75t_L g808 ( 
.A1(n_700),
.A2(n_659),
.B(n_674),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_675),
.B(n_643),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_L g810 ( 
.A1(n_704),
.A2(n_610),
.B(n_616),
.Y(n_810)
);

AO21x1_ASAP7_75t_L g811 ( 
.A1(n_773),
.A2(n_674),
.B(n_543),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_693),
.B(n_577),
.Y(n_812)
);

INVx4_ASAP7_75t_L g813 ( 
.A(n_802),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_682),
.B(n_643),
.Y(n_814)
);

AO21x1_ASAP7_75t_L g815 ( 
.A1(n_773),
.A2(n_781),
.B(n_684),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_679),
.A2(n_590),
.B1(n_656),
.B2(n_586),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_682),
.B(n_656),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_690),
.A2(n_547),
.B(n_555),
.C(n_568),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_728),
.A2(n_616),
.B(n_584),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_786),
.B(n_607),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_737),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_760),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_680),
.B(n_634),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_729),
.A2(n_584),
.B(n_578),
.Y(n_824)
);

AOI33xp33_ASAP7_75t_L g825 ( 
.A1(n_753),
.A2(n_590),
.A3(n_579),
.B1(n_580),
.B2(n_589),
.B3(n_591),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_705),
.A2(n_583),
.B(n_542),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_696),
.B(n_644),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_690),
.B(n_656),
.Y(n_828)
);

BUFx2_ASAP7_75t_L g829 ( 
.A(n_742),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_768),
.Y(n_830)
);

O2A1O1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_677),
.A2(n_654),
.B(n_594),
.C(n_597),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_797),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_685),
.A2(n_619),
.B1(n_637),
.B2(n_559),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_697),
.B(n_660),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_681),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_677),
.A2(n_654),
.B(n_671),
.C(n_663),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_733),
.A2(n_583),
.B(n_551),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_707),
.B(n_657),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_708),
.B(n_671),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_735),
.A2(n_711),
.B(n_698),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_691),
.A2(n_735),
.B(n_730),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_698),
.A2(n_565),
.B(n_559),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_779),
.A2(n_663),
.B(n_637),
.C(n_562),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_785),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_678),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_689),
.B(n_608),
.Y(n_846)
);

OAI21xp5_ASAP7_75t_L g847 ( 
.A1(n_749),
.A2(n_567),
.B(n_569),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_750),
.B(n_582),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_774),
.A2(n_554),
.B(n_652),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_695),
.A2(n_608),
.B(n_582),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_712),
.B(n_582),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_712),
.B(n_582),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_734),
.B(n_582),
.Y(n_853)
);

BUFx10_ASAP7_75t_L g854 ( 
.A(n_726),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_734),
.B(n_608),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_745),
.B(n_608),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_741),
.A2(n_554),
.B(n_652),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_766),
.A2(n_243),
.B(n_241),
.Y(n_858)
);

INVx1_ASAP7_75t_SL g859 ( 
.A(n_694),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_766),
.A2(n_335),
.B(n_229),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_745),
.B(n_670),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_769),
.A2(n_335),
.B(n_229),
.Y(n_862)
);

INVx5_ASAP7_75t_L g863 ( 
.A(n_802),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_706),
.B(n_566),
.Y(n_864)
);

NAND3xp33_ASAP7_75t_SL g865 ( 
.A(n_676),
.B(n_40),
.C(n_41),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_686),
.B(n_41),
.Y(n_866)
);

AO22x1_ASAP7_75t_L g867 ( 
.A1(n_686),
.A2(n_229),
.B1(n_335),
.B2(n_46),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_754),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_706),
.A2(n_776),
.B(n_739),
.C(n_716),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_769),
.A2(n_42),
.B(n_43),
.Y(n_870)
);

AOI21x1_ASAP7_75t_L g871 ( 
.A1(n_756),
.A2(n_94),
.B(n_175),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_770),
.A2(n_50),
.B(n_57),
.Y(n_872)
);

NOR2xp67_ASAP7_75t_L g873 ( 
.A(n_722),
.B(n_754),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_805),
.A2(n_714),
.B1(n_782),
.B2(n_699),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_776),
.A2(n_62),
.B(n_70),
.C(n_73),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_770),
.A2(n_76),
.B(n_77),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_714),
.B(n_78),
.Y(n_877)
);

AO21x1_ASAP7_75t_L g878 ( 
.A1(n_804),
.A2(n_806),
.B(n_793),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_709),
.A2(n_81),
.B(n_93),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_692),
.B(n_764),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_782),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_748),
.Y(n_882)
);

NOR2x1_ASAP7_75t_L g883 ( 
.A(n_761),
.B(n_117),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_723),
.B(n_126),
.Y(n_884)
);

AOI21xp33_ASAP7_75t_L g885 ( 
.A1(n_740),
.A2(n_784),
.B(n_746),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_804),
.A2(n_129),
.B(n_144),
.Y(n_886)
);

O2A1O1Ixp5_ASAP7_75t_L g887 ( 
.A1(n_767),
.A2(n_146),
.B(n_149),
.C(n_157),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_737),
.B(n_159),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_752),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_715),
.A2(n_725),
.B1(n_718),
.B2(n_771),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_687),
.B(n_701),
.Y(n_891)
);

AOI33xp33_ASAP7_75t_L g892 ( 
.A1(n_772),
.A2(n_740),
.A3(n_792),
.B1(n_794),
.B2(n_777),
.B3(n_787),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_713),
.B(n_787),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_746),
.B(n_702),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_703),
.B(n_778),
.Y(n_895)
);

INVx4_ASAP7_75t_L g896 ( 
.A(n_737),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_743),
.A2(n_762),
.B1(n_683),
.B2(n_688),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_744),
.B(n_755),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_768),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_801),
.A2(n_798),
.B(n_790),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_747),
.B(n_720),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_727),
.B(n_731),
.Y(n_902)
);

AO21x1_ASAP7_75t_L g903 ( 
.A1(n_806),
.A2(n_759),
.B(n_688),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_801),
.A2(n_795),
.B(n_791),
.Y(n_904)
);

NAND2x1p5_ASAP7_75t_L g905 ( 
.A(n_737),
.B(n_758),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_736),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_796),
.A2(n_803),
.B(n_765),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_732),
.B(n_683),
.Y(n_908)
);

NAND3xp33_ASAP7_75t_L g909 ( 
.A(n_763),
.B(n_751),
.C(n_775),
.Y(n_909)
);

AOI33xp33_ASAP7_75t_L g910 ( 
.A1(n_717),
.A2(n_807),
.A3(n_800),
.B1(n_799),
.B2(n_789),
.B3(n_783),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_780),
.B(n_789),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_719),
.A2(n_757),
.B1(n_721),
.B2(n_736),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_710),
.A2(n_724),
.B(n_738),
.C(n_788),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_757),
.A2(n_704),
.B(n_675),
.Y(n_914)
);

NOR2x1p5_ASAP7_75t_SL g915 ( 
.A(n_757),
.B(n_678),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_757),
.A2(n_675),
.B(n_705),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_757),
.B(n_675),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_675),
.B(n_545),
.Y(n_918)
);

BUFx12f_ASAP7_75t_L g919 ( 
.A(n_742),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_675),
.A2(n_705),
.B(n_728),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_675),
.A2(n_679),
.B1(n_685),
.B2(n_684),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_742),
.Y(n_922)
);

O2A1O1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_675),
.A2(n_677),
.B(n_546),
.C(n_558),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_675),
.A2(n_679),
.B1(n_685),
.B2(n_684),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_680),
.B(n_593),
.Y(n_925)
);

A2O1A1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_675),
.A2(n_773),
.B(n_545),
.C(n_682),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_768),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_675),
.B(n_545),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_714),
.A2(n_746),
.B1(n_740),
.B2(n_666),
.Y(n_929)
);

AO22x1_ASAP7_75t_L g930 ( 
.A1(n_742),
.A2(n_380),
.B1(n_383),
.B2(n_382),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_675),
.A2(n_773),
.B(n_545),
.C(n_682),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_675),
.A2(n_729),
.B(n_728),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_675),
.A2(n_729),
.B(n_728),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_675),
.B(n_545),
.Y(n_934)
);

OAI321xp33_ASAP7_75t_L g935 ( 
.A1(n_675),
.A2(n_740),
.A3(n_714),
.B1(n_639),
.B2(n_700),
.C(n_391),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_768),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_786),
.B(n_675),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_675),
.A2(n_729),
.B(n_728),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_675),
.B(n_380),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_786),
.B(n_675),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_675),
.B(n_545),
.Y(n_941)
);

NOR2x1_ASAP7_75t_L g942 ( 
.A(n_754),
.B(n_761),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_737),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_704),
.A2(n_675),
.B(n_691),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_675),
.A2(n_729),
.B(n_728),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_737),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_675),
.A2(n_679),
.B1(n_685),
.B2(n_684),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_680),
.B(n_593),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_675),
.A2(n_729),
.B(n_728),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_675),
.A2(n_729),
.B(n_728),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_675),
.A2(n_773),
.B(n_545),
.C(n_682),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_737),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_675),
.B(n_545),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_680),
.B(n_593),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_737),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_926),
.A2(n_951),
.B(n_931),
.Y(n_956)
);

O2A1O1Ixp5_ASAP7_75t_L g957 ( 
.A1(n_808),
.A2(n_815),
.B(n_811),
.C(n_869),
.Y(n_957)
);

BUFx8_ASAP7_75t_SL g958 ( 
.A(n_919),
.Y(n_958)
);

OAI21x1_ASAP7_75t_L g959 ( 
.A1(n_819),
.A2(n_824),
.B(n_826),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_822),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_925),
.B(n_948),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_934),
.A2(n_953),
.B(n_941),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_932),
.A2(n_938),
.B(n_933),
.Y(n_963)
);

NOR2x1_ASAP7_75t_L g964 ( 
.A(n_868),
.B(n_829),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_809),
.B(n_814),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_832),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_921),
.B(n_924),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_830),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_954),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_947),
.B(n_894),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_938),
.A2(n_949),
.B(n_945),
.Y(n_971)
);

A2O1A1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_935),
.A2(n_939),
.B(n_923),
.C(n_897),
.Y(n_972)
);

OAI21x1_ASAP7_75t_L g973 ( 
.A1(n_819),
.A2(n_824),
.B(n_810),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_864),
.B(n_861),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_895),
.A2(n_839),
.B(n_898),
.C(n_901),
.Y(n_975)
);

AOI21x1_ASAP7_75t_SL g976 ( 
.A1(n_902),
.A2(n_817),
.B(n_828),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_945),
.A2(n_950),
.B(n_949),
.Y(n_977)
);

BUFx12f_ASAP7_75t_L g978 ( 
.A(n_854),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_950),
.A2(n_914),
.B(n_916),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_929),
.B(n_937),
.Y(n_980)
);

CKINVDCx20_ASAP7_75t_R g981 ( 
.A(n_854),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_859),
.B(n_882),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_940),
.B(n_825),
.Y(n_983)
);

INVxp67_ASAP7_75t_L g984 ( 
.A(n_866),
.Y(n_984)
);

INVx4_ASAP7_75t_L g985 ( 
.A(n_863),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_812),
.B(n_893),
.Y(n_986)
);

AOI21x1_ASAP7_75t_L g987 ( 
.A1(n_900),
.A2(n_904),
.B(n_907),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_836),
.A2(n_843),
.B(n_827),
.C(n_834),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_844),
.A2(n_909),
.B1(n_874),
.B2(n_877),
.Y(n_989)
);

AO21x1_ASAP7_75t_L g990 ( 
.A1(n_917),
.A2(n_904),
.B(n_900),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_846),
.A2(n_849),
.B(n_840),
.Y(n_991)
);

NAND2xp33_ASAP7_75t_L g992 ( 
.A(n_863),
.B(n_830),
.Y(n_992)
);

INVx5_ASAP7_75t_L g993 ( 
.A(n_863),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_830),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_823),
.Y(n_995)
);

AO21x1_ASAP7_75t_L g996 ( 
.A1(n_848),
.A2(n_856),
.B(n_855),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_908),
.B(n_845),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_885),
.B(n_889),
.Y(n_998)
);

NOR2x1_ASAP7_75t_L g999 ( 
.A(n_873),
.B(n_942),
.Y(n_999)
);

AO31x2_ASAP7_75t_L g1000 ( 
.A1(n_903),
.A2(n_878),
.A3(n_816),
.B(n_818),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_835),
.B(n_892),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_930),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_833),
.B(n_863),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_906),
.B(n_884),
.Y(n_1004)
);

AO31x2_ASAP7_75t_L g1005 ( 
.A1(n_857),
.A2(n_890),
.A3(n_913),
.B(n_860),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_944),
.A2(n_838),
.B(n_853),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_911),
.B(n_851),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_891),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_841),
.A2(n_831),
.B(n_837),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_880),
.B(n_820),
.Y(n_1010)
);

OA21x2_ASAP7_75t_L g1011 ( 
.A1(n_860),
.A2(n_862),
.B(n_879),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_852),
.B(n_910),
.Y(n_1012)
);

AOI221x1_ASAP7_75t_L g1013 ( 
.A1(n_879),
.A2(n_870),
.B1(n_872),
.B2(n_862),
.C(n_865),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_899),
.B(n_936),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_842),
.A2(n_850),
.B(n_847),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_876),
.A2(n_875),
.B(n_886),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_871),
.A2(n_905),
.B(n_887),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_905),
.A2(n_872),
.B(n_888),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_912),
.A2(n_936),
.B1(n_927),
.B2(n_899),
.Y(n_1019)
);

AO31x2_ASAP7_75t_L g1020 ( 
.A1(n_881),
.A2(n_858),
.A3(n_915),
.B(n_896),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_899),
.B(n_936),
.Y(n_1021)
);

NAND2xp33_ASAP7_75t_L g1022 ( 
.A(n_927),
.B(n_955),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_927),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_858),
.A2(n_883),
.B(n_955),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_821),
.B(n_952),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_867),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_821),
.A2(n_943),
.B(n_946),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_943),
.A2(n_952),
.B(n_946),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_896),
.A2(n_931),
.B(n_926),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_918),
.B(n_928),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_819),
.A2(n_824),
.B(n_826),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_SL g1032 ( 
.A1(n_815),
.A2(n_811),
.B(n_808),
.Y(n_1032)
);

AOI22x1_ASAP7_75t_L g1033 ( 
.A1(n_907),
.A2(n_904),
.B1(n_900),
.B2(n_920),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_925),
.B(n_948),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_918),
.B(n_928),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_819),
.A2(n_824),
.B(n_826),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_939),
.B(n_380),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_918),
.B(n_928),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_925),
.B(n_948),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_813),
.Y(n_1040)
);

INVx4_ASAP7_75t_L g1041 ( 
.A(n_863),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_863),
.B(n_786),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_939),
.B(n_786),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_819),
.A2(n_824),
.B(n_826),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_819),
.A2(n_824),
.B(n_826),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_918),
.A2(n_934),
.B(n_928),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_SL g1047 ( 
.A1(n_815),
.A2(n_811),
.B(n_808),
.Y(n_1047)
);

INVxp67_ASAP7_75t_L g1048 ( 
.A(n_832),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_918),
.A2(n_934),
.B(n_928),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_918),
.A2(n_934),
.B(n_928),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_918),
.A2(n_675),
.B1(n_953),
.B2(n_934),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_926),
.A2(n_931),
.B(n_951),
.C(n_935),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_926),
.A2(n_951),
.B(n_931),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_819),
.A2(n_824),
.B(n_826),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_868),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_918),
.B(n_928),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_918),
.A2(n_934),
.B(n_928),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_926),
.A2(n_951),
.B(n_931),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_918),
.B(n_928),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_926),
.A2(n_951),
.B(n_931),
.Y(n_1060)
);

NOR2xp67_ASAP7_75t_L g1061 ( 
.A(n_922),
.B(n_726),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_819),
.A2(n_824),
.B(n_826),
.Y(n_1062)
);

BUFx4f_ASAP7_75t_L g1063 ( 
.A(n_919),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_918),
.B(n_928),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_868),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_918),
.A2(n_934),
.B(n_928),
.Y(n_1066)
);

O2A1O1Ixp5_ASAP7_75t_L g1067 ( 
.A1(n_808),
.A2(n_931),
.B(n_951),
.C(n_926),
.Y(n_1067)
);

AO31x2_ASAP7_75t_L g1068 ( 
.A1(n_811),
.A2(n_808),
.A3(n_815),
.B(n_903),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_813),
.Y(n_1069)
);

AOI21x1_ASAP7_75t_SL g1070 ( 
.A1(n_918),
.A2(n_675),
.B(n_679),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_819),
.A2(n_824),
.B(n_826),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_819),
.A2(n_824),
.B(n_826),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_819),
.A2(n_824),
.B(n_826),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_918),
.A2(n_934),
.B(n_928),
.Y(n_1074)
);

AOI21xp33_ASAP7_75t_L g1075 ( 
.A1(n_935),
.A2(n_931),
.B(n_926),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_830),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_926),
.A2(n_931),
.B(n_951),
.C(n_935),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_918),
.A2(n_934),
.B(n_928),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_918),
.A2(n_934),
.B(n_928),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_819),
.A2(n_824),
.B(n_826),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_819),
.A2(n_824),
.B(n_826),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1051),
.B(n_965),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_SL g1083 ( 
.A(n_1063),
.B(n_1065),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_967),
.A2(n_972),
.B(n_1037),
.C(n_1077),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_985),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_961),
.B(n_1034),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_960),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_985),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_1042),
.B(n_993),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1039),
.B(n_974),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_1055),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_1041),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_958),
.Y(n_1093)
);

NOR2xp67_ASAP7_75t_L g1094 ( 
.A(n_1048),
.B(n_1061),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_988),
.A2(n_975),
.B(n_970),
.C(n_1079),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_962),
.A2(n_1050),
.B(n_1049),
.C(n_1078),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_979),
.A2(n_1052),
.B(n_1053),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_956),
.A2(n_1053),
.B(n_1058),
.Y(n_1098)
);

NOR2xp67_ASAP7_75t_L g1099 ( 
.A(n_966),
.B(n_969),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_986),
.B(n_982),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1001),
.B(n_1002),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_964),
.Y(n_1102)
);

NOR2x1_ASAP7_75t_SL g1103 ( 
.A(n_1003),
.B(n_968),
.Y(n_1103)
);

NAND2xp33_ASAP7_75t_L g1104 ( 
.A(n_1030),
.B(n_1035),
.Y(n_1104)
);

NAND3xp33_ASAP7_75t_L g1105 ( 
.A(n_956),
.B(n_1058),
.C(n_1060),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1030),
.A2(n_1064),
.B1(n_1038),
.B2(n_1059),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_978),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_981),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1008),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_968),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_995),
.Y(n_1111)
);

NOR2x1_ASAP7_75t_L g1112 ( 
.A(n_1043),
.B(n_999),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1056),
.B(n_1059),
.Y(n_1113)
);

CKINVDCx11_ASAP7_75t_R g1114 ( 
.A(n_968),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_1064),
.A2(n_1046),
.B1(n_1057),
.B2(n_1066),
.Y(n_1115)
);

OR2x2_ASAP7_75t_L g1116 ( 
.A(n_984),
.B(n_1074),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_1040),
.B(n_1069),
.Y(n_1117)
);

INVx1_ASAP7_75t_SL g1118 ( 
.A(n_1004),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_965),
.B(n_980),
.Y(n_1119)
);

NOR2xp67_ASAP7_75t_SL g1120 ( 
.A(n_1040),
.B(n_1069),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1075),
.A2(n_971),
.B(n_977),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_994),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_994),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_1010),
.B(n_1026),
.Y(n_1124)
);

INVx3_ASAP7_75t_L g1125 ( 
.A(n_994),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_R g1126 ( 
.A(n_992),
.B(n_1076),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_1023),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_997),
.B(n_983),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_SL g1129 ( 
.A1(n_963),
.A2(n_1029),
.B(n_1009),
.C(n_1024),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_997),
.B(n_983),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_1067),
.A2(n_989),
.B(n_1029),
.C(n_957),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_1019),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1012),
.B(n_1007),
.Y(n_1133)
);

BUFx12f_ASAP7_75t_L g1134 ( 
.A(n_1023),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1023),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1012),
.B(n_1007),
.Y(n_1136)
);

CKINVDCx11_ASAP7_75t_R g1137 ( 
.A(n_1076),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_1076),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_SL g1139 ( 
.A1(n_963),
.A2(n_1009),
.B(n_1024),
.C(n_991),
.Y(n_1139)
);

NOR2x1_ASAP7_75t_L g1140 ( 
.A(n_1021),
.B(n_1025),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1006),
.A2(n_1033),
.B(n_1015),
.Y(n_1141)
);

NOR2x1_ASAP7_75t_SL g1142 ( 
.A(n_1014),
.B(n_1021),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1032),
.A2(n_1047),
.B1(n_998),
.B2(n_996),
.Y(n_1143)
);

AO21x1_ASAP7_75t_L g1144 ( 
.A1(n_987),
.A2(n_1018),
.B(n_973),
.Y(n_1144)
);

INVx2_ASAP7_75t_SL g1145 ( 
.A(n_1028),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_1027),
.B(n_1020),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_1020),
.B(n_1013),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1020),
.B(n_1000),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1000),
.B(n_1068),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_990),
.A2(n_959),
.B(n_1081),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1000),
.B(n_1022),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1031),
.A2(n_1044),
.B(n_1073),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1005),
.B(n_1036),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1045),
.A2(n_1080),
.B(n_1062),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1054),
.A2(n_1072),
.B(n_1071),
.Y(n_1155)
);

O2A1O1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1070),
.A2(n_1011),
.B(n_976),
.C(n_1005),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1011),
.B(n_1017),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1037),
.B(n_380),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_960),
.Y(n_1159)
);

NOR2x1_ASAP7_75t_L g1160 ( 
.A(n_1065),
.B(n_868),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_972),
.A2(n_931),
.B(n_926),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_958),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_967),
.A2(n_1016),
.B(n_931),
.Y(n_1163)
);

OR2x6_ASAP7_75t_L g1164 ( 
.A(n_1042),
.B(n_736),
.Y(n_1164)
);

BUFx3_ASAP7_75t_L g1165 ( 
.A(n_1065),
.Y(n_1165)
);

OR2x6_ASAP7_75t_L g1166 ( 
.A(n_1042),
.B(n_736),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_961),
.B(n_1034),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1051),
.B(n_965),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1042),
.B(n_993),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_985),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_1065),
.Y(n_1171)
);

AND2x6_ASAP7_75t_L g1172 ( 
.A(n_1026),
.B(n_1042),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_961),
.B(n_1034),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_985),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_967),
.A2(n_931),
.B1(n_951),
.B2(n_926),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1051),
.B(n_965),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_960),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_1019),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1037),
.B(n_380),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_967),
.A2(n_1016),
.B(n_931),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1051),
.B(n_965),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1019),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_972),
.A2(n_931),
.B(n_926),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1051),
.B(n_965),
.Y(n_1184)
);

O2A1O1Ixp5_ASAP7_75t_SL g1185 ( 
.A1(n_1075),
.A2(n_659),
.B(n_1053),
.C(n_956),
.Y(n_1185)
);

BUFx12f_ASAP7_75t_L g1186 ( 
.A(n_978),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_967),
.A2(n_1016),
.B(n_931),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1065),
.Y(n_1188)
);

BUFx12f_ASAP7_75t_L g1189 ( 
.A(n_978),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_960),
.Y(n_1190)
);

BUFx3_ASAP7_75t_L g1191 ( 
.A(n_1065),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_985),
.Y(n_1192)
);

BUFx2_ASAP7_75t_SL g1193 ( 
.A(n_1065),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_967),
.A2(n_1016),
.B(n_931),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_961),
.B(n_1034),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1172),
.B(n_1089),
.Y(n_1196)
);

BUFx2_ASAP7_75t_R g1197 ( 
.A(n_1093),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1087),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_1134),
.Y(n_1199)
);

BUFx2_ASAP7_75t_SL g1200 ( 
.A(n_1094),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1113),
.B(n_1098),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1127),
.Y(n_1202)
);

INVx4_ASAP7_75t_SL g1203 ( 
.A(n_1172),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_1114),
.Y(n_1204)
);

BUFx8_ASAP7_75t_SL g1205 ( 
.A(n_1162),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1146),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_SL g1207 ( 
.A1(n_1101),
.A2(n_1182),
.B1(n_1132),
.B2(n_1178),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1159),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_1137),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1177),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1118),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1152),
.A2(n_1155),
.B(n_1154),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1146),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1110),
.Y(n_1214)
);

CKINVDCx14_ASAP7_75t_R g1215 ( 
.A(n_1107),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1172),
.A2(n_1105),
.B1(n_1128),
.B2(n_1090),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1106),
.B(n_1104),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1190),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_1149),
.B(n_1082),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1110),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1172),
.A2(n_1111),
.B1(n_1100),
.B2(n_1106),
.Y(n_1221)
);

CKINVDCx11_ASAP7_75t_R g1222 ( 
.A(n_1186),
.Y(n_1222)
);

AOI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1152),
.A2(n_1155),
.B(n_1154),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1109),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1110),
.Y(n_1225)
);

BUFx8_ASAP7_75t_SL g1226 ( 
.A(n_1189),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1132),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1178),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1182),
.Y(n_1229)
);

OA21x2_ASAP7_75t_L g1230 ( 
.A1(n_1141),
.A2(n_1121),
.B(n_1150),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1116),
.Y(n_1231)
);

BUFx2_ASAP7_75t_R g1232 ( 
.A(n_1193),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1099),
.Y(n_1233)
);

BUFx2_ASAP7_75t_R g1234 ( 
.A(n_1165),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1098),
.B(n_1082),
.Y(n_1235)
);

OR2x6_ASAP7_75t_L g1236 ( 
.A(n_1151),
.B(n_1164),
.Y(n_1236)
);

CKINVDCx6p67_ASAP7_75t_R g1237 ( 
.A(n_1191),
.Y(n_1237)
);

HB1xp67_ASAP7_75t_L g1238 ( 
.A(n_1086),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_SL g1239 ( 
.A1(n_1161),
.A2(n_1183),
.B1(n_1181),
.B2(n_1184),
.Y(n_1239)
);

INVx11_ASAP7_75t_L g1240 ( 
.A(n_1083),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1124),
.A2(n_1195),
.B1(n_1173),
.B2(n_1167),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1140),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1130),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1133),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1148),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1136),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1168),
.B(n_1176),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1171),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1136),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1188),
.B(n_1091),
.Y(n_1250)
);

CKINVDCx11_ASAP7_75t_R g1251 ( 
.A(n_1108),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1123),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1147),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1138),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_1102),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1119),
.A2(n_1168),
.B1(n_1176),
.B2(n_1181),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1119),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1115),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1125),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1143),
.B(n_1097),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1084),
.A2(n_1095),
.B1(n_1175),
.B2(n_1131),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1115),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1142),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1084),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1103),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_1164),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1125),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1135),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1135),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1131),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1112),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1163),
.A2(n_1187),
.B1(n_1180),
.B2(n_1194),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_SL g1273 ( 
.A1(n_1166),
.A2(n_1180),
.B1(n_1194),
.B2(n_1187),
.Y(n_1273)
);

BUFx2_ASAP7_75t_SL g1274 ( 
.A(n_1169),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1143),
.B(n_1163),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1096),
.B(n_1185),
.Y(n_1276)
);

AOI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1144),
.A2(n_1153),
.B(n_1157),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_1126),
.Y(n_1278)
);

OA21x2_ASAP7_75t_L g1279 ( 
.A1(n_1145),
.A2(n_1139),
.B(n_1129),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1085),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1122),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1156),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1085),
.B(n_1088),
.Y(n_1283)
);

INVx2_ASAP7_75t_SL g1284 ( 
.A(n_1117),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1120),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1088),
.A2(n_1092),
.B1(n_1170),
.B2(n_1174),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_SL g1287 ( 
.A(n_1160),
.Y(n_1287)
);

AO21x1_ASAP7_75t_L g1288 ( 
.A1(n_1170),
.A2(n_1174),
.B(n_1192),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1113),
.B(n_1098),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1172),
.B(n_1089),
.Y(n_1290)
);

INVx1_ASAP7_75t_SL g1291 ( 
.A(n_1193),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1087),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1146),
.Y(n_1293)
);

AOI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1158),
.A2(n_1179),
.B1(n_1037),
.B2(n_939),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1172),
.B(n_1089),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1087),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1227),
.B(n_1228),
.Y(n_1297)
);

AO21x2_ASAP7_75t_L g1298 ( 
.A1(n_1276),
.A2(n_1282),
.B(n_1223),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1272),
.A2(n_1261),
.A3(n_1258),
.B(n_1262),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1235),
.B(n_1201),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1235),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1206),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1231),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1201),
.B(n_1289),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1227),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1228),
.Y(n_1306)
);

NOR2x1_ASAP7_75t_SL g1307 ( 
.A(n_1217),
.B(n_1236),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1229),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1219),
.Y(n_1309)
);

BUFx4f_ASAP7_75t_SL g1310 ( 
.A(n_1278),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1219),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1247),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1247),
.Y(n_1313)
);

OR2x6_ASAP7_75t_L g1314 ( 
.A(n_1206),
.B(n_1213),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1229),
.B(n_1213),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1243),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1260),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1260),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1239),
.B(n_1257),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1289),
.B(n_1275),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1252),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1275),
.B(n_1253),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1224),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1277),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1226),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1238),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1245),
.B(n_1198),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1259),
.Y(n_1328)
);

BUFx12f_ASAP7_75t_L g1329 ( 
.A(n_1222),
.Y(n_1329)
);

CKINVDCx8_ASAP7_75t_R g1330 ( 
.A(n_1274),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1296),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1245),
.B(n_1293),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1267),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1208),
.B(n_1210),
.Y(n_1334)
);

AO21x2_ASAP7_75t_L g1335 ( 
.A1(n_1276),
.A2(n_1223),
.B(n_1270),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1218),
.B(n_1292),
.Y(n_1336)
);

CKINVDCx8_ASAP7_75t_R g1337 ( 
.A(n_1200),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1233),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1293),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1293),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1211),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1244),
.Y(n_1342)
);

CKINVDCx20_ASAP7_75t_R g1343 ( 
.A(n_1205),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1246),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1230),
.Y(n_1345)
);

OA21x2_ASAP7_75t_L g1346 ( 
.A1(n_1212),
.A2(n_1256),
.B(n_1264),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1249),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1230),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1273),
.B(n_1241),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1279),
.A2(n_1288),
.B(n_1263),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1279),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1203),
.B(n_1196),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1207),
.B(n_1216),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_1205),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1242),
.Y(n_1355)
);

AOI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1280),
.A2(n_1285),
.B(n_1271),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1196),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1280),
.B(n_1221),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1284),
.B(n_1269),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1268),
.Y(n_1360)
);

AO21x2_ASAP7_75t_L g1361 ( 
.A1(n_1265),
.A2(n_1281),
.B(n_1294),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_1234),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_1202),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1331),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1310),
.B(n_1237),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1297),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1300),
.B(n_1250),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1305),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1331),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1320),
.B(n_1304),
.Y(n_1370)
);

INVxp67_ASAP7_75t_L g1371 ( 
.A(n_1361),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_1297),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1301),
.B(n_1254),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1320),
.B(n_1304),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1301),
.B(n_1291),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1317),
.B(n_1202),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_1302),
.Y(n_1377)
);

INVx4_ASAP7_75t_L g1378 ( 
.A(n_1314),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1318),
.B(n_1220),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1318),
.B(n_1220),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1309),
.B(n_1283),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1306),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1306),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1312),
.B(n_1313),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1312),
.B(n_1313),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1308),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1298),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1315),
.B(n_1209),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1322),
.B(n_1225),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1322),
.B(n_1220),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1315),
.B(n_1209),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1303),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1327),
.B(n_1214),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1357),
.B(n_1203),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1327),
.B(n_1214),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1298),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1311),
.B(n_1204),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1343),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1298),
.Y(n_1399)
);

INVx4_ASAP7_75t_L g1400 ( 
.A(n_1314),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1342),
.B(n_1286),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1314),
.B(n_1237),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_SL g1403 ( 
.A1(n_1349),
.A2(n_1196),
.B(n_1290),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1314),
.B(n_1204),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1314),
.B(n_1295),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1299),
.B(n_1248),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1335),
.Y(n_1407)
);

OAI21xp5_ASAP7_75t_SL g1408 ( 
.A1(n_1406),
.A2(n_1353),
.B(n_1319),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1370),
.B(n_1341),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1370),
.B(n_1326),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1374),
.B(n_1321),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1392),
.B(n_1344),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1367),
.B(n_1347),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1367),
.B(n_1355),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1368),
.B(n_1338),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1403),
.A2(n_1330),
.B1(n_1337),
.B2(n_1358),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1384),
.B(n_1351),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1368),
.B(n_1323),
.Y(n_1418)
);

OAI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1401),
.A2(n_1356),
.B(n_1350),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1366),
.B(n_1316),
.Y(n_1420)
);

OAI221xp5_ASAP7_75t_SL g1421 ( 
.A1(n_1403),
.A2(n_1358),
.B1(n_1351),
.B2(n_1332),
.C(n_1362),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1366),
.B(n_1361),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1384),
.B(n_1335),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_SL g1424 ( 
.A(n_1398),
.B(n_1329),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1401),
.B(n_1363),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1397),
.A2(n_1337),
.B1(n_1363),
.B2(n_1248),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1402),
.A2(n_1215),
.B(n_1329),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1385),
.B(n_1335),
.Y(n_1428)
);

OA21x2_ASAP7_75t_L g1429 ( 
.A1(n_1371),
.A2(n_1350),
.B(n_1348),
.Y(n_1429)
);

NAND3xp33_ASAP7_75t_L g1430 ( 
.A(n_1387),
.B(n_1399),
.C(n_1396),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1372),
.B(n_1328),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1385),
.B(n_1346),
.Y(n_1432)
);

NAND3xp33_ASAP7_75t_L g1433 ( 
.A(n_1407),
.B(n_1333),
.C(n_1360),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1376),
.B(n_1389),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1376),
.B(n_1346),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_SL g1436 ( 
.A1(n_1404),
.A2(n_1329),
.B1(n_1266),
.B2(n_1354),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1389),
.B(n_1346),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1397),
.A2(n_1332),
.B1(n_1232),
.B2(n_1240),
.Y(n_1438)
);

NAND3xp33_ASAP7_75t_L g1439 ( 
.A(n_1387),
.B(n_1340),
.C(n_1339),
.Y(n_1439)
);

AOI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1396),
.A2(n_1356),
.B(n_1345),
.Y(n_1440)
);

NAND4xp25_ASAP7_75t_L g1441 ( 
.A(n_1388),
.B(n_1334),
.C(n_1336),
.D(n_1359),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_SL g1442 ( 
.A1(n_1394),
.A2(n_1307),
.B(n_1352),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1372),
.B(n_1373),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1404),
.B(n_1394),
.Y(n_1444)
);

NAND3xp33_ASAP7_75t_L g1445 ( 
.A(n_1399),
.B(n_1339),
.C(n_1340),
.Y(n_1445)
);

NOR2x1_ASAP7_75t_L g1446 ( 
.A(n_1378),
.B(n_1324),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1390),
.B(n_1299),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1373),
.B(n_1336),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1383),
.B(n_1299),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1382),
.B(n_1386),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1390),
.B(n_1393),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1365),
.B(n_1251),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1388),
.B(n_1251),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1393),
.B(n_1299),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1382),
.B(n_1299),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1391),
.A2(n_1240),
.B1(n_1255),
.B2(n_1287),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1395),
.B(n_1299),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1364),
.Y(n_1458)
);

AND2x2_ASAP7_75t_SL g1459 ( 
.A(n_1378),
.B(n_1352),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1454),
.B(n_1378),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1458),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1440),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1440),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1429),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1443),
.B(n_1375),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1458),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1450),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1449),
.B(n_1375),
.Y(n_1468)
);

NAND2x1_ASAP7_75t_L g1469 ( 
.A(n_1442),
.B(n_1400),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1423),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1428),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1424),
.B(n_1215),
.Y(n_1472)
);

INVxp67_ASAP7_75t_SL g1473 ( 
.A(n_1455),
.Y(n_1473)
);

INVxp67_ASAP7_75t_SL g1474 ( 
.A(n_1422),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1429),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1418),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1433),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1433),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1452),
.B(n_1325),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1457),
.B(n_1379),
.Y(n_1480)
);

INVx4_ASAP7_75t_L g1481 ( 
.A(n_1459),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1457),
.B(n_1379),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1432),
.B(n_1380),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1415),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1447),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1459),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1432),
.B(n_1364),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1447),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1439),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1437),
.B(n_1369),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1451),
.B(n_1417),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1448),
.B(n_1381),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1451),
.B(n_1400),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1445),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1430),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1435),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1420),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1413),
.B(n_1410),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1435),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1437),
.B(n_1380),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1461),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1461),
.Y(n_1502)
);

NAND2xp33_ASAP7_75t_L g1503 ( 
.A(n_1486),
.B(n_1436),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1468),
.B(n_1431),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1466),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1480),
.B(n_1434),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1481),
.Y(n_1507)
);

OAI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1489),
.A2(n_1408),
.B(n_1419),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1489),
.B(n_1412),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1464),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1466),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1494),
.B(n_1409),
.Y(n_1512)
);

NOR2x1_ASAP7_75t_L g1513 ( 
.A(n_1472),
.B(n_1427),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1497),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1497),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1476),
.Y(n_1516)
);

BUFx2_ASAP7_75t_L g1517 ( 
.A(n_1481),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1480),
.B(n_1459),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1476),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_1494),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1484),
.B(n_1414),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1464),
.Y(n_1522)
);

INVx2_ASAP7_75t_SL g1523 ( 
.A(n_1493),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1465),
.Y(n_1524)
);

INVxp67_ASAP7_75t_L g1525 ( 
.A(n_1495),
.Y(n_1525)
);

NAND2x1p5_ASAP7_75t_L g1526 ( 
.A(n_1469),
.B(n_1446),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1481),
.B(n_1402),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1468),
.B(n_1411),
.Y(n_1528)
);

NAND2x1_ASAP7_75t_L g1529 ( 
.A(n_1481),
.B(n_1442),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1480),
.B(n_1453),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1490),
.B(n_1441),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1465),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1464),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1486),
.B(n_1444),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1492),
.Y(n_1535)
);

AND2x4_ASAP7_75t_L g1536 ( 
.A(n_1486),
.B(n_1405),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1492),
.Y(n_1537)
);

CKINVDCx16_ASAP7_75t_R g1538 ( 
.A(n_1479),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1490),
.B(n_1421),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1484),
.B(n_1425),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1482),
.B(n_1377),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1475),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1518),
.B(n_1506),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_SL g1544 ( 
.A(n_1538),
.B(n_1486),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1501),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1520),
.B(n_1477),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1502),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1510),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1525),
.B(n_1477),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1518),
.B(n_1496),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1505),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1512),
.B(n_1478),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1508),
.A2(n_1478),
.B(n_1495),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1535),
.B(n_1487),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1511),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1517),
.B(n_1496),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1514),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1506),
.B(n_1482),
.Y(n_1558)
);

AOI221xp5_ASAP7_75t_L g1559 ( 
.A1(n_1539),
.A2(n_1473),
.B1(n_1470),
.B2(n_1474),
.C(n_1488),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1537),
.B(n_1487),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1510),
.Y(n_1561)
);

BUFx2_ASAP7_75t_L g1562 ( 
.A(n_1513),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1509),
.B(n_1467),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1517),
.B(n_1482),
.Y(n_1564)
);

NAND2x1p5_ASAP7_75t_L g1565 ( 
.A(n_1529),
.B(n_1469),
.Y(n_1565)
);

NOR3xp33_ASAP7_75t_L g1566 ( 
.A(n_1503),
.B(n_1463),
.C(n_1462),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1523),
.B(n_1491),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1524),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1532),
.B(n_1531),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1521),
.B(n_1467),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1523),
.B(n_1534),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1522),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1534),
.B(n_1491),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1516),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1519),
.B(n_1473),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1515),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1528),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1528),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1530),
.B(n_1222),
.Y(n_1579)
);

NOR4xp25_ASAP7_75t_L g1580 ( 
.A(n_1503),
.B(n_1539),
.C(n_1540),
.D(n_1531),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1534),
.B(n_1499),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1504),
.B(n_1485),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1536),
.B(n_1499),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1504),
.B(n_1485),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1522),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1530),
.B(n_1470),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1507),
.B(n_1488),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1545),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1545),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1562),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1547),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1543),
.B(n_1527),
.Y(n_1592)
);

OAI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1562),
.A2(n_1529),
.B1(n_1527),
.B2(n_1507),
.Y(n_1593)
);

CKINVDCx16_ASAP7_75t_R g1594 ( 
.A(n_1580),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1547),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1553),
.A2(n_1527),
.B1(n_1507),
.B2(n_1526),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1551),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1543),
.B(n_1536),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1573),
.B(n_1536),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1579),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1576),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1566),
.A2(n_1526),
.B1(n_1436),
.B2(n_1416),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1577),
.B(n_1483),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1551),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1573),
.B(n_1541),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1565),
.Y(n_1606)
);

OR2x6_ASAP7_75t_L g1607 ( 
.A(n_1565),
.B(n_1533),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1571),
.B(n_1460),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1558),
.B(n_1541),
.Y(n_1609)
);

NOR2x1_ASAP7_75t_L g1610 ( 
.A(n_1546),
.B(n_1456),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1558),
.B(n_1493),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1567),
.B(n_1500),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1578),
.B(n_1483),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1555),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1564),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1557),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1557),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1569),
.B(n_1498),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1567),
.B(n_1500),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1549),
.B(n_1483),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1564),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1581),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1552),
.B(n_1471),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1574),
.Y(n_1624)
);

OAI22xp33_ASAP7_75t_SL g1625 ( 
.A1(n_1594),
.A2(n_1569),
.B1(n_1565),
.B2(n_1544),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1588),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1594),
.Y(n_1627)
);

OAI21xp33_ASAP7_75t_L g1628 ( 
.A1(n_1610),
.A2(n_1559),
.B(n_1571),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1602),
.A2(n_1561),
.B1(n_1572),
.B2(n_1548),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1588),
.Y(n_1630)
);

OAI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1618),
.A2(n_1586),
.B1(n_1550),
.B2(n_1563),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1589),
.Y(n_1632)
);

A2O1A1Ixp33_ASAP7_75t_L g1633 ( 
.A1(n_1600),
.A2(n_1590),
.B(n_1596),
.C(n_1618),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1592),
.B(n_1550),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1589),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1591),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1601),
.B(n_1568),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_1622),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1591),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1595),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1615),
.B(n_1570),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1615),
.B(n_1554),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1622),
.Y(n_1643)
);

XOR2x2_ASAP7_75t_L g1644 ( 
.A(n_1606),
.B(n_1438),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1595),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1621),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1597),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1592),
.B(n_1226),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1621),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1597),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1604),
.Y(n_1651)
);

INVx3_ASAP7_75t_L g1652 ( 
.A(n_1627),
.Y(n_1652)
);

OAI21xp33_ASAP7_75t_L g1653 ( 
.A1(n_1628),
.A2(n_1598),
.B(n_1620),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1634),
.B(n_1599),
.Y(n_1654)
);

NAND3xp33_ASAP7_75t_L g1655 ( 
.A(n_1633),
.B(n_1624),
.C(n_1614),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1646),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1646),
.Y(n_1657)
);

NOR2x1_ASAP7_75t_L g1658 ( 
.A(n_1648),
.B(n_1606),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1649),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1638),
.Y(n_1660)
);

AND2x4_ASAP7_75t_SL g1661 ( 
.A(n_1648),
.B(n_1608),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1638),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1649),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1626),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1643),
.B(n_1612),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1642),
.B(n_1599),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_1637),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1630),
.Y(n_1668)
);

NAND2xp33_ASAP7_75t_L g1669 ( 
.A(n_1633),
.B(n_1593),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1644),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1644),
.Y(n_1671)
);

OAI211xp5_ASAP7_75t_L g1672 ( 
.A1(n_1652),
.A2(n_1629),
.B(n_1635),
.C(n_1632),
.Y(n_1672)
);

NOR3xp33_ASAP7_75t_L g1673 ( 
.A(n_1652),
.B(n_1625),
.C(n_1641),
.Y(n_1673)
);

OAI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1671),
.A2(n_1669),
.B1(n_1652),
.B2(n_1629),
.C(n_1670),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_SL g1675 ( 
.A(n_1658),
.B(n_1197),
.Y(n_1675)
);

OAI221xp5_ASAP7_75t_SL g1676 ( 
.A1(n_1653),
.A2(n_1607),
.B1(n_1650),
.B2(n_1647),
.C(n_1645),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_SL g1677 ( 
.A(n_1670),
.B(n_1556),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1669),
.A2(n_1631),
.B1(n_1607),
.B2(n_1585),
.Y(n_1678)
);

O2A1O1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1655),
.A2(n_1636),
.B(n_1640),
.C(n_1639),
.Y(n_1679)
);

AOI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1663),
.A2(n_1607),
.B1(n_1585),
.B2(n_1561),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1666),
.B(n_1612),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1665),
.B(n_1603),
.Y(n_1682)
);

NOR3x1_ASAP7_75t_L g1683 ( 
.A(n_1664),
.B(n_1651),
.C(n_1624),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1677),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1681),
.B(n_1654),
.Y(n_1685)
);

NOR4xp25_ASAP7_75t_L g1686 ( 
.A(n_1674),
.B(n_1662),
.C(n_1667),
.D(n_1657),
.Y(n_1686)
);

NAND3xp33_ASAP7_75t_L g1687 ( 
.A(n_1673),
.B(n_1660),
.C(n_1662),
.Y(n_1687)
);

NOR3xp33_ASAP7_75t_L g1688 ( 
.A(n_1672),
.B(n_1663),
.C(n_1657),
.Y(n_1688)
);

NAND3xp33_ASAP7_75t_L g1689 ( 
.A(n_1678),
.B(n_1659),
.C(n_1656),
.Y(n_1689)
);

NAND2x1_ASAP7_75t_L g1690 ( 
.A(n_1680),
.B(n_1666),
.Y(n_1690)
);

OAI322xp33_ASAP7_75t_L g1691 ( 
.A1(n_1679),
.A2(n_1656),
.A3(n_1659),
.B1(n_1668),
.B2(n_1604),
.C1(n_1616),
.C2(n_1617),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1683),
.B(n_1654),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1682),
.Y(n_1693)
);

NAND3xp33_ASAP7_75t_L g1694 ( 
.A(n_1676),
.B(n_1617),
.C(n_1616),
.Y(n_1694)
);

NAND4xp25_ASAP7_75t_L g1695 ( 
.A(n_1687),
.B(n_1675),
.C(n_1598),
.D(n_1614),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1685),
.Y(n_1696)
);

NOR2xp67_ASAP7_75t_L g1697 ( 
.A(n_1684),
.B(n_1608),
.Y(n_1697)
);

NAND3xp33_ASAP7_75t_L g1698 ( 
.A(n_1688),
.B(n_1607),
.C(n_1556),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1693),
.B(n_1686),
.Y(n_1699)
);

OA211x2_ASAP7_75t_L g1700 ( 
.A1(n_1690),
.A2(n_1661),
.B(n_1623),
.C(n_1613),
.Y(n_1700)
);

NAND3xp33_ASAP7_75t_L g1701 ( 
.A(n_1689),
.B(n_1607),
.C(n_1556),
.Y(n_1701)
);

NAND4xp25_ASAP7_75t_SL g1702 ( 
.A(n_1692),
.B(n_1661),
.C(n_1581),
.D(n_1605),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1696),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1697),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1699),
.A2(n_1694),
.B1(n_1608),
.B2(n_1572),
.Y(n_1705)
);

AOI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1695),
.A2(n_1608),
.B1(n_1548),
.B2(n_1605),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1700),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1701),
.B(n_1619),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1698),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1702),
.Y(n_1710)
);

NAND3xp33_ASAP7_75t_SL g1711 ( 
.A(n_1704),
.B(n_1705),
.C(n_1707),
.Y(n_1711)
);

XOR2x1_ASAP7_75t_L g1712 ( 
.A(n_1703),
.B(n_1691),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1706),
.B(n_1619),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1708),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1709),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1710),
.B(n_1609),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1715),
.B(n_1609),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_SL g1718 ( 
.A1(n_1711),
.A2(n_1199),
.B(n_1287),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1712),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1716),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1719),
.B(n_1714),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1721),
.A2(n_1720),
.B1(n_1713),
.B2(n_1717),
.Y(n_1722)
);

AO22x2_ASAP7_75t_L g1723 ( 
.A1(n_1722),
.A2(n_1717),
.B1(n_1718),
.B2(n_1587),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1722),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1724),
.A2(n_1554),
.B1(n_1560),
.B2(n_1575),
.Y(n_1725)
);

INVxp33_ASAP7_75t_L g1726 ( 
.A(n_1723),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1726),
.A2(n_1560),
.B1(n_1587),
.B2(n_1583),
.Y(n_1727)
);

NAND2xp33_ASAP7_75t_SL g1728 ( 
.A(n_1725),
.B(n_1611),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1728),
.A2(n_1199),
.B(n_1583),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1729),
.A2(n_1727),
.B1(n_1611),
.B2(n_1533),
.Y(n_1730)
);

OAI221xp5_ASAP7_75t_L g1731 ( 
.A1(n_1730),
.A2(n_1584),
.B1(n_1582),
.B2(n_1426),
.C(n_1542),
.Y(n_1731)
);

AOI211xp5_ASAP7_75t_L g1732 ( 
.A1(n_1731),
.A2(n_1584),
.B(n_1582),
.C(n_1542),
.Y(n_1732)
);


endmodule