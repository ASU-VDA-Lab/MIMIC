module real_jpeg_32748_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g289 ( 
.A(n_0),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_1),
.B(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_1),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_1),
.B(n_169),
.Y(n_266)
);

OAI32xp33_ASAP7_75t_L g300 ( 
.A1(n_1),
.A2(n_301),
.A3(n_304),
.B1(n_309),
.B2(n_315),
.Y(n_300)
);

OAI21xp33_ASAP7_75t_L g380 ( 
.A1(n_1),
.A2(n_174),
.B(n_381),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_1),
.A2(n_244),
.B1(n_434),
.B2(n_438),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_2),
.A2(n_186),
.B1(n_191),
.B2(n_192),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_2),
.Y(n_191)
);

AO22x1_ASAP7_75t_L g269 ( 
.A1(n_2),
.A2(n_191),
.B1(n_270),
.B2(n_273),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_3),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_3),
.Y(n_149)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_4),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_4),
.Y(n_111)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_5),
.Y(n_199)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_5),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_6),
.A2(n_177),
.B1(n_180),
.B2(n_183),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_6),
.Y(n_183)
);

OAI22x1_ASAP7_75t_L g59 ( 
.A1(n_7),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_59)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_7),
.A2(n_65),
.B1(n_221),
.B2(n_225),
.Y(n_220)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_8),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_8),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_8),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_8),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_10),
.A2(n_125),
.B1(n_128),
.B2(n_129),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_10),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_10),
.A2(n_128),
.B1(n_135),
.B2(n_139),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_10),
.A2(n_128),
.B1(n_232),
.B2(n_234),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_10),
.A2(n_128),
.B1(n_293),
.B2(n_298),
.Y(n_292)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_11),
.Y(n_202)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_11),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_11),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_12),
.A2(n_87),
.B1(n_91),
.B2(n_92),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_12),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_12),
.A2(n_91),
.B1(n_322),
.B2(n_324),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g342 ( 
.A1(n_12),
.A2(n_91),
.B1(n_343),
.B2(n_346),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_13),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_14),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_14),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_15),
.A2(n_163),
.B1(n_164),
.B2(n_166),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_15),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_15),
.A2(n_163),
.B1(n_248),
.B2(n_251),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_15),
.A2(n_163),
.B1(n_336),
.B2(n_338),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_15),
.A2(n_163),
.B1(n_409),
.B2(n_412),
.Y(n_408)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_278),
.B1(n_453),
.B2(n_454),
.Y(n_17)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_18),
.Y(n_454)
);

NAND2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_276),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_257),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_21),
.B(n_257),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_171),
.Y(n_21)
);

XNOR2x1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_83),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_51),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_24),
.B(n_51),
.Y(n_260)
);

AOI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.A3(n_34),
.B1(n_39),
.B2(n_43),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_29),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_29),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_29),
.Y(n_437)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_32),
.Y(n_145)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_33),
.Y(n_158)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g165 ( 
.A(n_37),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_38),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_38),
.Y(n_144)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_39),
.Y(n_245)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp33_ASAP7_75t_R g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_45),
.Y(n_160)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_50),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_59),
.B1(n_71),
.B2(n_75),
.Y(n_51)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_52),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_52),
.B(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_52),
.A2(n_275),
.B1(n_334),
.B2(n_341),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_53),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_173)
);

INVx3_ASAP7_75t_SL g275 ( 
.A(n_53),
.Y(n_275)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_55),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_55),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_55),
.Y(n_426)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_58),
.Y(n_179)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_58),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_58),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_59),
.B(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_69),
.Y(n_204)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_70),
.Y(n_367)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_74),
.Y(n_392)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_75),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g340 ( 
.A(n_82),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_132),
.B2(n_170),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_97),
.B(n_122),
.Y(n_85)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_86),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_90),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OA21x2_ASAP7_75t_L g432 ( 
.A1(n_97),
.A2(n_122),
.B(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22x1_ASAP7_75t_L g246 ( 
.A1(n_98),
.A2(n_247),
.B1(n_252),
.B2(n_253),
.Y(n_246)
);

NAND2xp33_ASAP7_75t_SL g265 ( 
.A(n_98),
.B(n_124),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_112),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_104),
.B1(n_107),
.B2(n_109),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_101),
.Y(n_318)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_102),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_108),
.Y(n_323)
);

INVx5_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_115),
.B1(n_118),
.B2(n_121),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_114),
.Y(n_250)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_114),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_117),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_123),
.Y(n_254)
);

INVxp67_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_161),
.Y(n_132)
);

NAND2x1_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_141),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_134),
.B(n_169),
.Y(n_240)
);

INVx3_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_139),
.Y(n_243)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_141),
.B(n_242),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_153),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_145),
.B1(n_146),
.B2(n_150),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

AOI22x1_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_169),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_228),
.B1(n_255),
.B2(n_256),
.Y(n_171)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_172),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_184),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_174),
.A2(n_269),
.B(n_274),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_174),
.A2(n_342),
.B(n_381),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_177),
.B(n_388),
.Y(n_387)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_182),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_195),
.B1(n_220),
.B2(n_227),
.Y(n_184)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_185),
.Y(n_237)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx4f_ASAP7_75t_SL g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_190),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_190),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_194),
.Y(n_236)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_195),
.A2(n_321),
.B(n_325),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_207),
.Y(n_195)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

OAI22x1_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_200),
.B1(n_203),
.B2(n_205),
.Y(n_196)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_197),
.Y(n_345)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_199),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_199),
.Y(n_337)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_202),
.Y(n_206)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_210),
.B1(n_214),
.B2(n_217),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx6_ASAP7_75t_L g362 ( 
.A(n_212),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_219),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_219),
.Y(n_411)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_224),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_226),
.Y(n_233)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_227),
.Y(n_430)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_228),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_239),
.C(n_246),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_246),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_237),
.B2(n_238),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_230),
.B(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_230),
.B(n_231),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_230),
.A2(n_429),
.B1(n_430),
.B2(n_431),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_231),
.B(n_238),
.Y(n_325)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_236),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_238),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B(n_245),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_244),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_244),
.B(n_307),
.Y(n_354)
);

OAI21xp33_ASAP7_75t_L g373 ( 
.A1(n_244),
.A2(n_354),
.B(n_374),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_244),
.B(n_389),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_244),
.B(n_395),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_244),
.B(n_254),
.Y(n_406)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_254),
.A2(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.C(n_261),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_266),
.C(n_267),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_263),
.B(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_266),
.B(n_268),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_R g286 ( 
.A(n_269),
.B(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_269),
.A2(n_291),
.B(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_272),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_278),
.Y(n_453)
);

OAI21x1_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_329),
.B(n_451),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_280),
.Y(n_452)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_284),
.B(n_452),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_319),
.C(n_326),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_285),
.A2(n_319),
.B1(n_320),
.B2(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_285),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_290),
.B(n_300),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx8_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVxp67_ASAP7_75t_SL g290 ( 
.A(n_291),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_SL g396 ( 
.A1(n_291),
.A2(n_335),
.B(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_292),
.B(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_297),
.Y(n_350)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_300),
.B(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_303),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_321),
.Y(n_431)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_325),
.B(n_372),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_327),
.B(n_445),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_442),
.B(n_450),
.Y(n_329)
);

O2A1O1Ixp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_401),
.B(n_417),
.C(n_418),
.Y(n_330)
);

AOI21x1_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_378),
.B(n_400),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_351),
.Y(n_332)
);

NOR2xp67_ASAP7_75t_L g400 ( 
.A(n_333),
.B(n_351),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVxp33_ASAP7_75t_SL g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_371),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_352),
.B(n_371),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_355),
.B1(n_363),
.B2(n_368),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_358),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_358),
.B(n_369),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

OAI21xp33_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_393),
.B(n_399),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_387),
.Y(n_379)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_392),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_396),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_394),
.B(n_396),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_395),
.A2(n_408),
.B(n_416),
.Y(n_407)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

NOR2xp67_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_402),
.B(n_403),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_404),
.B(n_420),
.C(n_421),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_406),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_407),
.Y(n_420)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_408),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_410),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_413),
.Y(n_412)
);

INVx4_ASAP7_75t_SL g413 ( 
.A(n_414),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_422),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_419),
.B(n_422),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_427),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_423),
.Y(n_448)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_432),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_432),
.C(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_443),
.B(n_449),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_447),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g450 ( 
.A(n_444),
.B(n_447),
.Y(n_450)
);


endmodule