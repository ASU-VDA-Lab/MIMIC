module fake_aes_3057_n_681 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_681);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_681;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_529;
wire n_312;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_466;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_SL g77 ( .A(n_17), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_54), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_3), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_39), .Y(n_80) );
INVx3_ASAP7_75t_L g81 ( .A(n_29), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_18), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_61), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_40), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_16), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_71), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_2), .Y(n_87) );
CKINVDCx20_ASAP7_75t_R g88 ( .A(n_9), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_66), .Y(n_89) );
INVxp33_ASAP7_75t_SL g90 ( .A(n_58), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_47), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_2), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_5), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_37), .Y(n_94) );
BUFx3_ASAP7_75t_L g95 ( .A(n_36), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_14), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_10), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_64), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_60), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_4), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_3), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_31), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_19), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_11), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_49), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_30), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_73), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_9), .Y(n_108) );
BUFx3_ASAP7_75t_L g109 ( .A(n_21), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_45), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_52), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_15), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_8), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_4), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_67), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_10), .B(n_76), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_62), .Y(n_117) );
INVxp33_ASAP7_75t_SL g118 ( .A(n_22), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_74), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_24), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_57), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_33), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_13), .Y(n_123) );
AND2x4_ASAP7_75t_L g124 ( .A(n_81), .B(n_0), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_104), .B(n_0), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_81), .Y(n_126) );
INVx4_ASAP7_75t_L g127 ( .A(n_81), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_123), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_80), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_83), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_92), .B(n_1), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_90), .A2(n_1), .B1(n_5), .B2(n_6), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_92), .B(n_6), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_93), .B(n_7), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_95), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_80), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_117), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_95), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_78), .B(n_7), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_117), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_85), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_85), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_99), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_86), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_79), .B(n_8), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_101), .B(n_11), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_93), .B(n_12), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_86), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_113), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_108), .B(n_12), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_91), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_91), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_115), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_109), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_98), .B(n_13), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_115), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_113), .B(n_14), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_119), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_114), .B(n_20), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_119), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_120), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_120), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_109), .Y(n_164) );
CKINVDCx16_ASAP7_75t_R g165 ( .A(n_88), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_121), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_144), .B(n_99), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_144), .B(n_105), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_127), .B(n_105), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_135), .Y(n_170) );
NOR3xp33_ASAP7_75t_L g171 ( .A(n_146), .B(n_87), .C(n_97), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_127), .B(n_118), .Y(n_172) );
NAND3xp33_ASAP7_75t_L g173 ( .A(n_125), .B(n_123), .C(n_114), .Y(n_173) );
INVx2_ASAP7_75t_SL g174 ( .A(n_127), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_124), .B(n_90), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_130), .B(n_118), .Y(n_176) );
BUFx8_ASAP7_75t_L g177 ( .A(n_125), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_130), .B(n_102), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_124), .B(n_106), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_138), .B(n_110), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_128), .B(n_96), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_135), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_124), .B(n_100), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_135), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_135), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_134), .Y(n_186) );
INVxp67_ASAP7_75t_L g187 ( .A(n_160), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_138), .B(n_111), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_142), .B(n_121), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_135), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_142), .B(n_122), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_134), .Y(n_192) );
INVxp67_ASAP7_75t_L g193 ( .A(n_160), .Y(n_193) );
BUFx6f_ASAP7_75t_SL g194 ( .A(n_134), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_147), .A2(n_94), .B(n_82), .C(n_107), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_131), .A2(n_112), .B1(n_89), .B2(n_84), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g197 ( .A1(n_132), .A2(n_103), .B1(n_77), .B2(n_116), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_150), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_139), .Y(n_199) );
OAI221xp5_ASAP7_75t_L g200 ( .A1(n_149), .A2(n_23), .B1(n_25), .B2(n_26), .C(n_27), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_139), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_150), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_150), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_149), .B(n_28), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_126), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_126), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_131), .Y(n_207) );
NOR3xp33_ASAP7_75t_L g208 ( .A(n_151), .B(n_32), .C(n_34), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_152), .B(n_35), .Y(n_209) );
INVxp67_ASAP7_75t_L g210 ( .A(n_133), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_133), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_152), .B(n_38), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_148), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_148), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_153), .B(n_41), .Y(n_215) );
BUFx5_ASAP7_75t_L g216 ( .A(n_153), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_154), .B(n_42), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_154), .B(n_43), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_163), .B(n_44), .Y(n_219) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_158), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_163), .B(n_46), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_143), .B(n_48), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_143), .B(n_50), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_198), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_220), .B(n_158), .Y(n_225) );
INVx2_ASAP7_75t_SL g226 ( .A(n_220), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_210), .B(n_165), .Y(n_227) );
BUFx3_ASAP7_75t_L g228 ( .A(n_184), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_210), .B(n_162), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_216), .Y(n_230) );
BUFx3_ASAP7_75t_L g231 ( .A(n_185), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_202), .Y(n_232) );
INVx2_ASAP7_75t_SL g233 ( .A(n_186), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_182), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_203), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_205), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_187), .B(n_156), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_216), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_216), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_206), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_216), .Y(n_241) );
INVx3_ASAP7_75t_L g242 ( .A(n_194), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_187), .B(n_145), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_216), .B(n_166), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_192), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_193), .B(n_145), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_193), .B(n_157), .Y(n_247) );
INVx2_ASAP7_75t_SL g248 ( .A(n_216), .Y(n_248) );
AND2x4_ASAP7_75t_L g249 ( .A(n_207), .B(n_157), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_211), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_213), .B(n_162), .Y(n_251) );
AND2x6_ASAP7_75t_L g252 ( .A(n_214), .B(n_161), .Y(n_252) );
INVx2_ASAP7_75t_SL g253 ( .A(n_181), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_176), .B(n_140), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_170), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_189), .Y(n_256) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_177), .Y(n_257) );
NAND2x1_ASAP7_75t_L g258 ( .A(n_174), .B(n_159), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_173), .B(n_159), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_191), .B(n_161), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_179), .Y(n_261) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_177), .Y(n_262) );
AND3x1_ASAP7_75t_SL g263 ( .A(n_200), .B(n_166), .C(n_141), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_172), .B(n_129), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_175), .B(n_129), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_169), .Y(n_266) );
BUFx3_ASAP7_75t_L g267 ( .A(n_182), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_178), .B(n_141), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_196), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_180), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_204), .B(n_166), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_195), .A2(n_137), .B(n_136), .C(n_166), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_171), .A2(n_166), .B1(n_164), .B2(n_155), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_190), .Y(n_274) );
INVxp67_ASAP7_75t_L g275 ( .A(n_183), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_221), .B(n_164), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_188), .B(n_137), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_195), .B(n_136), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_171), .B(n_164), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_167), .B(n_164), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_168), .B(n_164), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_194), .A2(n_155), .B1(n_139), .B2(n_55), .Y(n_282) );
AOI22x1_ASAP7_75t_L g283 ( .A1(n_199), .A2(n_155), .B1(n_139), .B2(n_56), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_223), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_209), .B(n_155), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_223), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_270), .B(n_197), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_226), .A2(n_208), .B1(n_219), .B2(n_217), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_256), .B(n_208), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_230), .Y(n_290) );
A2O1A1Ixp33_ASAP7_75t_L g291 ( .A1(n_254), .A2(n_215), .B(n_222), .C(n_218), .Y(n_291) );
CKINVDCx6p67_ASAP7_75t_R g292 ( .A(n_257), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_226), .B(n_155), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g294 ( .A1(n_233), .A2(n_212), .B1(n_139), .B2(n_201), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_246), .B(n_237), .Y(n_295) );
INVx1_ASAP7_75t_SL g296 ( .A(n_225), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_227), .B(n_182), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_262), .Y(n_298) );
NAND3xp33_ASAP7_75t_L g299 ( .A(n_272), .B(n_182), .C(n_53), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_230), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_246), .B(n_75), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_238), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_229), .B(n_51), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_224), .Y(n_304) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_284), .A2(n_59), .B(n_63), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_271), .A2(n_65), .B(n_68), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_232), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_235), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_242), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_260), .B(n_69), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_252), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_238), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_239), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_254), .B(n_70), .Y(n_314) );
INVx1_ASAP7_75t_SL g315 ( .A(n_252), .Y(n_315) );
NOR2xp67_ASAP7_75t_L g316 ( .A(n_233), .B(n_72), .Y(n_316) );
NOR2xp67_ASAP7_75t_L g317 ( .A(n_275), .B(n_242), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_236), .Y(n_318) );
A2O1A1Ixp33_ASAP7_75t_SL g319 ( .A1(n_265), .A2(n_273), .B(n_286), .C(n_242), .Y(n_319) );
NOR2x1_ASAP7_75t_SL g320 ( .A(n_248), .B(n_266), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_252), .Y(n_321) );
INVx2_ASAP7_75t_SL g322 ( .A(n_252), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_249), .B(n_251), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_253), .B(n_247), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_228), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_249), .B(n_251), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_250), .A2(n_245), .B1(n_243), .B2(n_253), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_252), .Y(n_328) );
INVx4_ASAP7_75t_L g329 ( .A(n_252), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_228), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_249), .B(n_251), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_264), .A2(n_265), .B1(n_279), .B2(n_259), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_240), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_268), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_239), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_261), .B(n_259), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_241), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_290), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_334), .B(n_259), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_334), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_296), .Y(n_341) );
INVx3_ASAP7_75t_L g342 ( .A(n_329), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_304), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_304), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_329), .Y(n_345) );
OAI21x1_ASAP7_75t_L g346 ( .A1(n_305), .A2(n_276), .B(n_271), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_290), .Y(n_347) );
NOR2xp33_ASAP7_75t_SL g348 ( .A(n_292), .B(n_269), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_295), .B(n_277), .Y(n_349) );
HB1xp67_ASAP7_75t_SL g350 ( .A(n_298), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_300), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_329), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_324), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_307), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_307), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_308), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_324), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_308), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_318), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_318), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_298), .B(n_269), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_333), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_333), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_289), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_331), .Y(n_365) );
BUFx2_ASAP7_75t_R g366 ( .A(n_309), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_300), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_323), .Y(n_368) );
BUFx3_ASAP7_75t_L g369 ( .A(n_325), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_343), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_338), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_369), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_340), .B(n_323), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_340), .Y(n_374) );
INVx3_ASAP7_75t_L g375 ( .A(n_342), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_343), .Y(n_376) );
INVxp67_ASAP7_75t_SL g377 ( .A(n_353), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_357), .Y(n_378) );
OAI221xp5_ASAP7_75t_L g379 ( .A1(n_349), .A2(n_287), .B1(n_327), .B2(n_272), .C(n_297), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_344), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_344), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_354), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_364), .B(n_326), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_364), .A2(n_326), .B1(n_336), .B2(n_317), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_339), .B(n_336), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_361), .B(n_292), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_354), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_342), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_339), .B(n_336), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_355), .B(n_310), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_355), .B(n_310), .Y(n_391) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_342), .Y(n_392) );
INVx3_ASAP7_75t_L g393 ( .A(n_342), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_356), .B(n_320), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_356), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_358), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_358), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_373), .B(n_341), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_371), .Y(n_399) );
OA21x2_ASAP7_75t_L g400 ( .A1(n_370), .A2(n_346), .B(n_299), .Y(n_400) );
INVx2_ASAP7_75t_SL g401 ( .A(n_372), .Y(n_401) );
NAND4xp25_ASAP7_75t_L g402 ( .A(n_384), .B(n_348), .C(n_297), .D(n_368), .Y(n_402) );
AO22x1_ASAP7_75t_L g403 ( .A1(n_377), .A2(n_359), .B1(n_360), .B2(n_363), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_370), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_376), .Y(n_405) );
OA21x2_ASAP7_75t_L g406 ( .A1(n_376), .A2(n_346), .B(n_291), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_378), .Y(n_407) );
INVx3_ASAP7_75t_L g408 ( .A(n_388), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_371), .Y(n_409) );
INVx1_ASAP7_75t_SL g410 ( .A(n_378), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_380), .B(n_362), .Y(n_411) );
INVx3_ASAP7_75t_SL g412 ( .A(n_372), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_371), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_377), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_374), .A2(n_350), .B1(n_362), .B2(n_359), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_380), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_397), .B(n_363), .Y(n_417) );
BUFx3_ASAP7_75t_L g418 ( .A(n_372), .Y(n_418) );
OAI33xp33_ASAP7_75t_L g419 ( .A1(n_381), .A2(n_332), .A3(n_278), .B1(n_281), .B2(n_280), .B3(n_360), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_374), .B(n_368), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_381), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_382), .B(n_365), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_382), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g424 ( .A1(n_383), .A2(n_365), .B1(n_309), .B2(n_319), .C(n_288), .Y(n_424) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_383), .A2(n_314), .B1(n_301), .B2(n_303), .C(n_266), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_387), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_387), .Y(n_427) );
AO21x2_ASAP7_75t_L g428 ( .A1(n_395), .A2(n_285), .B(n_276), .Y(n_428) );
CKINVDCx5p33_ASAP7_75t_R g429 ( .A(n_386), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_395), .Y(n_430) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_394), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_416), .B(n_397), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_416), .B(n_396), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_404), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_414), .B(n_396), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_404), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_416), .B(n_394), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_399), .Y(n_438) );
NOR2xp33_ASAP7_75t_SL g439 ( .A(n_429), .B(n_366), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_415), .A2(n_379), .B1(n_391), .B2(n_390), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_398), .B(n_373), .Y(n_441) );
BUFx2_ASAP7_75t_L g442 ( .A(n_412), .Y(n_442) );
INVx2_ASAP7_75t_SL g443 ( .A(n_412), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_405), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_405), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_426), .B(n_385), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_431), .B(n_385), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_426), .B(n_389), .Y(n_448) );
AOI21xp33_ASAP7_75t_SL g449 ( .A1(n_403), .A2(n_379), .B(n_322), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_421), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_421), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_423), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_411), .B(n_417), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_411), .B(n_390), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_417), .B(n_391), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_410), .B(n_389), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_423), .Y(n_457) );
OAI211xp5_ASAP7_75t_L g458 ( .A1(n_402), .A2(n_306), .B(n_282), .C(n_321), .Y(n_458) );
INVx1_ASAP7_75t_SL g459 ( .A(n_412), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_430), .B(n_347), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_426), .B(n_375), .Y(n_461) );
NAND2x1p5_ASAP7_75t_L g462 ( .A(n_418), .B(n_369), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_424), .A2(n_293), .B(n_316), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_430), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_427), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_427), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_427), .B(n_367), .Y(n_467) );
AND2x4_ASAP7_75t_L g468 ( .A(n_418), .B(n_375), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_407), .B(n_347), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_422), .B(n_351), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_422), .Y(n_471) );
NOR2x1p5_ASAP7_75t_SL g472 ( .A(n_399), .B(n_351), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_399), .Y(n_473) );
AND2x4_ASAP7_75t_L g474 ( .A(n_418), .B(n_375), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_420), .B(n_413), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_409), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_420), .B(n_367), .Y(n_477) );
NAND2xp33_ASAP7_75t_L g478 ( .A(n_401), .B(n_392), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_409), .B(n_338), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_434), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_442), .B(n_401), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_436), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g483 ( .A(n_439), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_453), .B(n_475), .Y(n_484) );
NAND4xp25_ASAP7_75t_L g485 ( .A(n_440), .B(n_402), .C(n_425), .D(n_293), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_437), .B(n_403), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_437), .B(n_413), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_447), .B(n_413), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_471), .B(n_409), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_444), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_432), .B(n_406), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_445), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_450), .Y(n_493) );
AND2x4_ASAP7_75t_SL g494 ( .A(n_443), .B(n_408), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_451), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_435), .B(n_408), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_432), .B(n_406), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_452), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_438), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_433), .B(n_406), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_454), .B(n_408), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_457), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_464), .Y(n_503) );
NAND3xp33_ASAP7_75t_L g504 ( .A(n_469), .B(n_406), .C(n_400), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_433), .Y(n_505) );
NOR2xp67_ASAP7_75t_SL g506 ( .A(n_443), .B(n_369), .Y(n_506) );
INVx3_ASAP7_75t_L g507 ( .A(n_459), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_465), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_466), .B(n_400), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_455), .B(n_400), .Y(n_510) );
AND2x4_ASAP7_75t_L g511 ( .A(n_468), .B(n_474), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_446), .A2(n_419), .B1(n_375), .B2(n_393), .Y(n_512) );
BUFx3_ASAP7_75t_L g513 ( .A(n_462), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_438), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_446), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_473), .B(n_400), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_448), .B(n_408), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_473), .B(n_428), .Y(n_518) );
INVx2_ASAP7_75t_SL g519 ( .A(n_477), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_448), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_460), .Y(n_521) );
BUFx2_ASAP7_75t_L g522 ( .A(n_462), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_476), .Y(n_523) );
NOR2xp67_ASAP7_75t_SL g524 ( .A(n_458), .B(n_476), .Y(n_524) );
BUFx2_ASAP7_75t_L g525 ( .A(n_468), .Y(n_525) );
XNOR2x1_ASAP7_75t_L g526 ( .A(n_456), .B(n_315), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_467), .B(n_428), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_467), .B(n_428), .Y(n_528) );
INVx1_ASAP7_75t_SL g529 ( .A(n_478), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_470), .B(n_392), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_441), .B(n_392), .Y(n_531) );
INVx3_ASAP7_75t_L g532 ( .A(n_468), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_479), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_479), .B(n_392), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_461), .B(n_393), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_461), .B(n_393), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_517), .B(n_461), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_480), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_482), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_519), .B(n_474), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_485), .B(n_449), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_490), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_533), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_484), .B(n_474), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_515), .B(n_478), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_481), .B(n_472), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_492), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_493), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_495), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_508), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_520), .B(n_392), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_483), .B(n_463), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_505), .B(n_393), .Y(n_553) );
NAND2x1_ASAP7_75t_L g554 ( .A(n_507), .B(n_392), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_498), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_499), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_502), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_503), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_488), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_489), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_486), .B(n_388), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_489), .Y(n_562) );
INVxp67_ASAP7_75t_SL g563 ( .A(n_516), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_521), .B(n_388), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_487), .B(n_388), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_523), .B(n_388), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_511), .B(n_388), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_501), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_507), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_531), .B(n_320), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_514), .B(n_311), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_510), .B(n_311), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_510), .B(n_311), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_496), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_525), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_491), .B(n_328), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_491), .B(n_328), .Y(n_577) );
INVxp67_ASAP7_75t_SL g578 ( .A(n_516), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_509), .Y(n_579) );
CKINVDCx16_ASAP7_75t_R g580 ( .A(n_511), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_532), .B(n_328), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_530), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_509), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_494), .Y(n_584) );
INVxp67_ASAP7_75t_L g585 ( .A(n_524), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_497), .B(n_322), .Y(n_586) );
OAI21xp5_ASAP7_75t_SL g587 ( .A1(n_522), .A2(n_345), .B(n_352), .Y(n_587) );
AND2x4_ASAP7_75t_L g588 ( .A(n_532), .B(n_352), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_580), .B(n_534), .Y(n_589) );
OAI21xp5_ASAP7_75t_SL g590 ( .A1(n_585), .A2(n_481), .B(n_529), .Y(n_590) );
NOR3xp33_ASAP7_75t_L g591 ( .A(n_541), .B(n_504), .C(n_518), .Y(n_591) );
OAI211xp5_ASAP7_75t_L g592 ( .A1(n_541), .A2(n_513), .B(n_529), .C(n_512), .Y(n_592) );
AO21x1_ASAP7_75t_L g593 ( .A1(n_546), .A2(n_526), .B(n_518), .Y(n_593) );
NOR3xp33_ASAP7_75t_L g594 ( .A(n_552), .B(n_536), .C(n_535), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_568), .B(n_497), .Y(n_595) );
NAND4xp25_ASAP7_75t_L g596 ( .A(n_552), .B(n_536), .C(n_535), .D(n_528), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_559), .B(n_528), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_538), .Y(n_598) );
OAI21xp5_ASAP7_75t_SL g599 ( .A1(n_585), .A2(n_500), .B(n_527), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_560), .B(n_500), .Y(n_600) );
NOR2x1_ASAP7_75t_L g601 ( .A(n_587), .B(n_527), .Y(n_601) );
NAND4xp75_ASAP7_75t_L g602 ( .A(n_546), .B(n_506), .C(n_316), .D(n_263), .Y(n_602) );
NOR2x1_ASAP7_75t_L g603 ( .A(n_584), .B(n_352), .Y(n_603) );
AOI221xp5_ASAP7_75t_L g604 ( .A1(n_563), .A2(n_294), .B1(n_345), .B2(n_244), .C(n_352), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_537), .B(n_330), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_539), .Y(n_606) );
NOR3xp33_ASAP7_75t_SL g607 ( .A(n_540), .B(n_244), .C(n_283), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_562), .B(n_325), .Y(n_608) );
NOR3xp33_ASAP7_75t_L g609 ( .A(n_569), .B(n_330), .C(n_335), .Y(n_609) );
AOI311xp33_ASAP7_75t_L g610 ( .A1(n_574), .A2(n_258), .A3(n_267), .B(n_234), .C(n_274), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_563), .B(n_337), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_556), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_578), .B(n_337), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_578), .B(n_335), .Y(n_614) );
NOR3xp33_ASAP7_75t_SL g615 ( .A(n_572), .B(n_573), .C(n_576), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_537), .B(n_267), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_544), .B(n_234), .Y(n_617) );
NAND3xp33_ASAP7_75t_SL g618 ( .A(n_554), .B(n_313), .C(n_312), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_582), .B(n_313), .Y(n_619) );
OA211x2_ASAP7_75t_L g620 ( .A1(n_570), .A2(n_234), .B(n_231), .C(n_312), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_543), .B(n_302), .Y(n_621) );
OAI211xp5_ASAP7_75t_SL g622 ( .A1(n_575), .A2(n_255), .B(n_274), .C(n_302), .Y(n_622) );
NAND3xp33_ASAP7_75t_SL g623 ( .A(n_542), .B(n_241), .C(n_255), .Y(n_623) );
NAND3xp33_ASAP7_75t_SL g624 ( .A(n_547), .B(n_231), .C(n_234), .Y(n_624) );
NOR2x1_ASAP7_75t_L g625 ( .A(n_548), .B(n_248), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_594), .A2(n_545), .B1(n_561), .B2(n_588), .Y(n_626) );
NAND4xp25_ASAP7_75t_SL g627 ( .A(n_593), .B(n_549), .C(n_558), .D(n_557), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_591), .B(n_556), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_590), .A2(n_543), .B1(n_555), .B2(n_550), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_598), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_603), .A2(n_550), .B1(n_565), .B2(n_579), .Y(n_631) );
OAI21xp5_ASAP7_75t_L g632 ( .A1(n_625), .A2(n_564), .B(n_588), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_606), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_597), .B(n_595), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_612), .Y(n_635) );
INVxp67_ASAP7_75t_L g636 ( .A(n_601), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_589), .B(n_567), .Y(n_637) );
OAI21xp5_ASAP7_75t_SL g638 ( .A1(n_599), .A2(n_588), .B(n_551), .Y(n_638) );
INVx1_ASAP7_75t_SL g639 ( .A(n_605), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_600), .B(n_596), .Y(n_640) );
AND3x2_ASAP7_75t_L g641 ( .A(n_609), .B(n_581), .C(n_583), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_623), .A2(n_566), .B(n_579), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_611), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_613), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_623), .A2(n_583), .B(n_553), .Y(n_645) );
OAI21xp5_ASAP7_75t_L g646 ( .A1(n_592), .A2(n_577), .B(n_571), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_614), .B(n_586), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_615), .B(n_619), .Y(n_648) );
NAND4xp75_ASAP7_75t_L g649 ( .A(n_628), .B(n_620), .C(n_616), .D(n_604), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_640), .B(n_592), .Y(n_650) );
XNOR2x1_ASAP7_75t_L g651 ( .A(n_641), .B(n_602), .Y(n_651) );
NOR4xp75_ASAP7_75t_SL g652 ( .A(n_629), .B(n_608), .C(n_621), .D(n_610), .Y(n_652) );
OAI221xp5_ASAP7_75t_L g653 ( .A1(n_636), .A2(n_604), .B1(n_624), .B2(n_618), .C(n_617), .Y(n_653) );
NOR2x1_ASAP7_75t_L g654 ( .A(n_627), .B(n_624), .Y(n_654) );
NOR2x1p5_ASAP7_75t_L g655 ( .A(n_648), .B(n_607), .Y(n_655) );
XNOR2xp5_ASAP7_75t_L g656 ( .A(n_639), .B(n_622), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_637), .B(n_626), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_636), .B(n_630), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_634), .B(n_638), .Y(n_659) );
OAI211xp5_ASAP7_75t_SL g660 ( .A1(n_646), .A2(n_644), .B(n_643), .C(n_647), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_633), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_635), .B(n_631), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_661), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_662), .Y(n_664) );
NOR3xp33_ASAP7_75t_SL g665 ( .A(n_649), .B(n_632), .C(n_645), .Y(n_665) );
NOR3xp33_ASAP7_75t_SL g666 ( .A(n_650), .B(n_641), .C(n_642), .Y(n_666) );
A2O1A1Ixp33_ASAP7_75t_L g667 ( .A1(n_654), .A2(n_650), .B(n_659), .C(n_660), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_658), .Y(n_668) );
BUFx10_ASAP7_75t_L g669 ( .A(n_655), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_656), .Y(n_670) );
AOI211xp5_ASAP7_75t_L g671 ( .A1(n_667), .A2(n_653), .B(n_652), .C(n_657), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_664), .Y(n_672) );
NOR3xp33_ASAP7_75t_L g673 ( .A(n_670), .B(n_653), .C(n_651), .Y(n_673) );
XNOR2xp5_ASAP7_75t_L g674 ( .A(n_665), .B(n_666), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_672), .Y(n_675) );
NOR3x1_ASAP7_75t_L g676 ( .A(n_674), .B(n_669), .C(n_671), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_673), .Y(n_677) );
OAI21xp33_ASAP7_75t_L g678 ( .A1(n_677), .A2(n_666), .B(n_668), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_675), .A2(n_663), .B1(n_669), .B2(n_676), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_679), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_680), .A2(n_678), .B(n_675), .Y(n_681) );
endmodule