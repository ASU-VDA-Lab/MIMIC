module fake_jpeg_3708_n_401 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_401);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_401;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_4),
.B(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_0),
.B(n_12),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_45),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_14),
.B(n_1),
.C(n_4),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_46),
.B(n_84),
.Y(n_103)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_51),
.Y(n_142)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_55),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_14),
.B(n_1),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_56),
.B(n_64),
.Y(n_124)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_57),
.Y(n_147)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_58),
.Y(n_144)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_5),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_74),
.Y(n_116)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_37),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_75),
.B(n_76),
.Y(n_122)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx12_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_78),
.B(n_79),
.Y(n_139)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_80),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_44),
.B(n_5),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_82),
.Y(n_101)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_41),
.B(n_5),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_83),
.B(n_88),
.Y(n_107)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_21),
.B(n_7),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_86),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_36),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_89),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_31),
.B(n_7),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_15),
.B(n_30),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_91),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_94),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_38),
.B(n_15),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_95),
.Y(n_127)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_53),
.A2(n_43),
.B1(n_38),
.B2(n_27),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_98),
.A2(n_102),
.B1(n_110),
.B2(n_117),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_45),
.A2(n_20),
.B1(n_34),
.B2(n_33),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_54),
.A2(n_39),
.B1(n_40),
.B2(n_27),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_105),
.A2(n_125),
.B1(n_130),
.B2(n_146),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_65),
.A2(n_20),
.B1(n_34),
.B2(n_33),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_106),
.A2(n_109),
.B1(n_139),
.B2(n_135),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_79),
.A2(n_40),
.B1(n_32),
.B2(n_30),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_61),
.A2(n_95),
.B1(n_91),
.B2(n_90),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_66),
.A2(n_32),
.B1(n_18),
.B2(n_39),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_54),
.A2(n_18),
.B1(n_9),
.B2(n_10),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_63),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_130)
);

AND2x4_ASAP7_75t_L g132 ( 
.A(n_68),
.B(n_8),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_132),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_74),
.B(n_9),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_148),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_62),
.B(n_9),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_136),
.B(n_132),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_50),
.B(n_11),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_141),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_57),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_50),
.B(n_11),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_55),
.B(n_12),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_150),
.B(n_113),
.Y(n_182)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_152),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_106),
.A2(n_60),
.B1(n_86),
.B2(n_58),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_153),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_80),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_155),
.B(n_162),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_78),
.B1(n_71),
.B2(n_69),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_156),
.A2(n_180),
.B1(n_188),
.B2(n_190),
.Y(n_194)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_103),
.A2(n_70),
.B1(n_52),
.B2(n_67),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_158),
.A2(n_161),
.B1(n_156),
.B2(n_177),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_107),
.B(n_59),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_172),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_116),
.B(n_73),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_161),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_141),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_109),
.A2(n_84),
.B1(n_70),
.B2(n_13),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_132),
.A2(n_122),
.B1(n_116),
.B2(n_147),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_166),
.Y(n_227)
);

AO22x2_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_13),
.B1(n_141),
.B2(n_147),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_167),
.A2(n_129),
.B(n_140),
.Y(n_215)
);

BUFx6f_ASAP7_75t_SL g168 ( 
.A(n_111),
.Y(n_168)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_171),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_122),
.Y(n_172)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_174),
.Y(n_224)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_186),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_122),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_181),
.Y(n_199)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_178),
.B(n_184),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_101),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_189),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_97),
.A2(n_149),
.B1(n_99),
.B2(n_100),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_124),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_183),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_96),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

OR2x2_ASAP7_75t_SL g185 ( 
.A(n_104),
.B(n_118),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_129),
.B(n_120),
.C(n_108),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_99),
.B(n_118),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_142),
.A2(n_113),
.B1(n_145),
.B2(n_119),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_139),
.A2(n_112),
.B1(n_135),
.B2(n_121),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_142),
.B(n_139),
.C(n_144),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_120),
.Y(n_223)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_138),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_193),
.A2(n_140),
.B1(n_96),
.B2(n_137),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_155),
.A2(n_121),
.B1(n_112),
.B2(n_143),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_195),
.A2(n_200),
.B1(n_206),
.B2(n_211),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_104),
.B(n_113),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_205),
.A2(n_218),
.B(n_192),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_210),
.A2(n_173),
.B(n_172),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_193),
.A2(n_143),
.B1(n_140),
.B2(n_137),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_161),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_119),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_222),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_187),
.A2(n_129),
.B(n_108),
.Y(n_218)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

BUFx24_ASAP7_75t_SL g222 ( 
.A(n_181),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_176),
.C(n_191),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_228),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_162),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_232),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_194),
.A2(n_154),
.B1(n_157),
.B2(n_171),
.Y(n_231)
);

INVx11_ASAP7_75t_L g272 ( 
.A(n_231),
.Y(n_272)
);

AO21x1_ASAP7_75t_L g232 ( 
.A1(n_227),
.A2(n_160),
.B(n_151),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_226),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_241),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_186),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_238),
.Y(n_265)
);

O2A1O1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_215),
.A2(n_185),
.B(n_178),
.C(n_170),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_239),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_220),
.C(n_219),
.Y(n_269)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_167),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_252),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_200),
.A2(n_158),
.B1(n_179),
.B2(n_159),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_244),
.A2(n_198),
.B1(n_220),
.B2(n_202),
.Y(n_263)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_246),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_226),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_199),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_247),
.B(n_250),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_201),
.Y(n_248)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_248),
.Y(n_258)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_213),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_207),
.B(n_214),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_215),
.A2(n_227),
.B1(n_223),
.B2(n_198),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_197),
.A2(n_167),
.B1(n_183),
.B2(n_189),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_254),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_205),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_270),
.B1(n_271),
.B2(n_252),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_217),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_266),
.C(n_269),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_217),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_254),
.A2(n_218),
.B(n_210),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_267),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_244),
.A2(n_204),
.B1(n_212),
.B2(n_211),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_230),
.A2(n_204),
.B1(n_212),
.B2(n_195),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_237),
.B(n_167),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_167),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_233),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_279),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_233),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_273),
.Y(n_280)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_280),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_281),
.A2(n_287),
.B1(n_288),
.B2(n_257),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_268),
.Y(n_282)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_282),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_247),
.Y(n_284)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_284),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_276),
.A2(n_230),
.B1(n_236),
.B2(n_243),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_286),
.A2(n_298),
.B1(n_281),
.B2(n_267),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_276),
.A2(n_242),
.B1(n_236),
.B2(n_243),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_261),
.A2(n_243),
.B1(n_251),
.B2(n_254),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_235),
.B1(n_246),
.B2(n_250),
.Y(n_289)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_289),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_278),
.B(n_234),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_290),
.Y(n_303)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_291),
.Y(n_314)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_292),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_228),
.C(n_239),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_296),
.C(n_300),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_263),
.B(n_234),
.Y(n_295)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_295),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_241),
.C(n_245),
.Y(n_296)
);

OAI32xp33_ASAP7_75t_L g297 ( 
.A1(n_265),
.A2(n_238),
.A3(n_249),
.B1(n_232),
.B2(n_184),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_265),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_277),
.A2(n_238),
.B1(n_232),
.B2(n_196),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_260),
.Y(n_299)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_299),
.Y(n_320)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_255),
.Y(n_301)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_302),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_288),
.A2(n_262),
.B1(n_256),
.B2(n_277),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_304),
.B(n_279),
.Y(n_336)
);

AOI21x1_ASAP7_75t_SL g334 ( 
.A1(n_305),
.A2(n_312),
.B(n_316),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_283),
.B(n_266),
.C(n_256),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_313),
.C(n_287),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_310),
.A2(n_272),
.B1(n_258),
.B2(n_248),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_294),
.A2(n_261),
.B(n_260),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_283),
.B(n_296),
.C(n_293),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_294),
.A2(n_297),
.B(n_298),
.Y(n_316)
);

O2A1O1Ixp33_ASAP7_75t_L g319 ( 
.A1(n_292),
.A2(n_272),
.B(n_270),
.C(n_271),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_319),
.A2(n_286),
.B(n_285),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_259),
.Y(n_322)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_322),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_323),
.B(n_328),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_280),
.Y(n_325)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_325),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_326),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_300),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_327),
.B(n_329),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_306),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_274),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_312),
.B(n_291),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_330),
.B(n_320),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_311),
.A2(n_285),
.B(n_301),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_331),
.A2(n_337),
.B1(n_338),
.B2(n_315),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_224),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_332),
.B(n_333),
.C(n_320),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_304),
.B(n_224),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_336),
.A2(n_305),
.B1(n_310),
.B2(n_309),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_311),
.A2(n_275),
.B(n_255),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_322),
.Y(n_339)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_339),
.Y(n_347)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_317),
.Y(n_340)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_340),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_342),
.B(n_314),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_344),
.B(n_333),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_346),
.A2(n_349),
.B1(n_351),
.B2(n_330),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_324),
.A2(n_316),
.B1(n_318),
.B2(n_317),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_335),
.Y(n_350)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_350),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_326),
.A2(n_318),
.B1(n_303),
.B2(n_319),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_309),
.C(n_321),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_352),
.B(n_327),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_353),
.A2(n_319),
.B1(n_334),
.B2(n_307),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_356),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_357),
.A2(n_349),
.B1(n_346),
.B2(n_344),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_341),
.A2(n_334),
.B(n_323),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_358),
.A2(n_343),
.B(n_225),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_345),
.A2(n_332),
.B(n_338),
.Y(n_359)
);

AOI21x1_ASAP7_75t_SL g371 ( 
.A1(n_359),
.A2(n_347),
.B(n_348),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_362),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_352),
.B(n_329),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_361),
.B(n_364),
.C(n_365),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_351),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_363),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_354),
.B(n_314),
.C(n_307),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_354),
.B(n_315),
.C(n_225),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_363),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_374),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_365),
.B(n_364),
.C(n_361),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_375),
.Y(n_383)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_370),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_371),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_357),
.A2(n_343),
.B(n_258),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_373),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_377),
.B(n_380),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_369),
.B(n_356),
.C(n_359),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_368),
.B(n_366),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_381),
.B(n_382),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_368),
.B(n_248),
.Y(n_382)
);

AOI21x1_ASAP7_75t_L g385 ( 
.A1(n_379),
.A2(n_372),
.B(n_374),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_385),
.A2(n_386),
.B(n_389),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_383),
.A2(n_371),
.B(n_367),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_378),
.A2(n_376),
.B(n_201),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_380),
.B(n_201),
.C(n_165),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_390),
.B(n_164),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_387),
.A2(n_384),
.B(n_221),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_391),
.A2(n_392),
.B(n_221),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_388),
.B(n_384),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_393),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_395),
.A2(n_397),
.B(n_114),
.Y(n_399)
);

AOI21x1_ASAP7_75t_L g397 ( 
.A1(n_394),
.A2(n_174),
.B(n_175),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_396),
.A2(n_152),
.B1(n_203),
.B2(n_138),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_398),
.B(n_399),
.C(n_203),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_400),
.A2(n_114),
.B1(n_168),
.B2(n_138),
.Y(n_401)
);


endmodule