module fake_netlist_5_2435_n_3389 (n_137, n_924, n_676, n_294, n_431, n_318, n_380, n_419, n_977, n_653, n_611, n_444, n_642, n_469, n_615, n_851, n_82, n_194, n_316, n_785, n_389, n_843, n_855, n_549, n_684, n_850, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_705, n_619, n_408, n_865, n_61, n_913, n_678, n_664, n_376, n_697, n_503, n_967, n_127, n_75, n_235, n_226, n_605, n_74, n_776, n_928, n_667, n_515, n_790, n_57, n_353, n_351, n_367, n_620, n_643, n_916, n_452, n_885, n_397, n_493, n_111, n_525, n_880, n_703, n_698, n_980, n_483, n_544, n_683, n_155, n_780, n_649, n_552, n_547, n_43, n_721, n_116, n_841, n_956, n_22, n_467, n_564, n_802, n_423, n_840, n_284, n_46, n_245, n_21, n_501, n_823, n_725, n_983, n_139, n_38, n_105, n_280, n_744, n_590, n_629, n_672, n_4, n_873, n_378, n_551, n_762, n_17, n_581, n_688, n_382, n_554, n_800, n_898, n_254, n_690, n_33, n_23, n_583, n_671, n_718, n_819, n_302, n_265, n_526, n_915, n_719, n_293, n_372, n_443, n_244, n_677, n_47, n_173, n_859, n_864, n_951, n_821, n_198, n_714, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_909, n_625, n_854, n_949, n_621, n_753, n_100, n_455, n_674, n_932, n_417, n_946, n_612, n_212, n_385, n_498, n_516, n_933, n_788, n_507, n_119, n_497, n_689, n_738, n_912, n_606, n_559, n_275, n_640, n_968, n_252, n_624, n_825, n_26, n_295, n_133, n_330, n_877, n_508, n_739, n_506, n_2, n_737, n_610, n_972, n_692, n_986, n_755, n_6, n_509, n_568, n_936, n_39, n_147, n_373, n_820, n_757, n_947, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_758, n_668, n_733, n_991, n_375, n_301, n_828, n_779, n_576, n_941, n_929, n_981, n_68, n_804, n_93, n_867, n_186, n_537, n_134, n_902, n_191, n_587, n_945, n_659, n_51, n_63, n_492, n_792, n_563, n_171, n_153, n_756, n_878, n_524, n_943, n_399, n_341, n_204, n_394, n_250, n_579, n_992, n_938, n_741, n_548, n_543, n_260, n_812, n_842, n_298, n_650, n_984, n_320, n_694, n_518, n_505, n_286, n_883, n_122, n_282, n_752, n_331, n_10, n_905, n_906, n_24, n_406, n_519, n_470, n_908, n_782, n_919, n_325, n_449, n_132, n_862, n_90, n_900, n_724, n_856, n_546, n_101, n_760, n_658, n_281, n_918, n_240, n_942, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_731, n_31, n_456, n_13, n_371, n_959, n_481, n_535, n_709, n_152, n_540, n_317, n_618, n_940, n_896, n_9, n_323, n_569, n_769, n_195, n_42, n_356, n_227, n_592, n_45, n_920, n_894, n_271, n_934, n_94, n_831, n_826, n_335, n_123, n_886, n_978, n_964, n_654, n_370, n_167, n_976, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_833, n_297, n_156, n_5, n_853, n_603, n_225, n_377, n_751, n_484, n_775, n_219, n_988, n_442, n_157, n_814, n_131, n_192, n_636, n_786, n_600, n_660, n_223, n_392, n_158, n_655, n_704, n_787, n_138, n_264, n_109, n_669, n_472, n_742, n_750, n_454, n_961, n_955, n_387, n_771, n_374, n_163, n_276, n_339, n_95, n_882, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_763, n_169, n_59, n_522, n_550, n_255, n_696, n_897, n_215, n_350, n_196, n_798, n_662, n_459, n_646, n_211, n_218, n_400, n_930, n_181, n_436, n_962, n_3, n_290, n_580, n_221, n_178, n_622, n_723, n_386, n_578, n_926, n_287, n_344, n_848, n_555, n_783, n_473, n_422, n_475, n_777, n_72, n_661, n_104, n_41, n_682, n_415, n_56, n_141, n_485, n_496, n_355, n_958, n_849, n_486, n_670, n_15, n_816, n_336, n_584, n_681, n_591, n_922, n_145, n_48, n_521, n_614, n_663, n_845, n_50, n_337, n_430, n_313, n_631, n_673, n_837, n_88, n_479, n_528, n_510, n_216, n_680, n_168, n_974, n_395, n_164, n_432, n_553, n_727, n_839, n_901, n_311, n_813, n_957, n_830, n_773, n_208, n_142, n_743, n_214, n_328, n_140, n_801, n_299, n_303, n_369, n_675, n_888, n_296, n_613, n_871, n_241, n_637, n_357, n_875, n_598, n_685, n_608, n_184, n_446, n_445, n_65, n_78, n_749, n_829, n_144, n_858, n_114, n_96, n_923, n_772, n_691, n_881, n_717, n_165, n_468, n_499, n_939, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_789, n_363, n_402, n_413, n_734, n_638, n_700, n_197, n_796, n_107, n_573, n_69, n_866, n_969, n_236, n_388, n_761, n_1, n_249, n_903, n_740, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_889, n_80, n_973, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_693, n_309, n_30, n_512, n_14, n_836, n_990, n_84, n_462, n_975, n_130, n_322, n_567, n_258, n_652, n_778, n_29, n_79, n_151, n_25, n_306, n_907, n_722, n_458, n_288, n_770, n_188, n_190, n_844, n_201, n_263, n_471, n_609, n_852, n_989, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_711, n_781, n_834, n_474, n_112, n_765, n_542, n_85, n_463, n_488, n_595, n_736, n_502, n_892, n_893, n_891, n_239, n_466, n_420, n_630, n_489, n_632, n_699, n_55, n_979, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_748, n_586, n_846, n_874, n_465, n_838, n_76, n_358, n_362, n_876, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_953, n_601, n_279, n_917, n_966, n_70, n_987, n_253, n_261, n_174, n_289, n_745, n_963, n_954, n_627, n_767, n_172, n_206, n_217, n_440, n_726, n_478, n_793, n_545, n_982, n_441, n_860, n_450, n_648, n_312, n_476, n_818, n_429, n_861, n_534, n_948, n_884, n_899, n_345, n_210, n_944, n_494, n_641, n_628, n_365, n_774, n_91, n_729, n_730, n_176, n_970, n_911, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_679, n_707, n_710, n_795, n_695, n_832, n_180, n_857, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_937, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_879, n_16, n_720, n_0, n_58, n_623, n_405, n_824, n_18, n_359, n_863, n_910, n_971, n_490, n_805, n_117, n_326, n_794, n_768, n_921, n_233, n_404, n_686, n_205, n_366, n_572, n_113, n_712, n_754, n_847, n_815, n_246, n_596, n_179, n_125, n_410, n_558, n_708, n_269, n_529, n_128, n_735, n_702, n_285, n_822, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_728, n_895, n_202, n_266, n_272, n_491, n_427, n_791, n_732, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_808, n_409, n_797, n_887, n_589, n_716, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_809, n_870, n_931, n_159, n_334, n_599, n_766, n_811, n_952, n_541, n_807, n_391, n_701, n_434, n_645, n_539, n_835, n_175, n_538, n_666, n_262, n_803, n_868, n_238, n_639, n_799, n_914, n_99, n_687, n_715, n_411, n_414, n_319, n_364, n_965, n_927, n_20, n_536, n_531, n_935, n_121, n_242, n_817, n_872, n_360, n_36, n_594, n_764, n_200, n_890, n_162, n_960, n_64, n_759, n_222, n_28, n_89, n_438, n_806, n_115, n_713, n_904, n_985, n_869, n_324, n_810, n_634, n_416, n_199, n_827, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_925, n_424, n_7, n_706, n_746, n_256, n_305, n_533, n_950, n_747, n_52, n_278, n_784, n_110, n_3389);

input n_137;
input n_924;
input n_676;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_977;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_851;
input n_82;
input n_194;
input n_316;
input n_785;
input n_389;
input n_843;
input n_855;
input n_549;
input n_684;
input n_850;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_705;
input n_619;
input n_408;
input n_865;
input n_61;
input n_913;
input n_678;
input n_664;
input n_376;
input n_697;
input n_503;
input n_967;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_776;
input n_928;
input n_667;
input n_515;
input n_790;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_916;
input n_452;
input n_885;
input n_397;
input n_493;
input n_111;
input n_525;
input n_880;
input n_703;
input n_698;
input n_980;
input n_483;
input n_544;
input n_683;
input n_155;
input n_780;
input n_649;
input n_552;
input n_547;
input n_43;
input n_721;
input n_116;
input n_841;
input n_956;
input n_22;
input n_467;
input n_564;
input n_802;
input n_423;
input n_840;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_823;
input n_725;
input n_983;
input n_139;
input n_38;
input n_105;
input n_280;
input n_744;
input n_590;
input n_629;
input n_672;
input n_4;
input n_873;
input n_378;
input n_551;
input n_762;
input n_17;
input n_581;
input n_688;
input n_382;
input n_554;
input n_800;
input n_898;
input n_254;
input n_690;
input n_33;
input n_23;
input n_583;
input n_671;
input n_718;
input n_819;
input n_302;
input n_265;
input n_526;
input n_915;
input n_719;
input n_293;
input n_372;
input n_443;
input n_244;
input n_677;
input n_47;
input n_173;
input n_859;
input n_864;
input n_951;
input n_821;
input n_198;
input n_714;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_909;
input n_625;
input n_854;
input n_949;
input n_621;
input n_753;
input n_100;
input n_455;
input n_674;
input n_932;
input n_417;
input n_946;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_933;
input n_788;
input n_507;
input n_119;
input n_497;
input n_689;
input n_738;
input n_912;
input n_606;
input n_559;
input n_275;
input n_640;
input n_968;
input n_252;
input n_624;
input n_825;
input n_26;
input n_295;
input n_133;
input n_330;
input n_877;
input n_508;
input n_739;
input n_506;
input n_2;
input n_737;
input n_610;
input n_972;
input n_692;
input n_986;
input n_755;
input n_6;
input n_509;
input n_568;
input n_936;
input n_39;
input n_147;
input n_373;
input n_820;
input n_757;
input n_947;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_758;
input n_668;
input n_733;
input n_991;
input n_375;
input n_301;
input n_828;
input n_779;
input n_576;
input n_941;
input n_929;
input n_981;
input n_68;
input n_804;
input n_93;
input n_867;
input n_186;
input n_537;
input n_134;
input n_902;
input n_191;
input n_587;
input n_945;
input n_659;
input n_51;
input n_63;
input n_492;
input n_792;
input n_563;
input n_171;
input n_153;
input n_756;
input n_878;
input n_524;
input n_943;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_992;
input n_938;
input n_741;
input n_548;
input n_543;
input n_260;
input n_812;
input n_842;
input n_298;
input n_650;
input n_984;
input n_320;
input n_694;
input n_518;
input n_505;
input n_286;
input n_883;
input n_122;
input n_282;
input n_752;
input n_331;
input n_10;
input n_905;
input n_906;
input n_24;
input n_406;
input n_519;
input n_470;
input n_908;
input n_782;
input n_919;
input n_325;
input n_449;
input n_132;
input n_862;
input n_90;
input n_900;
input n_724;
input n_856;
input n_546;
input n_101;
input n_760;
input n_658;
input n_281;
input n_918;
input n_240;
input n_942;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_731;
input n_31;
input n_456;
input n_13;
input n_371;
input n_959;
input n_481;
input n_535;
input n_709;
input n_152;
input n_540;
input n_317;
input n_618;
input n_940;
input n_896;
input n_9;
input n_323;
input n_569;
input n_769;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_920;
input n_894;
input n_271;
input n_934;
input n_94;
input n_831;
input n_826;
input n_335;
input n_123;
input n_886;
input n_978;
input n_964;
input n_654;
input n_370;
input n_167;
input n_976;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_833;
input n_297;
input n_156;
input n_5;
input n_853;
input n_603;
input n_225;
input n_377;
input n_751;
input n_484;
input n_775;
input n_219;
input n_988;
input n_442;
input n_157;
input n_814;
input n_131;
input n_192;
input n_636;
input n_786;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_704;
input n_787;
input n_138;
input n_264;
input n_109;
input n_669;
input n_472;
input n_742;
input n_750;
input n_454;
input n_961;
input n_955;
input n_387;
input n_771;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_882;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_763;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_696;
input n_897;
input n_215;
input n_350;
input n_196;
input n_798;
input n_662;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_930;
input n_181;
input n_436;
input n_962;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_723;
input n_386;
input n_578;
input n_926;
input n_287;
input n_344;
input n_848;
input n_555;
input n_783;
input n_473;
input n_422;
input n_475;
input n_777;
input n_72;
input n_661;
input n_104;
input n_41;
input n_682;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_958;
input n_849;
input n_486;
input n_670;
input n_15;
input n_816;
input n_336;
input n_584;
input n_681;
input n_591;
input n_922;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_845;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_673;
input n_837;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_680;
input n_168;
input n_974;
input n_395;
input n_164;
input n_432;
input n_553;
input n_727;
input n_839;
input n_901;
input n_311;
input n_813;
input n_957;
input n_830;
input n_773;
input n_208;
input n_142;
input n_743;
input n_214;
input n_328;
input n_140;
input n_801;
input n_299;
input n_303;
input n_369;
input n_675;
input n_888;
input n_296;
input n_613;
input n_871;
input n_241;
input n_637;
input n_357;
input n_875;
input n_598;
input n_685;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_749;
input n_829;
input n_144;
input n_858;
input n_114;
input n_96;
input n_923;
input n_772;
input n_691;
input n_881;
input n_717;
input n_165;
input n_468;
input n_499;
input n_939;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_789;
input n_363;
input n_402;
input n_413;
input n_734;
input n_638;
input n_700;
input n_197;
input n_796;
input n_107;
input n_573;
input n_69;
input n_866;
input n_969;
input n_236;
input n_388;
input n_761;
input n_1;
input n_249;
input n_903;
input n_740;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_889;
input n_80;
input n_973;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_693;
input n_309;
input n_30;
input n_512;
input n_14;
input n_836;
input n_990;
input n_84;
input n_462;
input n_975;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_778;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_907;
input n_722;
input n_458;
input n_288;
input n_770;
input n_188;
input n_190;
input n_844;
input n_201;
input n_263;
input n_471;
input n_609;
input n_852;
input n_989;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_711;
input n_781;
input n_834;
input n_474;
input n_112;
input n_765;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_736;
input n_502;
input n_892;
input n_893;
input n_891;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_699;
input n_55;
input n_979;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_748;
input n_586;
input n_846;
input n_874;
input n_465;
input n_838;
input n_76;
input n_358;
input n_362;
input n_876;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_953;
input n_601;
input n_279;
input n_917;
input n_966;
input n_70;
input n_987;
input n_253;
input n_261;
input n_174;
input n_289;
input n_745;
input n_963;
input n_954;
input n_627;
input n_767;
input n_172;
input n_206;
input n_217;
input n_440;
input n_726;
input n_478;
input n_793;
input n_545;
input n_982;
input n_441;
input n_860;
input n_450;
input n_648;
input n_312;
input n_476;
input n_818;
input n_429;
input n_861;
input n_534;
input n_948;
input n_884;
input n_899;
input n_345;
input n_210;
input n_944;
input n_494;
input n_641;
input n_628;
input n_365;
input n_774;
input n_91;
input n_729;
input n_730;
input n_176;
input n_970;
input n_911;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_679;
input n_707;
input n_710;
input n_795;
input n_695;
input n_832;
input n_180;
input n_857;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_937;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_879;
input n_16;
input n_720;
input n_0;
input n_58;
input n_623;
input n_405;
input n_824;
input n_18;
input n_359;
input n_863;
input n_910;
input n_971;
input n_490;
input n_805;
input n_117;
input n_326;
input n_794;
input n_768;
input n_921;
input n_233;
input n_404;
input n_686;
input n_205;
input n_366;
input n_572;
input n_113;
input n_712;
input n_754;
input n_847;
input n_815;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_708;
input n_269;
input n_529;
input n_128;
input n_735;
input n_702;
input n_285;
input n_822;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_728;
input n_895;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_791;
input n_732;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_808;
input n_409;
input n_797;
input n_887;
input n_589;
input n_716;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_809;
input n_870;
input n_931;
input n_159;
input n_334;
input n_599;
input n_766;
input n_811;
input n_952;
input n_541;
input n_807;
input n_391;
input n_701;
input n_434;
input n_645;
input n_539;
input n_835;
input n_175;
input n_538;
input n_666;
input n_262;
input n_803;
input n_868;
input n_238;
input n_639;
input n_799;
input n_914;
input n_99;
input n_687;
input n_715;
input n_411;
input n_414;
input n_319;
input n_364;
input n_965;
input n_927;
input n_20;
input n_536;
input n_531;
input n_935;
input n_121;
input n_242;
input n_817;
input n_872;
input n_360;
input n_36;
input n_594;
input n_764;
input n_200;
input n_890;
input n_162;
input n_960;
input n_64;
input n_759;
input n_222;
input n_28;
input n_89;
input n_438;
input n_806;
input n_115;
input n_713;
input n_904;
input n_985;
input n_869;
input n_324;
input n_810;
input n_634;
input n_416;
input n_199;
input n_827;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_925;
input n_424;
input n_7;
input n_706;
input n_746;
input n_256;
input n_305;
input n_533;
input n_950;
input n_747;
input n_52;
input n_278;
input n_784;
input n_110;

output n_3389;

wire n_1263;
wire n_3304;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_1423;
wire n_1126;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_3241;
wire n_2617;
wire n_2200;
wire n_3261;
wire n_3006;
wire n_1161;
wire n_3027;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_3179;
wire n_3127;
wire n_1780;
wire n_3256;
wire n_1488;
wire n_2899;
wire n_2955;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_3086;
wire n_3297;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_3088;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_2853;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_3246;
wire n_3202;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_1545;
wire n_2374;
wire n_3341;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_3019;
wire n_3039;
wire n_2011;
wire n_2096;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_3163;
wire n_1118;
wire n_1686;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1728;
wire n_1107;
wire n_2076;
wire n_2031;
wire n_2482;
wire n_3036;
wire n_2677;
wire n_1230;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_3010;
wire n_3180;
wire n_3379;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_3188;
wire n_3325;
wire n_3107;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_1098;
wire n_2963;
wire n_2142;
wire n_3186;
wire n_3082;
wire n_1154;
wire n_2189;
wire n_3332;
wire n_1242;
wire n_3283;
wire n_1135;
wire n_3048;
wire n_3258;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_2959;
wire n_3340;
wire n_2047;
wire n_1280;
wire n_3277;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_1483;
wire n_2888;
wire n_1314;
wire n_1512;
wire n_3157;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2983;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_3214;
wire n_2306;
wire n_2515;
wire n_3022;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2635;
wire n_2652;
wire n_2715;
wire n_3087;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_3060;
wire n_2651;
wire n_1484;
wire n_2071;
wire n_2643;
wire n_1374;
wire n_1328;
wire n_2561;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_3183;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_3353;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_3049;
wire n_1723;
wire n_1850;
wire n_3028;
wire n_1146;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_3156;
wire n_3101;
wire n_3376;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_2976;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_3089;
wire n_1547;
wire n_1070;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_3222;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_1801;
wire n_1391;
wire n_1034;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_3361;
wire n_1600;
wire n_2235;
wire n_1862;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_3291;
wire n_1473;
wire n_1587;
wire n_2682;
wire n_2432;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_2934;
wire n_1672;
wire n_2506;
wire n_2699;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_2079;
wire n_2238;
wire n_2118;
wire n_1151;
wire n_2985;
wire n_2944;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_2932;
wire n_2753;
wire n_2980;
wire n_1582;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_3262;
wire n_3136;
wire n_1836;
wire n_2868;
wire n_1450;
wire n_3141;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_3164;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_2358;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_3191;
wire n_1585;
wire n_2684;
wire n_2712;
wire n_3193;
wire n_1971;
wire n_1599;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_3367;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_1447;
wire n_2251;
wire n_3096;
wire n_1377;
wire n_2370;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_3339;
wire n_2055;
wire n_3025;
wire n_3349;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_3320;
wire n_3007;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_3071;
wire n_3310;
wire n_2258;
wire n_1667;
wire n_1058;
wire n_3359;
wire n_2784;
wire n_2919;
wire n_3092;
wire n_1053;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_3146;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_1052;
wire n_1385;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_2987;
wire n_1527;
wire n_2042;
wire n_3106;
wire n_1882;
wire n_3328;
wire n_1754;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2674;
wire n_2606;
wire n_3187;
wire n_1565;
wire n_2828;
wire n_3371;
wire n_1809;
wire n_1856;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_3208;
wire n_1319;
wire n_2379;
wire n_3331;
wire n_2616;
wire n_2911;
wire n_3305;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_3257;
wire n_1027;
wire n_1156;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2293;
wire n_2837;
wire n_1393;
wire n_2319;
wire n_1775;
wire n_2979;
wire n_3296;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_2808;
wire n_1276;
wire n_3009;
wire n_2548;
wire n_1412;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_2108;
wire n_1538;
wire n_1162;
wire n_2930;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_2967;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_1905;
wire n_2553;
wire n_3207;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_3224;
wire n_2698;
wire n_1711;
wire n_1891;
wire n_1662;
wire n_1481;
wire n_2626;
wire n_3042;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_3047;
wire n_2454;
wire n_2804;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_3120;
wire n_1876;
wire n_1743;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_2222;
wire n_1892;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_3218;
wire n_1477;
wire n_3142;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_3119;
wire n_1189;
wire n_2690;
wire n_3370;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_1649;
wire n_3150;
wire n_2064;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_3279;
wire n_2621;
wire n_1759;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_1537;
wire n_2227;
wire n_2671;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_3346;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_3133;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_2992;
wire n_1674;
wire n_1833;
wire n_3138;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_3128;
wire n_1734;
wire n_3038;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_3068;
wire n_1767;
wire n_3144;
wire n_2943;
wire n_2913;
wire n_2336;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_3317;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_3355;
wire n_2007;
wire n_3220;
wire n_2539;
wire n_3263;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_3158;
wire n_1624;
wire n_3000;
wire n_1510;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_1406;
wire n_1279;
wire n_3113;
wire n_3108;
wire n_3111;
wire n_2718;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_2577;
wire n_1760;
wire n_2875;
wire n_1500;
wire n_2960;
wire n_1090;
wire n_2796;
wire n_3280;
wire n_2342;
wire n_2856;
wire n_1832;
wire n_1851;
wire n_999;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_2937;
wire n_3003;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_3288;
wire n_1158;
wire n_3095;
wire n_2045;
wire n_3369;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_3199;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_3030;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_1163;
wire n_3271;
wire n_2039;
wire n_1207;
wire n_2412;
wire n_2406;
wire n_2846;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_2035;
wire n_2061;
wire n_3075;
wire n_3173;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_3236;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_2459;
wire n_3031;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_3243;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_2982;
wire n_3385;
wire n_1017;
wire n_2481;
wire n_2947;
wire n_2171;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_3343;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_1079;
wire n_2320;
wire n_2339;
wire n_1045;
wire n_1208;
wire n_2473;
wire n_2038;
wire n_3287;
wire n_2137;
wire n_3378;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_2029;
wire n_995;
wire n_3221;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_3021;
wire n_1989;
wire n_2359;
wire n_2941;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_3098;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_2312;
wire n_1215;
wire n_3015;
wire n_1171;
wire n_1578;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_3058;
wire n_2812;
wire n_2048;
wire n_3197;
wire n_3109;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_3002;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_3276;
wire n_1355;
wire n_2565;
wire n_1159;
wire n_2124;
wire n_3001;
wire n_2081;
wire n_3149;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_3268;
wire n_2418;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_3301;
wire n_1237;
wire n_1420;
wire n_3185;
wire n_1132;
wire n_3330;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_3248;
wire n_2277;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_2090;
wire n_3374;
wire n_3153;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_2896;
wire n_1111;
wire n_3213;
wire n_1365;
wire n_1927;
wire n_3065;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_1041;
wire n_1265;
wire n_3223;
wire n_1909;
wire n_3077;
wire n_2681;
wire n_1562;
wire n_3103;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_1015;
wire n_1140;
wire n_1651;
wire n_1965;
wire n_3387;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_1823;
wire n_2464;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_3189;
wire n_1846;
wire n_3037;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_3154;
wire n_3229;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_1849;
wire n_2410;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_1935;
wire n_2922;
wire n_1430;
wire n_3275;
wire n_2645;
wire n_2467;
wire n_3366;
wire n_2727;
wire n_1094;
wire n_1534;
wire n_1354;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1205;
wire n_1044;
wire n_2436;
wire n_1209;
wire n_3029;
wire n_1552;
wire n_2508;
wire n_3242;
wire n_2593;
wire n_1435;
wire n_2416;
wire n_2405;
wire n_3286;
wire n_2088;
wire n_2953;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_996;
wire n_1684;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_3097;
wire n_1821;
wire n_2929;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_3388;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2890;
wire n_3059;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_3215;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_1436;
wire n_1691;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_3171;
wire n_1229;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_2216;
wire n_3020;
wire n_1757;
wire n_1897;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_2933;
wire n_2308;
wire n_1893;
wire n_2910;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_1206;
wire n_2647;
wire n_3160;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_2969;
wire n_3195;
wire n_1519;
wire n_3190;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_1346;
wire n_3053;
wire n_1299;
wire n_3244;
wire n_2158;
wire n_1808;
wire n_3290;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_3130;
wire n_2465;
wire n_2824;
wire n_3033;
wire n_2650;
wire n_3298;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_3334;
wire n_1442;
wire n_2923;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_3264;
wire n_2333;
wire n_2916;
wire n_3166;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_1632;
wire n_3110;
wire n_2998;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_2402;
wire n_1157;
wire n_3073;
wire n_2403;
wire n_1050;
wire n_1954;
wire n_2265;
wire n_3162;
wire n_1608;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_3377;
wire n_2870;
wire n_1305;
wire n_3178;
wire n_1826;
wire n_1112;
wire n_3134;
wire n_2304;
wire n_2999;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_3362;
wire n_2881;
wire n_1631;
wire n_1203;
wire n_3282;
wire n_2472;
wire n_1763;
wire n_2341;
wire n_3105;
wire n_3231;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_2993;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_3274;
wire n_3041;
wire n_3299;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_3209;
wire n_2037;
wire n_2685;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_3203;
wire n_1301;
wire n_1668;
wire n_1363;
wire n_1185;
wire n_2903;
wire n_1967;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_3255;
wire n_1439;
wire n_1312;
wire n_2827;
wire n_1688;
wire n_3052;
wire n_2997;
wire n_3327;
wire n_1504;
wire n_3326;
wire n_3067;
wire n_1932;
wire n_3375;
wire n_2755;
wire n_3237;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_1983;
wire n_3167;
wire n_1594;
wire n_1400;
wire n_1342;
wire n_1214;
wire n_2362;
wire n_2609;
wire n_1793;
wire n_3382;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1422;
wire n_1077;
wire n_3196;
wire n_3078;
wire n_2364;
wire n_2533;
wire n_3094;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_3316;
wire n_2291;
wire n_3099;
wire n_2596;
wire n_1636;
wire n_2056;
wire n_3253;
wire n_1730;
wire n_2280;
wire n_2192;
wire n_3363;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_2973;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_2974;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_3372;
wire n_2971;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_3240;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_3147;
wire n_2758;
wire n_1458;
wire n_2471;
wire n_1472;
wire n_1176;
wire n_2298;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_2559;
wire n_3230;
wire n_1020;
wire n_1062;
wire n_3342;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_3386;
wire n_1204;
wire n_2840;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_2893;
wire n_1188;
wire n_2588;
wire n_2962;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_2600;
wire n_2795;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_2002;
wire n_2282;
wire n_2800;
wire n_2371;
wire n_2935;
wire n_3233;
wire n_3380;
wire n_3177;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_3085;
wire n_2444;
wire n_2068;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_3123;
wire n_3137;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_1603;
wire n_1232;
wire n_2638;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_2270;
wire n_1506;
wire n_3206;
wire n_2653;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_1465;
wire n_3145;
wire n_3124;
wire n_1122;
wire n_3192;
wire n_2608;
wire n_2657;
wire n_2995;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2852;
wire n_2392;
wire n_3093;
wire n_1843;
wire n_1499;
wire n_3061;
wire n_3155;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_3324;
wire n_3356;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_3182;
wire n_1572;
wire n_1968;
wire n_3269;
wire n_2564;
wire n_2252;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_1714;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_3174;
wire n_2575;
wire n_2988;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_2373;
wire n_1970;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2722;
wire n_2117;
wire n_2745;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1514;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_1345;
wire n_1059;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_3226;
wire n_1410;
wire n_1005;
wire n_1003;
wire n_3090;
wire n_2067;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_2877;
wire n_3318;
wire n_2148;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_1584;
wire n_1726;
wire n_1835;
wire n_3035;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_3333;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_2811;
wire n_1496;
wire n_3348;
wire n_1125;
wire n_2547;
wire n_3014;
wire n_1812;
wire n_2501;
wire n_3079;
wire n_1915;
wire n_1109;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_3308;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_1533;
wire n_2224;
wire n_3368;
wire n_2924;
wire n_2484;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_3329;
wire n_2994;
wire n_1067;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_3135;
wire n_2003;
wire n_1457;
wire n_2692;
wire n_3148;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_2264;
wire n_2754;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_2012;
wire n_1291;
wire n_3381;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_3278;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_2965;
wire n_3217;
wire n_1703;
wire n_3312;
wire n_1352;
wire n_2926;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_3046;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_3249;
wire n_3211;
wire n_3285;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_2103;
wire n_2160;
wire n_3337;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_3074;
wire n_3204;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_2363;
wire n_2430;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_1235;
wire n_1115;
wire n_2433;
wire n_3293;
wire n_3129;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_2977;
wire n_2601;
wire n_3043;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_1334;
wire n_1907;
wire n_2686;
wire n_2528;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_1985;
wire n_3055;
wire n_1898;
wire n_2107;
wire n_3294;
wire n_3219;
wire n_3315;
wire n_2906;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_2817;
wire n_3172;
wire n_3139;
wire n_2773;
wire n_3239;
wire n_3292;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_3365;
wire n_1452;
wire n_2687;
wire n_3023;
wire n_1120;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_2850;
wire n_1683;
wire n_1817;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_2654;
wire n_997;
wire n_3104;
wire n_3169;
wire n_3151;
wire n_3131;
wire n_2078;
wire n_1409;
wire n_1326;
wire n_3070;
wire n_3284;
wire n_3176;
wire n_2884;
wire n_1268;
wire n_2996;
wire n_2819;
wire n_3126;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_1718;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_1922;
wire n_2966;
wire n_1376;
wire n_2326;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_2950;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_3140;
wire n_3170;
wire n_2104;
wire n_2748;
wire n_3311;
wire n_2057;
wire n_3272;
wire n_3011;
wire n_1772;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_3345;
wire n_1425;
wire n_1901;
wire n_3069;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_2889;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_3313;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_2939;
wire n_1745;
wire n_2735;
wire n_2497;
wire n_2006;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_1618;
wire n_2260;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_2014;
wire n_3056;
wire n_1221;
wire n_2345;
wire n_2986;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2726;
wire n_2774;
wire n_3295;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_2382;
wire n_1707;
wire n_3062;
wire n_3161;
wire n_2317;
wire n_3289;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_3017;
wire n_2476;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_2984;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_3364;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_1873;
wire n_1411;
wire n_3201;
wire n_3054;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_3344;
wire n_2194;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_3302;
wire n_3235;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_3102;
wire n_3122;
wire n_1648;
wire n_1536;
wire n_3050;
wire n_3265;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_2957;
wire n_1769;
wire n_1210;
wire n_2964;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_3314;
wire n_2360;
wire n_3254;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_2442;
wire n_3309;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_2018;
wire n_3260;
wire n_1555;
wire n_3117;
wire n_2834;
wire n_3245;
wire n_3357;
wire n_2531;
wire n_1589;
wire n_2961;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_1858;
wire n_3351;
wire n_1619;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_2883;
wire n_3115;
wire n_3352;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_3063;
wire n_2912;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_3251;
wire n_1910;
wire n_1298;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_2809;
wire n_2050;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_3118;
wire n_3227;
wire n_3300;
wire n_2321;
wire n_1226;
wire n_1277;
wire n_2591;
wire n_2146;
wire n_3384;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_3336;
wire n_2940;
wire n_1546;
wire n_2612;
wire n_1495;
wire n_1337;
wire n_1515;
wire n_2841;
wire n_3165;
wire n_1627;
wire n_2918;
wire n_3232;
wire n_3322;
wire n_1245;
wire n_2427;
wire n_2505;
wire n_2438;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_3250;
wire n_1739;
wire n_3181;
wire n_2958;
wire n_2278;
wire n_3114;
wire n_2594;
wire n_3125;
wire n_3234;
wire n_2394;
wire n_1914;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3004;
wire n_3323;
wire n_2569;
wire n_3112;
wire n_2349;
wire n_1103;
wire n_3132;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_3024;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_3238;
wire n_3210;
wire n_3175;
wire n_2036;
wire n_1325;
wire n_3267;
wire n_1595;
wire n_2161;
wire n_2404;
wire n_2083;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_3266;
wire n_2485;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_2210;
wire n_3247;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_3091;
wire n_2695;
wire n_1764;
wire n_2892;
wire n_3057;
wire n_3194;
wire n_3066;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_3347;
wire n_2004;
wire n_3216;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_1996;
wire n_1505;
wire n_1181;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_1340;
wire n_2274;
wire n_2972;
wire n_1558;
wire n_3225;
wire n_3321;
wire n_2166;
wire n_2938;
wire n_3212;
wire n_3319;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_3152;
wire n_3335;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2689;
wire n_2920;
wire n_3259;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_2991;
wire n_3383;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_2975;
wire n_2599;
wire n_2704;
wire n_2839;
wire n_3338;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_3360;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_3159;
wire n_2728;
wire n_2268;

INVx1_ASAP7_75t_L g993 ( 
.A(n_17),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_701),
.Y(n_994)
);

CKINVDCx16_ASAP7_75t_R g995 ( 
.A(n_135),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_788),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_928),
.Y(n_997)
);

CKINVDCx16_ASAP7_75t_R g998 ( 
.A(n_754),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_871),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_288),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_873),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_940),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_840),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_58),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_852),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_962),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_936),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_960),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_710),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_850),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_701),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_203),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_556),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_168),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_120),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_370),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_257),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_524),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_823),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_649),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_865),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_844),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_379),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_943),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_389),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_265),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_900),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_201),
.Y(n_1028)
);

BUFx10_ASAP7_75t_L g1029 ( 
.A(n_112),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_650),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_713),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_426),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_166),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_659),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_912),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_406),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_944),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_63),
.Y(n_1038)
);

CKINVDCx20_ASAP7_75t_R g1039 ( 
.A(n_129),
.Y(n_1039)
);

INVx4_ASAP7_75t_R g1040 ( 
.A(n_479),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_951),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_51),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_947),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_35),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_924),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_828),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_686),
.Y(n_1047)
);

CKINVDCx20_ASAP7_75t_R g1048 ( 
.A(n_927),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_918),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_740),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_806),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_552),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_734),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_306),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_141),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_80),
.Y(n_1056)
);

CKINVDCx20_ASAP7_75t_R g1057 ( 
.A(n_898),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_438),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_600),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_203),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_535),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_892),
.Y(n_1062)
);

INVx1_ASAP7_75t_SL g1063 ( 
.A(n_602),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_620),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_910),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_895),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_942),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_484),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_907),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_23),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_982),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_917),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_122),
.Y(n_1073)
);

CKINVDCx16_ASAP7_75t_R g1074 ( 
.A(n_948),
.Y(n_1074)
);

CKINVDCx16_ASAP7_75t_R g1075 ( 
.A(n_970),
.Y(n_1075)
);

INVx1_ASAP7_75t_SL g1076 ( 
.A(n_645),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_930),
.Y(n_1077)
);

BUFx5_ASAP7_75t_L g1078 ( 
.A(n_42),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_151),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_144),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_595),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_409),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_839),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_886),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_909),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_292),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_573),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_684),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_453),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_926),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_914),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_263),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_8),
.Y(n_1093)
);

BUFx10_ASAP7_75t_L g1094 ( 
.A(n_916),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_92),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_699),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_643),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_191),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_915),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_172),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_689),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_676),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_211),
.Y(n_1103)
);

BUFx10_ASAP7_75t_L g1104 ( 
.A(n_81),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_937),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_837),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_152),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_436),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_507),
.Y(n_1109)
);

CKINVDCx20_ASAP7_75t_R g1110 ( 
.A(n_487),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_956),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_237),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_964),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_966),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_135),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_959),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_266),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_988),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_699),
.Y(n_1119)
);

INVx1_ASAP7_75t_SL g1120 ( 
.A(n_279),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_466),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_679),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_653),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_697),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_706),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_722),
.Y(n_1126)
);

BUFx5_ASAP7_75t_L g1127 ( 
.A(n_737),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_794),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_43),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_91),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_935),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_429),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_961),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_317),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_680),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_132),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_695),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_314),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_796),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_450),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_138),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_320),
.Y(n_1142)
);

CKINVDCx20_ASAP7_75t_R g1143 ( 
.A(n_160),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_238),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_460),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_696),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_301),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_832),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_219),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_235),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_461),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_698),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_504),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_449),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_688),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_983),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_925),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_495),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_0),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_913),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_170),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_290),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_812),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_673),
.Y(n_1164)
);

CKINVDCx20_ASAP7_75t_R g1165 ( 
.A(n_934),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_370),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_922),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_617),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_485),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_318),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_954),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_901),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_938),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_887),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_423),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_463),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_183),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_953),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_905),
.Y(n_1179)
);

BUFx8_ASAP7_75t_SL g1180 ( 
.A(n_511),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_190),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_58),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_509),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_249),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_415),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_853),
.Y(n_1186)
);

INVxp67_ASAP7_75t_L g1187 ( 
.A(n_921),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_166),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_893),
.Y(n_1189)
);

CKINVDCx16_ASAP7_75t_R g1190 ( 
.A(n_902),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_933),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_771),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_678),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_633),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_702),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_950),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_499),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_919),
.Y(n_1198)
);

BUFx10_ASAP7_75t_L g1199 ( 
.A(n_680),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_677),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_248),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_920),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_322),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_574),
.Y(n_1204)
);

CKINVDCx20_ASAP7_75t_R g1205 ( 
.A(n_785),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_949),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_764),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_353),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_894),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_474),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_86),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_387),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_449),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_305),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_134),
.Y(n_1215)
);

CKINVDCx16_ASAP7_75t_R g1216 ( 
.A(n_890),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_383),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_360),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_958),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_123),
.Y(n_1220)
);

CKINVDCx16_ASAP7_75t_R g1221 ( 
.A(n_691),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_719),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_609),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_145),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_515),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_581),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_770),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_285),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_911),
.Y(n_1229)
);

INVxp67_ASAP7_75t_L g1230 ( 
.A(n_904),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_711),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_651),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_478),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_228),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_412),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_24),
.Y(n_1236)
);

HB1xp67_ASAP7_75t_L g1237 ( 
.A(n_75),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_897),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_827),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_976),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_693),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_277),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_923),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_210),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_675),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_550),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_331),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_276),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_632),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_600),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_702),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_12),
.Y(n_1252)
);

CKINVDCx16_ASAP7_75t_R g1253 ( 
.A(n_646),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_456),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_602),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_128),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_931),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_316),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_700),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_681),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_368),
.Y(n_1261)
);

INVxp67_ASAP7_75t_SL g1262 ( 
.A(n_442),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_26),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_687),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_525),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_75),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_831),
.Y(n_1267)
);

INVx1_ASAP7_75t_SL g1268 ( 
.A(n_533),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_625),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_199),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_582),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_683),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_929),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_548),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_685),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_29),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_682),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_118),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_903),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_946),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_808),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_316),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_782),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_343),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_420),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_617),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_773),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_896),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_94),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_704),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_874),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_123),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_690),
.Y(n_1293)
);

INVx1_ASAP7_75t_SL g1294 ( 
.A(n_939),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_43),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_694),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_855),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_987),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_703),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_305),
.Y(n_1300)
);

CKINVDCx16_ASAP7_75t_R g1301 ( 
.A(n_989),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_198),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_217),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_22),
.Y(n_1304)
);

BUFx2_ASAP7_75t_L g1305 ( 
.A(n_818),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_347),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_932),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_194),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_42),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_538),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_275),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_804),
.Y(n_1312)
);

BUFx8_ASAP7_75t_SL g1313 ( 
.A(n_550),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_92),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_486),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_952),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_102),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_168),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_349),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_240),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_292),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_908),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_301),
.Y(n_1323)
);

BUFx10_ASAP7_75t_L g1324 ( 
.A(n_906),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_963),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_231),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_665),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_758),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_691),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_538),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_158),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_18),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_242),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_692),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_38),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_672),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_14),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_97),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_278),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_945),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_330),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_124),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_60),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_700),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_655),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_955),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_941),
.Y(n_1347)
);

CKINVDCx20_ASAP7_75t_R g1348 ( 
.A(n_57),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_825),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_574),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_371),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_957),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_842),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_229),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_47),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_377),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_593),
.Y(n_1357)
);

CKINVDCx20_ASAP7_75t_R g1358 ( 
.A(n_82),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_250),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_530),
.Y(n_1360)
);

BUFx5_ASAP7_75t_L g1361 ( 
.A(n_591),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_899),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_426),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1078),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1078),
.Y(n_1365)
);

INVxp33_ASAP7_75t_L g1366 ( 
.A(n_1237),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1078),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1078),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1078),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1361),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1361),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1361),
.Y(n_1372)
);

INVxp67_ASAP7_75t_L g1373 ( 
.A(n_1089),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1361),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1180),
.Y(n_1375)
);

INVxp33_ASAP7_75t_SL g1376 ( 
.A(n_1327),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1361),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1318),
.Y(n_1378)
);

CKINVDCx16_ASAP7_75t_R g1379 ( 
.A(n_995),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1318),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1052),
.Y(n_1381)
);

INVxp67_ASAP7_75t_SL g1382 ( 
.A(n_1305),
.Y(n_1382)
);

INVxp67_ASAP7_75t_SL g1383 ( 
.A(n_1027),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1052),
.Y(n_1384)
);

INVxp33_ASAP7_75t_L g1385 ( 
.A(n_1313),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1052),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1070),
.Y(n_1387)
);

INVxp67_ASAP7_75t_L g1388 ( 
.A(n_1121),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1221),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_996),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1070),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_1048),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_997),
.Y(n_1393)
);

INVxp33_ASAP7_75t_SL g1394 ( 
.A(n_1000),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1070),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1101),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1101),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1094),
.Y(n_1398)
);

CKINVDCx16_ASAP7_75t_R g1399 ( 
.A(n_1253),
.Y(n_1399)
);

INVxp67_ASAP7_75t_SL g1400 ( 
.A(n_1041),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1101),
.Y(n_1401)
);

CKINVDCx14_ASAP7_75t_R g1402 ( 
.A(n_1094),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_1057),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1245),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_1067),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1156),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1245),
.Y(n_1407)
);

INVxp67_ASAP7_75t_SL g1408 ( 
.A(n_1125),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1245),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_1165),
.Y(n_1410)
);

INVxp33_ASAP7_75t_SL g1411 ( 
.A(n_1004),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1276),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1276),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_1029),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_SL g1415 ( 
.A(n_1029),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_999),
.Y(n_1416)
);

INVxp67_ASAP7_75t_SL g1417 ( 
.A(n_1297),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1276),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1023),
.Y(n_1419)
);

INVxp33_ASAP7_75t_L g1420 ( 
.A(n_993),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1032),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_1205),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1219),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1055),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1001),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1235),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1002),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1249),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_994),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1017),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1018),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1036),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1390),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_1392),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1395),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1376),
.A2(n_1382),
.B1(n_1373),
.B2(n_1366),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1407),
.Y(n_1437)
);

BUFx6f_ASAP7_75t_L g1438 ( 
.A(n_1418),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_SL g1439 ( 
.A1(n_1402),
.A2(n_1098),
.B1(n_1110),
.B2(n_1039),
.Y(n_1439)
);

INVx5_ASAP7_75t_L g1440 ( 
.A(n_1398),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1381),
.Y(n_1441)
);

INVx3_ASAP7_75t_L g1442 ( 
.A(n_1384),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1386),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1387),
.Y(n_1444)
);

BUFx6f_ASAP7_75t_L g1445 ( 
.A(n_1391),
.Y(n_1445)
);

OAI22x1_ASAP7_75t_L g1446 ( 
.A1(n_1414),
.A2(n_1076),
.B1(n_1112),
.B2(n_1063),
.Y(n_1446)
);

INVx2_ASAP7_75t_SL g1447 ( 
.A(n_1419),
.Y(n_1447)
);

AOI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1379),
.A2(n_1074),
.B1(n_1075),
.B2(n_998),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1393),
.Y(n_1449)
);

XNOR2xp5_ASAP7_75t_L g1450 ( 
.A(n_1403),
.B(n_1119),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1416),
.B(n_1037),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1396),
.Y(n_1452)
);

AOI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1399),
.A2(n_1216),
.B1(n_1301),
.B2(n_1190),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1397),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1401),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1394),
.A2(n_1316),
.B1(n_1322),
.B2(n_1238),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1404),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1409),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1389),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1415),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1383),
.B(n_1324),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1412),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1413),
.Y(n_1463)
);

BUFx12f_ASAP7_75t_L g1464 ( 
.A(n_1375),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1364),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1429),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1400),
.B(n_1187),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1365),
.Y(n_1468)
);

INVx5_ASAP7_75t_L g1469 ( 
.A(n_1415),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1367),
.Y(n_1470)
);

BUFx12f_ASAP7_75t_L g1471 ( 
.A(n_1425),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1368),
.Y(n_1472)
);

INVx5_ASAP7_75t_L g1473 ( 
.A(n_1411),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1369),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1370),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1427),
.B(n_1046),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1430),
.Y(n_1477)
);

OA21x2_ASAP7_75t_L g1478 ( 
.A1(n_1371),
.A2(n_1230),
.B(n_1019),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1420),
.A2(n_1087),
.B1(n_1012),
.B2(n_1014),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1421),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1385),
.B(n_1324),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1433),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_1461),
.Y(n_1483)
);

INVxp33_ASAP7_75t_SL g1484 ( 
.A(n_1450),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1466),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1449),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_R g1487 ( 
.A(n_1434),
.B(n_1405),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1471),
.Y(n_1488)
);

AND3x1_ASAP7_75t_L g1489 ( 
.A(n_1448),
.B(n_1224),
.C(n_1146),
.Y(n_1489)
);

CKINVDCx20_ASAP7_75t_R g1490 ( 
.A(n_1456),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1467),
.B(n_1408),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1464),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1473),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1473),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1469),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1469),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1451),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1476),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1459),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1436),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1440),
.Y(n_1501)
);

CKINVDCx20_ASAP7_75t_R g1502 ( 
.A(n_1453),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1440),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_1439),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_R g1505 ( 
.A(n_1472),
.B(n_1406),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1477),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1460),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1438),
.Y(n_1508)
);

BUFx2_ASAP7_75t_L g1509 ( 
.A(n_1446),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1445),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1475),
.B(n_1417),
.Y(n_1511)
);

NOR2xp67_ASAP7_75t_L g1512 ( 
.A(n_1480),
.B(n_1388),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1479),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1481),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1447),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1445),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1457),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1465),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1468),
.Y(n_1519)
);

NOR2xp67_ASAP7_75t_L g1520 ( 
.A(n_1441),
.B(n_1388),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1470),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1474),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1443),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1444),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1455),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1454),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1458),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1462),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_1442),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1463),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1452),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1435),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_R g1533 ( 
.A(n_1437),
.B(n_1410),
.Y(n_1533)
);

NAND2xp33_ASAP7_75t_R g1534 ( 
.A(n_1478),
.B(n_1013),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1433),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1433),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1433),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1433),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1438),
.Y(n_1539)
);

CKINVDCx20_ASAP7_75t_R g1540 ( 
.A(n_1434),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1433),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1459),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1466),
.Y(n_1543)
);

BUFx6f_ASAP7_75t_L g1544 ( 
.A(n_1438),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1476),
.B(n_1372),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1433),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1433),
.Y(n_1547)
);

CKINVDCx20_ASAP7_75t_R g1548 ( 
.A(n_1434),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1438),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1438),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1476),
.B(n_1374),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1433),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1524),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1545),
.A2(n_1114),
.B1(n_1192),
.B2(n_1065),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1517),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1551),
.A2(n_1291),
.B1(n_1347),
.B2(n_1283),
.Y(n_1556)
);

INVx3_ASAP7_75t_L g1557 ( 
.A(n_1544),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_SL g1558 ( 
.A1(n_1490),
.A2(n_1504),
.B1(n_1502),
.B2(n_1500),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1523),
.Y(n_1559)
);

INVx4_ASAP7_75t_L g1560 ( 
.A(n_1544),
.Y(n_1560)
);

INVx4_ASAP7_75t_L g1561 ( 
.A(n_1544),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1498),
.B(n_1497),
.Y(n_1562)
);

OAI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1513),
.A2(n_1423),
.B1(n_1422),
.B2(n_1262),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1518),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1519),
.Y(n_1565)
);

OAI221xp5_ASAP7_75t_L g1566 ( 
.A1(n_1511),
.A2(n_1236),
.B1(n_1042),
.B2(n_1056),
.C(n_1054),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1483),
.B(n_1294),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1526),
.B(n_1353),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1482),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1491),
.A2(n_1021),
.B1(n_1022),
.B2(n_1006),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1521),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1522),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1515),
.B(n_1003),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1529),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1527),
.B(n_1120),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1508),
.Y(n_1576)
);

INVx4_ASAP7_75t_L g1577 ( 
.A(n_1510),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1531),
.B(n_1377),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1516),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1485),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_1486),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1510),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_SL g1583 ( 
.A(n_1528),
.B(n_1005),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1530),
.B(n_1024),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1532),
.B(n_1007),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1514),
.B(n_1135),
.Y(n_1586)
);

INVx3_ASAP7_75t_L g1587 ( 
.A(n_1539),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1509),
.A2(n_1031),
.B1(n_1071),
.B2(n_1053),
.Y(n_1588)
);

NAND2xp33_ASAP7_75t_L g1589 ( 
.A(n_1510),
.B(n_1008),
.Y(n_1589)
);

NAND2xp33_ASAP7_75t_SL g1590 ( 
.A(n_1505),
.B(n_1143),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1499),
.B(n_1268),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1506),
.Y(n_1592)
);

INVxp67_ASAP7_75t_SL g1593 ( 
.A(n_1525),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1549),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1512),
.B(n_1072),
.Y(n_1595)
);

INVx3_ASAP7_75t_L g1596 ( 
.A(n_1550),
.Y(n_1596)
);

INVxp33_ASAP7_75t_L g1597 ( 
.A(n_1542),
.Y(n_1597)
);

BUFx6f_ASAP7_75t_SL g1598 ( 
.A(n_1543),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1525),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1520),
.Y(n_1600)
);

AND2x4_ASAP7_75t_L g1601 ( 
.A(n_1489),
.B(n_1431),
.Y(n_1601)
);

INVxp33_ASAP7_75t_L g1602 ( 
.A(n_1487),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1533),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1535),
.B(n_1424),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1493),
.B(n_1077),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1501),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1503),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1494),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1495),
.Y(n_1609)
);

NAND2xp33_ASAP7_75t_SL g1610 ( 
.A(n_1534),
.B(n_1176),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1536),
.B(n_1426),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1496),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1537),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1540),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1538),
.B(n_1009),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1541),
.Y(n_1616)
);

OR2x2_ASAP7_75t_SL g1617 ( 
.A(n_1484),
.B(n_1011),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1507),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1548),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1552),
.B(n_1084),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_L g1621 ( 
.A(n_1546),
.B(n_1319),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1547),
.A2(n_1105),
.B1(n_1157),
.B2(n_1085),
.Y(n_1622)
);

BUFx2_ASAP7_75t_L g1623 ( 
.A(n_1488),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1492),
.B(n_1432),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_1482),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1545),
.A2(n_1173),
.B1(n_1179),
.B2(n_1178),
.Y(n_1626)
);

NAND3xp33_ASAP7_75t_L g1627 ( 
.A(n_1513),
.B(n_1428),
.C(n_1016),
.Y(n_1627)
);

BUFx6f_ASAP7_75t_L g1628 ( 
.A(n_1544),
.Y(n_1628)
);

BUFx6f_ASAP7_75t_L g1629 ( 
.A(n_1544),
.Y(n_1629)
);

AND2x6_ASAP7_75t_L g1630 ( 
.A(n_1491),
.B(n_1196),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1508),
.B(n_1378),
.Y(n_1631)
);

INVx4_ASAP7_75t_L g1632 ( 
.A(n_1524),
.Y(n_1632)
);

BUFx6f_ASAP7_75t_L g1633 ( 
.A(n_1544),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1498),
.B(n_1010),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_SL g1635 ( 
.A(n_1482),
.B(n_1358),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1498),
.B(n_1015),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1517),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1523),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1483),
.B(n_1380),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1523),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1524),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1499),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1523),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1483),
.B(n_1104),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1499),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1498),
.B(n_1020),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1523),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1523),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1523),
.Y(n_1649)
);

OAI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1500),
.A2(n_1340),
.B1(n_1222),
.B2(n_1273),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1545),
.A2(n_1267),
.B1(n_1287),
.B2(n_1280),
.Y(n_1651)
);

INVx4_ASAP7_75t_L g1652 ( 
.A(n_1524),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1523),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_R g1654 ( 
.A(n_1482),
.B(n_1035),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1523),
.Y(n_1655)
);

BUFx3_ASAP7_75t_L g1656 ( 
.A(n_1524),
.Y(n_1656)
);

AO21x2_ASAP7_75t_L g1657 ( 
.A1(n_1545),
.A2(n_1362),
.B(n_1307),
.Y(n_1657)
);

BUFx6f_ASAP7_75t_L g1658 ( 
.A(n_1544),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1524),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1498),
.B(n_1043),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1498),
.B(n_1352),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1483),
.B(n_1104),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1498),
.B(n_1045),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1523),
.Y(n_1664)
);

BUFx6f_ASAP7_75t_L g1665 ( 
.A(n_1544),
.Y(n_1665)
);

BUFx4f_ASAP7_75t_L g1666 ( 
.A(n_1544),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1523),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1555),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1628),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1568),
.B(n_1660),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1575),
.B(n_1199),
.Y(n_1671)
);

INVx8_ASAP7_75t_L g1672 ( 
.A(n_1630),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1663),
.B(n_1049),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1636),
.B(n_1050),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_SL g1675 ( 
.A(n_1562),
.B(n_1051),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1610),
.A2(n_1066),
.B1(n_1069),
.B2(n_1062),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1559),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1637),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1586),
.B(n_1199),
.Y(n_1679)
);

BUFx3_ASAP7_75t_L g1680 ( 
.A(n_1553),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1621),
.B(n_1210),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1646),
.B(n_1083),
.Y(n_1682)
);

O2A1O1Ixp5_ASAP7_75t_L g1683 ( 
.A1(n_1638),
.A2(n_1246),
.B(n_1277),
.C(n_1144),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1597),
.B(n_1234),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1640),
.Y(n_1685)
);

INVxp33_ASAP7_75t_L g1686 ( 
.A(n_1591),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1578),
.B(n_1643),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1647),
.B(n_1090),
.Y(n_1688)
);

OR2x6_ASAP7_75t_L g1689 ( 
.A(n_1641),
.B(n_1044),
.Y(n_1689)
);

O2A1O1Ixp5_ASAP7_75t_L g1690 ( 
.A1(n_1648),
.A2(n_1317),
.B(n_1335),
.C(n_1302),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1611),
.B(n_1266),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1649),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1653),
.B(n_1091),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1655),
.B(n_1099),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1570),
.A2(n_1333),
.B1(n_1337),
.B2(n_1292),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1628),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1620),
.B(n_1345),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1602),
.B(n_1348),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1664),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1667),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1603),
.B(n_1604),
.Y(n_1701)
);

INVx3_ASAP7_75t_L g1702 ( 
.A(n_1629),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1564),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_SL g1704 ( 
.A(n_1569),
.B(n_1106),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1642),
.B(n_1111),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1645),
.B(n_1350),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1626),
.A2(n_1127),
.B1(n_1279),
.B2(n_1343),
.Y(n_1707)
);

AND2x6_ASAP7_75t_SL g1708 ( 
.A(n_1613),
.B(n_1351),
.Y(n_1708)
);

INVx3_ASAP7_75t_L g1709 ( 
.A(n_1629),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1619),
.B(n_1354),
.Y(n_1710)
);

OR2x6_ASAP7_75t_L g1711 ( 
.A(n_1656),
.B(n_1079),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_SL g1712 ( 
.A(n_1584),
.B(n_1113),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1565),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1639),
.B(n_1600),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1634),
.B(n_1025),
.Y(n_1715)
);

AOI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1630),
.A2(n_1118),
.B1(n_1126),
.B2(n_1116),
.Y(n_1716)
);

INVx2_ASAP7_75t_SL g1717 ( 
.A(n_1666),
.Y(n_1717)
);

INVx2_ASAP7_75t_SL g1718 ( 
.A(n_1633),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1571),
.B(n_1128),
.Y(n_1719)
);

OAI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1651),
.A2(n_1133),
.B1(n_1139),
.B2(n_1131),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1572),
.B(n_1148),
.Y(n_1721)
);

INVx2_ASAP7_75t_SL g1722 ( 
.A(n_1633),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1631),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_SL g1724 ( 
.A(n_1581),
.B(n_1625),
.Y(n_1724)
);

NAND3xp33_ASAP7_75t_L g1725 ( 
.A(n_1622),
.B(n_1028),
.C(n_1026),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1579),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1630),
.B(n_1160),
.Y(n_1727)
);

INVx2_ASAP7_75t_SL g1728 ( 
.A(n_1658),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_SL g1729 ( 
.A(n_1635),
.B(n_1163),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1627),
.B(n_1654),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1661),
.B(n_1030),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1595),
.B(n_1644),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1662),
.B(n_1167),
.Y(n_1733)
);

O2A1O1Ixp5_ASAP7_75t_L g1734 ( 
.A1(n_1567),
.A2(n_1359),
.B(n_1081),
.C(n_1092),
.Y(n_1734)
);

BUFx3_ASAP7_75t_L g1735 ( 
.A(n_1659),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1563),
.B(n_1033),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1594),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1618),
.B(n_1171),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_SL g1739 ( 
.A(n_1632),
.B(n_1172),
.Y(n_1739)
);

INVxp67_ASAP7_75t_L g1740 ( 
.A(n_1605),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1624),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1616),
.B(n_1583),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_SL g1743 ( 
.A(n_1623),
.B(n_1174),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1652),
.B(n_1186),
.Y(n_1744)
);

AND2x2_ASAP7_75t_SL g1745 ( 
.A(n_1606),
.B(n_1588),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1657),
.A2(n_1189),
.B1(n_1198),
.B2(n_1191),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1615),
.B(n_1034),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1582),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1554),
.B(n_1202),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1585),
.B(n_1038),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1556),
.B(n_1206),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1580),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1593),
.B(n_1577),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1592),
.Y(n_1754)
);

BUFx2_ASAP7_75t_L g1755 ( 
.A(n_1614),
.Y(n_1755)
);

INVxp67_ASAP7_75t_SL g1756 ( 
.A(n_1658),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1650),
.B(n_1207),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1574),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1573),
.B(n_1047),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1601),
.A2(n_1127),
.B1(n_1279),
.B2(n_1355),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1599),
.B(n_1058),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1576),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1587),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1596),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1558),
.B(n_1059),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1557),
.B(n_1209),
.Y(n_1766)
);

BUFx8_ASAP7_75t_L g1767 ( 
.A(n_1598),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1665),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1665),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1560),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_SL g1771 ( 
.A(n_1590),
.B(n_1227),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1561),
.B(n_1229),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1589),
.A2(n_1279),
.B(n_1239),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1608),
.A2(n_1231),
.B1(n_1243),
.B2(n_1240),
.Y(n_1774)
);

INVx5_ASAP7_75t_L g1775 ( 
.A(n_1606),
.Y(n_1775)
);

INVx2_ASAP7_75t_SL g1776 ( 
.A(n_1609),
.Y(n_1776)
);

NOR3xp33_ASAP7_75t_L g1777 ( 
.A(n_1566),
.B(n_1061),
.C(n_1060),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1617),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1612),
.B(n_1064),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1607),
.B(n_1257),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1568),
.B(n_1281),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_SL g1782 ( 
.A(n_1562),
.B(n_1288),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1568),
.B(n_1290),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1610),
.A2(n_1127),
.B1(n_1093),
.B2(n_1095),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_L g1785 ( 
.A(n_1562),
.B(n_1068),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1610),
.A2(n_1127),
.B1(n_1096),
.B2(n_1103),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1555),
.Y(n_1787)
);

AOI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1610),
.A2(n_1127),
.B1(n_1336),
.B2(n_1334),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1562),
.B(n_1073),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1562),
.B(n_1339),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1568),
.B(n_1298),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1568),
.B(n_1312),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1555),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_SL g1794 ( 
.A(n_1562),
.B(n_1325),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1555),
.Y(n_1795)
);

AND2x6_ASAP7_75t_SL g1796 ( 
.A(n_1621),
.B(n_1356),
.Y(n_1796)
);

AND2x6_ASAP7_75t_SL g1797 ( 
.A(n_1621),
.B(n_1082),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1562),
.B(n_1080),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1555),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1555),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1559),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1568),
.B(n_1328),
.Y(n_1802)
);

INVxp67_ASAP7_75t_SL g1803 ( 
.A(n_1628),
.Y(n_1803)
);

BUFx3_ASAP7_75t_L g1804 ( 
.A(n_1553),
.Y(n_1804)
);

INVx2_ASAP7_75t_SL g1805 ( 
.A(n_1645),
.Y(n_1805)
);

BUFx3_ASAP7_75t_L g1806 ( 
.A(n_1553),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1568),
.B(n_1346),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1562),
.B(n_1349),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1562),
.B(n_1086),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1559),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1555),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1645),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1559),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_L g1814 ( 
.A(n_1562),
.B(n_1088),
.Y(n_1814)
);

BUFx6f_ASAP7_75t_L g1815 ( 
.A(n_1628),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1555),
.Y(n_1816)
);

HB1xp67_ASAP7_75t_L g1817 ( 
.A(n_1645),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1562),
.B(n_1097),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1562),
.B(n_1100),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1559),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1610),
.A2(n_1330),
.B1(n_1342),
.B2(n_1326),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1562),
.B(n_1102),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1555),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1562),
.B(n_1331),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1568),
.B(n_1107),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1555),
.Y(n_1826)
);

AOI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1610),
.A2(n_1129),
.B1(n_1134),
.B2(n_1124),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1775),
.B(n_1145),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1670),
.B(n_1108),
.Y(n_1829)
);

AOI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1732),
.A2(n_1687),
.B(n_1673),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1740),
.B(n_1109),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_SL g1832 ( 
.A(n_1724),
.B(n_1115),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1685),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1753),
.A2(n_1164),
.B(n_1151),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1686),
.B(n_1117),
.Y(n_1835)
);

CKINVDCx10_ASAP7_75t_R g1836 ( 
.A(n_1689),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1785),
.B(n_1122),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1681),
.A2(n_1123),
.B1(n_1132),
.B2(n_1130),
.Y(n_1838)
);

OAI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1714),
.A2(n_1136),
.B1(n_1138),
.B2(n_1137),
.Y(n_1839)
);

OAI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1677),
.A2(n_1188),
.B(n_1181),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1674),
.A2(n_1203),
.B(n_1193),
.Y(n_1841)
);

OAI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1692),
.A2(n_1217),
.B(n_1204),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1682),
.A2(n_1220),
.B(n_1218),
.Y(n_1843)
);

OAI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1699),
.A2(n_1225),
.B(n_1223),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1815),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1781),
.A2(n_1248),
.B(n_1228),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1783),
.A2(n_1254),
.B(n_1251),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1789),
.B(n_1140),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1798),
.B(n_1141),
.Y(n_1849)
);

BUFx6f_ASAP7_75t_L g1850 ( 
.A(n_1815),
.Y(n_1850)
);

AOI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1791),
.A2(n_1270),
.B(n_1258),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1801),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1700),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1792),
.A2(n_1284),
.B(n_1282),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_SL g1855 ( 
.A(n_1742),
.B(n_1142),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1802),
.A2(n_1286),
.B(n_1285),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1697),
.B(n_1147),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1691),
.B(n_1149),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1809),
.B(n_1150),
.Y(n_1859)
);

AOI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1807),
.A2(n_1293),
.B(n_1289),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1810),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_SL g1862 ( 
.A(n_1701),
.B(n_1152),
.Y(n_1862)
);

AOI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1772),
.A2(n_1733),
.B(n_1693),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1813),
.Y(n_1864)
);

AO21x1_ASAP7_75t_L g1865 ( 
.A1(n_1715),
.A2(n_1304),
.B(n_1299),
.Y(n_1865)
);

O2A1O1Ixp33_ASAP7_75t_L g1866 ( 
.A1(n_1825),
.A2(n_1306),
.B(n_1310),
.C(n_1309),
.Y(n_1866)
);

CKINVDCx20_ASAP7_75t_R g1867 ( 
.A(n_1680),
.Y(n_1867)
);

AOI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1688),
.A2(n_1315),
.B(n_1314),
.Y(n_1868)
);

INVx2_ASAP7_75t_SL g1869 ( 
.A(n_1805),
.Y(n_1869)
);

A2O1A1Ixp33_ASAP7_75t_L g1870 ( 
.A1(n_1736),
.A2(n_1320),
.B(n_1153),
.C(n_1155),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1814),
.B(n_1154),
.Y(n_1871)
);

OAI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1820),
.A2(n_1159),
.B(n_1158),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1679),
.B(n_1161),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1671),
.B(n_1162),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1703),
.B(n_1713),
.Y(n_1875)
);

BUFx3_ASAP7_75t_L g1876 ( 
.A(n_1775),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1752),
.Y(n_1877)
);

INVx1_ASAP7_75t_SL g1878 ( 
.A(n_1812),
.Y(n_1878)
);

AOI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1694),
.A2(n_707),
.B(n_705),
.Y(n_1879)
);

BUFx4f_ASAP7_75t_L g1880 ( 
.A(n_1745),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1731),
.B(n_1166),
.Y(n_1881)
);

O2A1O1Ixp33_ASAP7_75t_L g1882 ( 
.A1(n_1778),
.A2(n_1040),
.B(n_1169),
.C(n_1168),
.Y(n_1882)
);

O2A1O1Ixp33_ASAP7_75t_SL g1883 ( 
.A1(n_1757),
.A2(n_709),
.B(n_712),
.C(n_708),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1668),
.Y(n_1884)
);

AOI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1675),
.A2(n_715),
.B(n_714),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1750),
.B(n_1170),
.Y(n_1886)
);

AOI21xp5_ASAP7_75t_L g1887 ( 
.A1(n_1782),
.A2(n_1808),
.B(n_1794),
.Y(n_1887)
);

AOI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1712),
.A2(n_717),
.B(n_716),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1790),
.B(n_1175),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1730),
.A2(n_720),
.B(n_718),
.Y(n_1890)
);

AOI21x1_ASAP7_75t_L g1891 ( 
.A1(n_1748),
.A2(n_1721),
.B(n_1719),
.Y(n_1891)
);

NOR3xp33_ASAP7_75t_L g1892 ( 
.A(n_1695),
.B(n_1182),
.C(n_1177),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1766),
.A2(n_723),
.B(n_721),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1698),
.B(n_1183),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1749),
.A2(n_725),
.B(n_724),
.Y(n_1895)
);

INVx2_ASAP7_75t_SL g1896 ( 
.A(n_1817),
.Y(n_1896)
);

HB1xp67_ASAP7_75t_L g1897 ( 
.A(n_1775),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1678),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1824),
.B(n_1184),
.Y(n_1899)
);

OAI21xp5_ASAP7_75t_L g1900 ( 
.A1(n_1784),
.A2(n_1194),
.B(n_1185),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1747),
.B(n_1195),
.Y(n_1901)
);

OAI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1786),
.A2(n_1788),
.B(n_1690),
.Y(n_1902)
);

AOI21x1_ASAP7_75t_L g1903 ( 
.A1(n_1738),
.A2(n_727),
.B(n_726),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1787),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1754),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1759),
.B(n_1197),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1751),
.A2(n_729),
.B(n_728),
.Y(n_1907)
);

AOI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1793),
.A2(n_731),
.B(n_730),
.Y(n_1908)
);

A2O1A1Ixp33_ASAP7_75t_L g1909 ( 
.A1(n_1779),
.A2(n_1201),
.B(n_1208),
.C(n_1200),
.Y(n_1909)
);

AOI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1795),
.A2(n_733),
.B(n_732),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_L g1911 ( 
.A(n_1684),
.B(n_1211),
.Y(n_1911)
);

AOI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1799),
.A2(n_1826),
.B(n_1823),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1800),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1811),
.B(n_1212),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1816),
.B(n_1213),
.Y(n_1915)
);

OAI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1683),
.A2(n_1215),
.B(n_1214),
.Y(n_1916)
);

A2O1A1Ixp33_ASAP7_75t_L g1917 ( 
.A1(n_1765),
.A2(n_1232),
.B(n_1233),
.C(n_1226),
.Y(n_1917)
);

BUFx6f_ASAP7_75t_L g1918 ( 
.A(n_1735),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1821),
.B(n_1241),
.Y(n_1919)
);

INVx3_ASAP7_75t_L g1920 ( 
.A(n_1804),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1780),
.A2(n_736),
.B(n_735),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1727),
.A2(n_739),
.B(n_738),
.Y(n_1922)
);

CKINVDCx16_ASAP7_75t_R g1923 ( 
.A(n_1806),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1726),
.Y(n_1924)
);

AO21x1_ASAP7_75t_L g1925 ( 
.A1(n_1746),
.A2(n_1771),
.B(n_1818),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1737),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1758),
.Y(n_1927)
);

OAI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1819),
.A2(n_1822),
.B(n_1827),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1756),
.A2(n_742),
.B(n_741),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1762),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_SL g1931 ( 
.A(n_1767),
.B(n_1704),
.Y(n_1931)
);

AOI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1803),
.A2(n_744),
.B(n_743),
.Y(n_1932)
);

AOI21x1_ASAP7_75t_L g1933 ( 
.A1(n_1773),
.A2(n_746),
.B(n_745),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1761),
.B(n_1242),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1705),
.A2(n_748),
.B(n_747),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1741),
.B(n_749),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1764),
.Y(n_1937)
);

BUFx12f_ASAP7_75t_L g1938 ( 
.A(n_1755),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1763),
.Y(n_1939)
);

AOI21xp5_ASAP7_75t_L g1940 ( 
.A1(n_1770),
.A2(n_751),
.B(n_750),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1776),
.B(n_1244),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1760),
.B(n_1247),
.Y(n_1942)
);

O2A1O1Ixp33_ASAP7_75t_SL g1943 ( 
.A1(n_1729),
.A2(n_753),
.B(n_755),
.C(n_752),
.Y(n_1943)
);

AOI21xp5_ASAP7_75t_L g1944 ( 
.A1(n_1739),
.A2(n_757),
.B(n_756),
.Y(n_1944)
);

AOI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1744),
.A2(n_1723),
.B(n_1672),
.Y(n_1945)
);

INVx2_ASAP7_75t_SL g1946 ( 
.A(n_1876),
.Y(n_1946)
);

A2O1A1Ixp33_ASAP7_75t_L g1947 ( 
.A1(n_1857),
.A2(n_1734),
.B(n_1777),
.C(n_1676),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1830),
.B(n_1743),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1863),
.A2(n_1672),
.B(n_1722),
.Y(n_1949)
);

AOI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1858),
.A2(n_1710),
.B1(n_1774),
.B2(n_1716),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_R g1951 ( 
.A(n_1867),
.B(n_1717),
.Y(n_1951)
);

AOI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1887),
.A2(n_1728),
.B(n_1718),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1837),
.B(n_1848),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1849),
.B(n_1768),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1852),
.Y(n_1955)
);

NAND2x1p5_ASAP7_75t_L g1956 ( 
.A(n_1920),
.B(n_1669),
.Y(n_1956)
);

NOR2xp33_ASAP7_75t_L g1957 ( 
.A(n_1859),
.B(n_1706),
.Y(n_1957)
);

AO22x1_ASAP7_75t_L g1958 ( 
.A1(n_1892),
.A2(n_1796),
.B1(n_1797),
.B2(n_1769),
.Y(n_1958)
);

A2O1A1Ixp33_ASAP7_75t_L g1959 ( 
.A1(n_1928),
.A2(n_1725),
.B(n_1707),
.C(n_1720),
.Y(n_1959)
);

AOI22xp33_ASAP7_75t_SL g1960 ( 
.A1(n_1880),
.A2(n_1711),
.B1(n_1689),
.B2(n_1702),
.Y(n_1960)
);

A2O1A1Ixp33_ASAP7_75t_L g1961 ( 
.A1(n_1894),
.A2(n_1709),
.B(n_1696),
.C(n_1252),
.Y(n_1961)
);

O2A1O1Ixp5_ASAP7_75t_L g1962 ( 
.A1(n_1925),
.A2(n_1708),
.B(n_1711),
.C(n_2),
.Y(n_1962)
);

OAI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1881),
.A2(n_1255),
.B1(n_1256),
.B2(n_1250),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1861),
.Y(n_1964)
);

AOI21xp5_ASAP7_75t_L g1965 ( 
.A1(n_1902),
.A2(n_760),
.B(n_759),
.Y(n_1965)
);

BUFx2_ASAP7_75t_L g1966 ( 
.A(n_1938),
.Y(n_1966)
);

INVx2_ASAP7_75t_SL g1967 ( 
.A(n_1918),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_1923),
.Y(n_1968)
);

A2O1A1Ixp33_ASAP7_75t_L g1969 ( 
.A1(n_1911),
.A2(n_1261),
.B(n_1263),
.C(n_1259),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1871),
.B(n_1260),
.Y(n_1970)
);

NAND3xp33_ASAP7_75t_SL g1971 ( 
.A(n_1886),
.B(n_1906),
.C(n_1901),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1864),
.Y(n_1972)
);

OAI22x1_ASAP7_75t_L g1973 ( 
.A1(n_1855),
.A2(n_1265),
.B1(n_1269),
.B2(n_1264),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1877),
.Y(n_1974)
);

NAND3xp33_ASAP7_75t_SL g1975 ( 
.A(n_1865),
.B(n_1272),
.C(n_1271),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1905),
.B(n_1875),
.Y(n_1976)
);

BUFx6f_ASAP7_75t_L g1977 ( 
.A(n_1918),
.Y(n_1977)
);

AOI21xp5_ASAP7_75t_L g1978 ( 
.A1(n_1895),
.A2(n_1907),
.B(n_1945),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1835),
.B(n_1274),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1872),
.B(n_1275),
.Y(n_1980)
);

OAI22x1_ASAP7_75t_L g1981 ( 
.A1(n_1829),
.A2(n_1295),
.B1(n_1296),
.B2(n_1278),
.Y(n_1981)
);

AND2x4_ASAP7_75t_L g1982 ( 
.A(n_1896),
.B(n_761),
.Y(n_1982)
);

AND2x4_ASAP7_75t_L g1983 ( 
.A(n_1869),
.B(n_1878),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1833),
.Y(n_1984)
);

O2A1O1Ixp5_ASAP7_75t_L g1985 ( 
.A1(n_1891),
.A2(n_2),
.B(n_0),
.C(n_1),
.Y(n_1985)
);

A2O1A1Ixp33_ASAP7_75t_L g1986 ( 
.A1(n_1840),
.A2(n_1303),
.B(n_1308),
.C(n_1300),
.Y(n_1986)
);

AOI21x1_ASAP7_75t_L g1987 ( 
.A1(n_1933),
.A2(n_763),
.B(n_762),
.Y(n_1987)
);

AOI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1921),
.A2(n_766),
.B(n_765),
.Y(n_1988)
);

OAI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1853),
.A2(n_1321),
.B1(n_1323),
.B2(n_1311),
.Y(n_1989)
);

NOR2xp33_ASAP7_75t_L g1990 ( 
.A(n_1873),
.B(n_1329),
.Y(n_1990)
);

HB1xp67_ASAP7_75t_L g1991 ( 
.A(n_1850),
.Y(n_1991)
);

AOI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1879),
.A2(n_768),
.B(n_767),
.Y(n_1992)
);

O2A1O1Ixp33_ASAP7_75t_SL g1993 ( 
.A1(n_1870),
.A2(n_772),
.B(n_774),
.C(n_769),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1924),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1884),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1831),
.B(n_1332),
.Y(n_1996)
);

INVx4_ASAP7_75t_L g1997 ( 
.A(n_1850),
.Y(n_1997)
);

BUFx6f_ASAP7_75t_L g1998 ( 
.A(n_1845),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_R g1999 ( 
.A(n_1931),
.B(n_775),
.Y(n_1999)
);

AND2x6_ASAP7_75t_L g2000 ( 
.A(n_1936),
.B(n_776),
.Y(n_2000)
);

HB1xp67_ASAP7_75t_L g2001 ( 
.A(n_1845),
.Y(n_2001)
);

AOI22xp33_ASAP7_75t_L g2002 ( 
.A1(n_1900),
.A2(n_1341),
.B1(n_1344),
.B2(n_1338),
.Y(n_2002)
);

A2O1A1Ixp33_ASAP7_75t_L g2003 ( 
.A1(n_1842),
.A2(n_1360),
.B(n_1363),
.C(n_1357),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1874),
.B(n_1),
.Y(n_2004)
);

AOI22xp33_ASAP7_75t_L g2005 ( 
.A1(n_1838),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1889),
.B(n_3),
.Y(n_2006)
);

OAI21xp33_ASAP7_75t_L g2007 ( 
.A1(n_1832),
.A2(n_4),
.B(n_5),
.Y(n_2007)
);

OAI21xp5_ASAP7_75t_L g2008 ( 
.A1(n_1912),
.A2(n_778),
.B(n_777),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1899),
.B(n_6),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1898),
.Y(n_2010)
);

A2O1A1Ixp33_ASAP7_75t_L g2011 ( 
.A1(n_1844),
.A2(n_1866),
.B(n_1843),
.C(n_1841),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1934),
.B(n_6),
.Y(n_2012)
);

OAI22xp5_ASAP7_75t_L g2013 ( 
.A1(n_1927),
.A2(n_1930),
.B1(n_1904),
.B2(n_1926),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_R g2014 ( 
.A(n_1845),
.B(n_779),
.Y(n_2014)
);

A2O1A1Ixp33_ASAP7_75t_L g2015 ( 
.A1(n_1882),
.A2(n_9),
.B(n_7),
.C(n_8),
.Y(n_2015)
);

O2A1O1Ixp33_ASAP7_75t_SL g2016 ( 
.A1(n_1917),
.A2(n_1909),
.B(n_1885),
.C(n_1890),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1913),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1939),
.Y(n_2018)
);

AND2x4_ASAP7_75t_L g2019 ( 
.A(n_1897),
.B(n_780),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_SL g2020 ( 
.A(n_1937),
.B(n_7),
.Y(n_2020)
);

AOI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_1922),
.A2(n_783),
.B(n_781),
.Y(n_2021)
);

AOI21x1_ASAP7_75t_L g2022 ( 
.A1(n_1903),
.A2(n_786),
.B(n_784),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1941),
.B(n_9),
.Y(n_2023)
);

OAI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_1942),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_2024)
);

NOR2xp33_ASAP7_75t_L g2025 ( 
.A(n_1862),
.B(n_10),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1914),
.Y(n_2026)
);

OR2x6_ASAP7_75t_SL g2027 ( 
.A(n_1919),
.B(n_11),
.Y(n_2027)
);

OAI22x1_ASAP7_75t_L g2028 ( 
.A1(n_1828),
.A2(n_15),
.B1(n_16),
.B2(n_14),
.Y(n_2028)
);

INVx3_ASAP7_75t_L g2029 ( 
.A(n_1915),
.Y(n_2029)
);

INVx5_ASAP7_75t_L g2030 ( 
.A(n_1836),
.Y(n_2030)
);

AOI22xp5_ASAP7_75t_L g2031 ( 
.A1(n_1839),
.A2(n_16),
.B1(n_13),
.B2(n_15),
.Y(n_2031)
);

AOI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_1893),
.A2(n_789),
.B(n_787),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_SL g2033 ( 
.A(n_1834),
.B(n_13),
.Y(n_2033)
);

OAI22x1_ASAP7_75t_L g2034 ( 
.A1(n_1883),
.A2(n_19),
.B1(n_20),
.B2(n_18),
.Y(n_2034)
);

NOR2xp33_ASAP7_75t_L g2035 ( 
.A(n_1846),
.B(n_17),
.Y(n_2035)
);

BUFx6f_ASAP7_75t_L g2036 ( 
.A(n_1943),
.Y(n_2036)
);

BUFx12f_ASAP7_75t_L g2037 ( 
.A(n_1868),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1847),
.B(n_19),
.Y(n_2038)
);

BUFx6f_ASAP7_75t_L g2039 ( 
.A(n_1935),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1851),
.B(n_20),
.Y(n_2040)
);

BUFx6f_ASAP7_75t_L g2041 ( 
.A(n_1888),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1854),
.B(n_21),
.Y(n_2042)
);

NOR3xp33_ASAP7_75t_SL g2043 ( 
.A(n_1856),
.B(n_21),
.C(n_22),
.Y(n_2043)
);

OAI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_1860),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1916),
.B(n_25),
.Y(n_2045)
);

NOR2xp33_ASAP7_75t_R g2046 ( 
.A(n_1944),
.B(n_790),
.Y(n_2046)
);

AOI21xp5_ASAP7_75t_L g2047 ( 
.A1(n_1940),
.A2(n_792),
.B(n_791),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_L g2048 ( 
.A(n_1929),
.B(n_26),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_L g2049 ( 
.A(n_1932),
.B(n_27),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1908),
.Y(n_2050)
);

AOI21xp5_ASAP7_75t_L g2051 ( 
.A1(n_1910),
.A2(n_795),
.B(n_793),
.Y(n_2051)
);

CKINVDCx8_ASAP7_75t_R g2052 ( 
.A(n_1923),
.Y(n_2052)
);

INVxp33_ASAP7_75t_L g2053 ( 
.A(n_1835),
.Y(n_2053)
);

O2A1O1Ixp33_ASAP7_75t_SL g2054 ( 
.A1(n_1870),
.A2(n_798),
.B(n_799),
.C(n_797),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1852),
.Y(n_2055)
);

INVx3_ASAP7_75t_L g2056 ( 
.A(n_1918),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1852),
.Y(n_2057)
);

INVx1_ASAP7_75t_SL g2058 ( 
.A(n_1878),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_1880),
.B(n_27),
.Y(n_2059)
);

AOI21x1_ASAP7_75t_L g2060 ( 
.A1(n_1891),
.A2(n_801),
.B(n_800),
.Y(n_2060)
);

BUFx6f_ASAP7_75t_L g2061 ( 
.A(n_1918),
.Y(n_2061)
);

BUFx2_ASAP7_75t_SL g2062 ( 
.A(n_1867),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_L g2063 ( 
.A(n_1857),
.B(n_28),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1852),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1880),
.B(n_28),
.Y(n_2065)
);

AOI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_1830),
.A2(n_803),
.B(n_802),
.Y(n_2066)
);

O2A1O1Ixp33_ASAP7_75t_L g2067 ( 
.A1(n_1857),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1857),
.B(n_30),
.Y(n_2068)
);

AOI22xp33_ASAP7_75t_L g2069 ( 
.A1(n_1892),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_2069)
);

AOI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_1830),
.A2(n_807),
.B(n_805),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_1880),
.B(n_32),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1857),
.B(n_33),
.Y(n_2072)
);

O2A1O1Ixp33_ASAP7_75t_L g2073 ( 
.A1(n_1857),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_2073)
);

OAI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_1880),
.A2(n_37),
.B1(n_34),
.B2(n_36),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1857),
.B(n_37),
.Y(n_2075)
);

AOI21xp5_ASAP7_75t_L g2076 ( 
.A1(n_1948),
.A2(n_986),
.B(n_985),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1972),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1994),
.Y(n_2078)
);

A2O1A1Ixp33_ASAP7_75t_L g2079 ( 
.A1(n_2063),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_2079)
);

AOI21xp5_ASAP7_75t_L g2080 ( 
.A1(n_1978),
.A2(n_992),
.B(n_991),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_2018),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1957),
.B(n_39),
.Y(n_2082)
);

OAI22x1_ASAP7_75t_L g2083 ( 
.A1(n_1950),
.A2(n_44),
.B1(n_40),
.B2(n_41),
.Y(n_2083)
);

OAI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_2011),
.A2(n_41),
.B(n_44),
.Y(n_2084)
);

NAND3xp33_ASAP7_75t_L g2085 ( 
.A(n_2068),
.B(n_2075),
.C(n_2072),
.Y(n_2085)
);

AO31x2_ASAP7_75t_L g2086 ( 
.A1(n_2034),
.A2(n_1949),
.A3(n_2045),
.B(n_2050),
.Y(n_2086)
);

NOR2xp67_ASAP7_75t_L g2087 ( 
.A(n_2029),
.B(n_809),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1955),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1964),
.Y(n_2089)
);

HB1xp67_ASAP7_75t_L g2090 ( 
.A(n_2058),
.Y(n_2090)
);

OAI21x1_ASAP7_75t_L g2091 ( 
.A1(n_1987),
.A2(n_811),
.B(n_810),
.Y(n_2091)
);

OAI21x1_ASAP7_75t_L g2092 ( 
.A1(n_2022),
.A2(n_814),
.B(n_813),
.Y(n_2092)
);

INVx2_ASAP7_75t_SL g2093 ( 
.A(n_1977),
.Y(n_2093)
);

AOI22xp5_ASAP7_75t_L g2094 ( 
.A1(n_1980),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_2094)
);

BUFx4f_ASAP7_75t_SL g2095 ( 
.A(n_1977),
.Y(n_2095)
);

NOR2xp33_ASAP7_75t_L g2096 ( 
.A(n_2053),
.B(n_1953),
.Y(n_2096)
);

A2O1A1Ixp33_ASAP7_75t_L g2097 ( 
.A1(n_2048),
.A2(n_48),
.B(n_45),
.C(n_46),
.Y(n_2097)
);

OA21x2_ASAP7_75t_L g2098 ( 
.A1(n_2008),
.A2(n_816),
.B(n_815),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2026),
.B(n_48),
.Y(n_2099)
);

OAI21x1_ASAP7_75t_L g2100 ( 
.A1(n_2060),
.A2(n_819),
.B(n_817),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2004),
.B(n_49),
.Y(n_2101)
);

OAI21x1_ASAP7_75t_L g2102 ( 
.A1(n_2066),
.A2(n_821),
.B(n_820),
.Y(n_2102)
);

AOI21xp5_ASAP7_75t_L g2103 ( 
.A1(n_1971),
.A2(n_977),
.B(n_975),
.Y(n_2103)
);

OAI22xp5_ASAP7_75t_L g2104 ( 
.A1(n_1990),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_2104)
);

OAI21x1_ASAP7_75t_L g2105 ( 
.A1(n_2070),
.A2(n_824),
.B(n_822),
.Y(n_2105)
);

AOI21xp5_ASAP7_75t_L g2106 ( 
.A1(n_2016),
.A2(n_981),
.B(n_980),
.Y(n_2106)
);

AOI21xp33_ASAP7_75t_L g2107 ( 
.A1(n_1947),
.A2(n_50),
.B(n_52),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2065),
.B(n_52),
.Y(n_2108)
);

INVx4_ASAP7_75t_L g2109 ( 
.A(n_2061),
.Y(n_2109)
);

OAI21xp5_ASAP7_75t_L g2110 ( 
.A1(n_1959),
.A2(n_53),
.B(n_54),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1974),
.Y(n_2111)
);

OAI21x1_ASAP7_75t_L g2112 ( 
.A1(n_1965),
.A2(n_829),
.B(n_826),
.Y(n_2112)
);

NOR2xp33_ASAP7_75t_SL g2113 ( 
.A(n_2052),
.B(n_1968),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2055),
.Y(n_2114)
);

AOI21xp5_ASAP7_75t_L g2115 ( 
.A1(n_2041),
.A2(n_990),
.B(n_833),
.Y(n_2115)
);

A2O1A1Ixp33_ASAP7_75t_L g2116 ( 
.A1(n_2049),
.A2(n_55),
.B(n_53),
.C(n_54),
.Y(n_2116)
);

AOI21xp5_ASAP7_75t_L g2117 ( 
.A1(n_2041),
.A2(n_972),
.B(n_971),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_1979),
.B(n_55),
.Y(n_2118)
);

AOI21xp5_ASAP7_75t_L g2119 ( 
.A1(n_2039),
.A2(n_974),
.B(n_973),
.Y(n_2119)
);

AOI21xp5_ASAP7_75t_L g2120 ( 
.A1(n_2039),
.A2(n_979),
.B(n_978),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1976),
.B(n_56),
.Y(n_2121)
);

AO31x2_ASAP7_75t_L g2122 ( 
.A1(n_2021),
.A2(n_834),
.A3(n_835),
.B(n_830),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2057),
.Y(n_2123)
);

AOI221x1_ASAP7_75t_L g2124 ( 
.A1(n_2007),
.A2(n_59),
.B1(n_56),
.B2(n_57),
.C(n_60),
.Y(n_2124)
);

NOR2xp33_ASAP7_75t_L g2125 ( 
.A(n_1970),
.B(n_836),
.Y(n_2125)
);

AOI21xp5_ASAP7_75t_L g2126 ( 
.A1(n_2047),
.A2(n_969),
.B(n_968),
.Y(n_2126)
);

INVx2_ASAP7_75t_SL g2127 ( 
.A(n_2061),
.Y(n_2127)
);

OAI21xp5_ASAP7_75t_L g2128 ( 
.A1(n_1969),
.A2(n_59),
.B(n_61),
.Y(n_2128)
);

AOI21xp5_ASAP7_75t_SL g2129 ( 
.A1(n_1954),
.A2(n_841),
.B(n_838),
.Y(n_2129)
);

OAI21x1_ASAP7_75t_L g2130 ( 
.A1(n_2032),
.A2(n_1992),
.B(n_1988),
.Y(n_2130)
);

NOR2x1_ASAP7_75t_SL g2131 ( 
.A(n_2036),
.B(n_843),
.Y(n_2131)
);

OAI22xp5_ASAP7_75t_L g2132 ( 
.A1(n_2002),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_2132)
);

OAI21xp5_ASAP7_75t_L g2133 ( 
.A1(n_1996),
.A2(n_62),
.B(n_64),
.Y(n_2133)
);

INVx1_ASAP7_75t_SL g2134 ( 
.A(n_1951),
.Y(n_2134)
);

OAI21xp5_ASAP7_75t_L g2135 ( 
.A1(n_2012),
.A2(n_64),
.B(n_65),
.Y(n_2135)
);

NOR2xp67_ASAP7_75t_L g2136 ( 
.A(n_1983),
.B(n_845),
.Y(n_2136)
);

AO21x2_ASAP7_75t_L g2137 ( 
.A1(n_1975),
.A2(n_847),
.B(n_846),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2025),
.B(n_1995),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2006),
.B(n_65),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2064),
.Y(n_2140)
);

AOI21xp5_ASAP7_75t_L g2141 ( 
.A1(n_2051),
.A2(n_984),
.B(n_849),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_2009),
.B(n_66),
.Y(n_2142)
);

BUFx12f_ASAP7_75t_L g2143 ( 
.A(n_1966),
.Y(n_2143)
);

AOI21xp5_ASAP7_75t_L g2144 ( 
.A1(n_1952),
.A2(n_967),
.B(n_965),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_SL g2145 ( 
.A(n_1960),
.B(n_66),
.Y(n_2145)
);

NOR2xp33_ASAP7_75t_L g2146 ( 
.A(n_2059),
.B(n_848),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_2010),
.Y(n_2147)
);

A2O1A1Ixp33_ASAP7_75t_L g2148 ( 
.A1(n_2035),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1958),
.B(n_67),
.Y(n_2149)
);

OAI21x1_ASAP7_75t_L g2150 ( 
.A1(n_1985),
.A2(n_854),
.B(n_851),
.Y(n_2150)
);

NOR2xp33_ASAP7_75t_L g2151 ( 
.A(n_2071),
.B(n_856),
.Y(n_2151)
);

OA21x2_ASAP7_75t_L g2152 ( 
.A1(n_1962),
.A2(n_858),
.B(n_857),
.Y(n_2152)
);

INVx4_ASAP7_75t_L g2153 ( 
.A(n_1998),
.Y(n_2153)
);

INVx1_ASAP7_75t_SL g2154 ( 
.A(n_2062),
.Y(n_2154)
);

OAI21xp5_ASAP7_75t_L g2155 ( 
.A1(n_1986),
.A2(n_68),
.B(n_69),
.Y(n_2155)
);

OAI21xp33_ASAP7_75t_L g2156 ( 
.A1(n_2069),
.A2(n_70),
.B(n_71),
.Y(n_2156)
);

O2A1O1Ixp5_ASAP7_75t_SL g2157 ( 
.A1(n_2024),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_2157)
);

AOI221x1_ASAP7_75t_L g2158 ( 
.A1(n_2015),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.C(n_76),
.Y(n_2158)
);

INVx2_ASAP7_75t_SL g2159 ( 
.A(n_2095),
.Y(n_2159)
);

NOR2xp67_ASAP7_75t_L g2160 ( 
.A(n_2085),
.B(n_1984),
.Y(n_2160)
);

OAI21x1_ASAP7_75t_L g2161 ( 
.A1(n_2130),
.A2(n_2013),
.B(n_2033),
.Y(n_2161)
);

AO21x2_ASAP7_75t_L g2162 ( 
.A1(n_2084),
.A2(n_2046),
.B(n_1993),
.Y(n_2162)
);

NAND2x1p5_ASAP7_75t_L g2163 ( 
.A(n_2154),
.B(n_1997),
.Y(n_2163)
);

OAI21x1_ASAP7_75t_SL g2164 ( 
.A1(n_2110),
.A2(n_2073),
.B(n_2067),
.Y(n_2164)
);

INVx2_ASAP7_75t_SL g2165 ( 
.A(n_2093),
.Y(n_2165)
);

NOR2xp33_ASAP7_75t_L g2166 ( 
.A(n_2096),
.B(n_2027),
.Y(n_2166)
);

NOR2xp33_ASAP7_75t_L g2167 ( 
.A(n_2134),
.B(n_2090),
.Y(n_2167)
);

A2O1A1Ixp33_ASAP7_75t_L g2168 ( 
.A1(n_2128),
.A2(n_2040),
.B(n_2038),
.C(n_2043),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2088),
.Y(n_2169)
);

OAI21x1_ASAP7_75t_L g2170 ( 
.A1(n_2100),
.A2(n_2080),
.B(n_2091),
.Y(n_2170)
);

INVxp67_ASAP7_75t_L g2171 ( 
.A(n_2138),
.Y(n_2171)
);

AOI22xp33_ASAP7_75t_L g2172 ( 
.A1(n_2156),
.A2(n_2074),
.B1(n_2044),
.B2(n_2037),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2121),
.B(n_2023),
.Y(n_2173)
);

BUFx3_ASAP7_75t_L g2174 ( 
.A(n_2127),
.Y(n_2174)
);

INVx3_ASAP7_75t_L g2175 ( 
.A(n_2109),
.Y(n_2175)
);

OAI21x1_ASAP7_75t_L g2176 ( 
.A1(n_2106),
.A2(n_2042),
.B(n_2017),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2077),
.Y(n_2177)
);

AOI221xp5_ASAP7_75t_L g2178 ( 
.A1(n_2107),
.A2(n_1963),
.B1(n_2005),
.B2(n_2028),
.C(n_2031),
.Y(n_2178)
);

INVx3_ASAP7_75t_L g2179 ( 
.A(n_2153),
.Y(n_2179)
);

INVx3_ASAP7_75t_L g2180 ( 
.A(n_2143),
.Y(n_2180)
);

CKINVDCx11_ASAP7_75t_R g2181 ( 
.A(n_2113),
.Y(n_2181)
);

NOR2xp33_ASAP7_75t_L g2182 ( 
.A(n_2125),
.B(n_2145),
.Y(n_2182)
);

OA21x2_ASAP7_75t_L g2183 ( 
.A1(n_2150),
.A2(n_2020),
.B(n_1961),
.Y(n_2183)
);

OAI21x1_ASAP7_75t_L g2184 ( 
.A1(n_2092),
.A2(n_1956),
.B(n_2054),
.Y(n_2184)
);

A2O1A1Ixp33_ASAP7_75t_L g2185 ( 
.A1(n_2155),
.A2(n_2003),
.B(n_2036),
.C(n_1982),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2082),
.B(n_2000),
.Y(n_2186)
);

OAI21x1_ASAP7_75t_L g2187 ( 
.A1(n_2102),
.A2(n_2001),
.B(n_1989),
.Y(n_2187)
);

INVx2_ASAP7_75t_SL g2188 ( 
.A(n_2081),
.Y(n_2188)
);

AOI22xp33_ASAP7_75t_L g2189 ( 
.A1(n_2133),
.A2(n_1973),
.B1(n_1981),
.B2(n_2000),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2135),
.B(n_2000),
.Y(n_2190)
);

NAND3xp33_ASAP7_75t_L g2191 ( 
.A(n_2079),
.B(n_2019),
.C(n_1991),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_2078),
.Y(n_2192)
);

INVx3_ASAP7_75t_L g2193 ( 
.A(n_2147),
.Y(n_2193)
);

AND2x4_ASAP7_75t_L g2194 ( 
.A(n_2136),
.B(n_1967),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2089),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2099),
.B(n_1999),
.Y(n_2196)
);

AO21x1_ASAP7_75t_L g2197 ( 
.A1(n_2132),
.A2(n_2104),
.B(n_2103),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2111),
.Y(n_2198)
);

OR2x6_ASAP7_75t_L g2199 ( 
.A(n_2129),
.B(n_1946),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2114),
.Y(n_2200)
);

NAND2x1p5_ASAP7_75t_L g2201 ( 
.A(n_2087),
.B(n_2056),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2123),
.Y(n_2202)
);

AO21x2_ASAP7_75t_L g2203 ( 
.A1(n_2144),
.A2(n_2014),
.B(n_1998),
.Y(n_2203)
);

OAI21x1_ASAP7_75t_L g2204 ( 
.A1(n_2105),
.A2(n_860),
.B(n_859),
.Y(n_2204)
);

AOI22xp33_ASAP7_75t_L g2205 ( 
.A1(n_2083),
.A2(n_2030),
.B1(n_76),
.B2(n_73),
.Y(n_2205)
);

HB1xp67_ASAP7_75t_L g2206 ( 
.A(n_2140),
.Y(n_2206)
);

AOI22xp33_ASAP7_75t_SL g2207 ( 
.A1(n_2146),
.A2(n_2030),
.B1(n_78),
.B2(n_74),
.Y(n_2207)
);

OAI21x1_ASAP7_75t_L g2208 ( 
.A1(n_2112),
.A2(n_862),
.B(n_861),
.Y(n_2208)
);

AO21x2_ASAP7_75t_L g2209 ( 
.A1(n_2126),
.A2(n_77),
.B(n_78),
.Y(n_2209)
);

OA21x2_ASAP7_75t_L g2210 ( 
.A1(n_2184),
.A2(n_2158),
.B(n_2124),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2206),
.Y(n_2211)
);

AO21x1_ASAP7_75t_L g2212 ( 
.A1(n_2182),
.A2(n_2149),
.B(n_2142),
.Y(n_2212)
);

AOI21xp5_ASAP7_75t_L g2213 ( 
.A1(n_2162),
.A2(n_2168),
.B(n_2164),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2195),
.Y(n_2214)
);

AOI21xp5_ASAP7_75t_L g2215 ( 
.A1(n_2164),
.A2(n_2098),
.B(n_2141),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2171),
.B(n_2139),
.Y(n_2216)
);

BUFx10_ASAP7_75t_L g2217 ( 
.A(n_2159),
.Y(n_2217)
);

OA21x2_ASAP7_75t_L g2218 ( 
.A1(n_2187),
.A2(n_2116),
.B(n_2097),
.Y(n_2218)
);

AO21x2_ASAP7_75t_L g2219 ( 
.A1(n_2161),
.A2(n_2076),
.B(n_2148),
.Y(n_2219)
);

INVx3_ASAP7_75t_L g2220 ( 
.A(n_2174),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2177),
.B(n_2101),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2169),
.Y(n_2222)
);

OR2x2_ASAP7_75t_L g2223 ( 
.A(n_2198),
.B(n_2086),
.Y(n_2223)
);

OAI21x1_ASAP7_75t_L g2224 ( 
.A1(n_2170),
.A2(n_2117),
.B(n_2115),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_2200),
.B(n_2086),
.Y(n_2225)
);

AND2x4_ASAP7_75t_L g2226 ( 
.A(n_2188),
.B(n_2131),
.Y(n_2226)
);

AOI21xp5_ASAP7_75t_L g2227 ( 
.A1(n_2185),
.A2(n_2120),
.B(n_2119),
.Y(n_2227)
);

BUFx2_ASAP7_75t_L g2228 ( 
.A(n_2163),
.Y(n_2228)
);

BUFx4f_ASAP7_75t_SL g2229 ( 
.A(n_2180),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_2202),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2192),
.B(n_2118),
.Y(n_2231)
);

OAI21x1_ASAP7_75t_L g2232 ( 
.A1(n_2176),
.A2(n_2204),
.B(n_2208),
.Y(n_2232)
);

CKINVDCx11_ASAP7_75t_R g2233 ( 
.A(n_2181),
.Y(n_2233)
);

A2O1A1Ixp33_ASAP7_75t_L g2234 ( 
.A1(n_2178),
.A2(n_2151),
.B(n_2094),
.C(n_2108),
.Y(n_2234)
);

OR2x2_ASAP7_75t_L g2235 ( 
.A(n_2173),
.B(n_2152),
.Y(n_2235)
);

OAI21x1_ASAP7_75t_L g2236 ( 
.A1(n_2183),
.A2(n_2157),
.B(n_2122),
.Y(n_2236)
);

INVx2_ASAP7_75t_SL g2237 ( 
.A(n_2165),
.Y(n_2237)
);

OA21x2_ASAP7_75t_L g2238 ( 
.A1(n_2190),
.A2(n_2122),
.B(n_2137),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2160),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2193),
.B(n_77),
.Y(n_2240)
);

OR2x6_ASAP7_75t_L g2241 ( 
.A(n_2199),
.B(n_2030),
.Y(n_2241)
);

OA21x2_ASAP7_75t_L g2242 ( 
.A1(n_2189),
.A2(n_79),
.B(n_80),
.Y(n_2242)
);

OA21x2_ASAP7_75t_L g2243 ( 
.A1(n_2186),
.A2(n_2191),
.B(n_2197),
.Y(n_2243)
);

OR2x2_ASAP7_75t_L g2244 ( 
.A(n_2196),
.B(n_79),
.Y(n_2244)
);

CKINVDCx5p33_ASAP7_75t_R g2245 ( 
.A(n_2167),
.Y(n_2245)
);

AO21x2_ASAP7_75t_L g2246 ( 
.A1(n_2209),
.A2(n_81),
.B(n_82),
.Y(n_2246)
);

OAI21x1_ASAP7_75t_L g2247 ( 
.A1(n_2183),
.A2(n_864),
.B(n_863),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2203),
.Y(n_2248)
);

AOI21xp33_ASAP7_75t_L g2249 ( 
.A1(n_2172),
.A2(n_2166),
.B(n_2199),
.Y(n_2249)
);

INVx3_ASAP7_75t_L g2250 ( 
.A(n_2175),
.Y(n_2250)
);

AOI21xp5_ASAP7_75t_L g2251 ( 
.A1(n_2201),
.A2(n_867),
.B(n_866),
.Y(n_2251)
);

INVx2_ASAP7_75t_SL g2252 ( 
.A(n_2179),
.Y(n_2252)
);

HB1xp67_ASAP7_75t_L g2253 ( 
.A(n_2194),
.Y(n_2253)
);

AO21x2_ASAP7_75t_L g2254 ( 
.A1(n_2207),
.A2(n_83),
.B(n_84),
.Y(n_2254)
);

CKINVDCx9p33_ASAP7_75t_R g2255 ( 
.A(n_2205),
.Y(n_2255)
);

A2O1A1Ixp33_ASAP7_75t_L g2256 ( 
.A1(n_2182),
.A2(n_85),
.B(n_83),
.C(n_84),
.Y(n_2256)
);

CKINVDCx20_ASAP7_75t_R g2257 ( 
.A(n_2181),
.Y(n_2257)
);

INVxp67_ASAP7_75t_L g2258 ( 
.A(n_2167),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2206),
.Y(n_2259)
);

AOI21xp5_ASAP7_75t_L g2260 ( 
.A1(n_2162),
.A2(n_869),
.B(n_868),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2195),
.Y(n_2261)
);

BUFx8_ASAP7_75t_L g2262 ( 
.A(n_2159),
.Y(n_2262)
);

AO21x2_ASAP7_75t_L g2263 ( 
.A1(n_2213),
.A2(n_85),
.B(n_86),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_2230),
.Y(n_2264)
);

OAI21x1_ASAP7_75t_L g2265 ( 
.A1(n_2215),
.A2(n_872),
.B(n_870),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2214),
.Y(n_2266)
);

OAI21x1_ASAP7_75t_L g2267 ( 
.A1(n_2232),
.A2(n_876),
.B(n_875),
.Y(n_2267)
);

BUFx2_ASAP7_75t_L g2268 ( 
.A(n_2228),
.Y(n_2268)
);

HB1xp67_ASAP7_75t_L g2269 ( 
.A(n_2211),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2222),
.Y(n_2270)
);

AOI21x1_ASAP7_75t_L g2271 ( 
.A1(n_2212),
.A2(n_87),
.B(n_88),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_2261),
.Y(n_2272)
);

BUFx3_ASAP7_75t_L g2273 ( 
.A(n_2262),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2259),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_2253),
.B(n_87),
.Y(n_2275)
);

OR2x2_ASAP7_75t_L g2276 ( 
.A(n_2223),
.B(n_88),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_2239),
.Y(n_2277)
);

BUFx2_ASAP7_75t_L g2278 ( 
.A(n_2241),
.Y(n_2278)
);

OAI21x1_ASAP7_75t_L g2279 ( 
.A1(n_2224),
.A2(n_878),
.B(n_877),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2225),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2225),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2248),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2235),
.Y(n_2283)
);

HB1xp67_ASAP7_75t_L g2284 ( 
.A(n_2243),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2238),
.Y(n_2285)
);

OR2x2_ASAP7_75t_L g2286 ( 
.A(n_2216),
.B(n_2231),
.Y(n_2286)
);

BUFx2_ASAP7_75t_L g2287 ( 
.A(n_2241),
.Y(n_2287)
);

HB1xp67_ASAP7_75t_L g2288 ( 
.A(n_2221),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2246),
.Y(n_2289)
);

BUFx6f_ASAP7_75t_L g2290 ( 
.A(n_2233),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2237),
.Y(n_2291)
);

OR2x2_ASAP7_75t_L g2292 ( 
.A(n_2258),
.B(n_89),
.Y(n_2292)
);

INVx4_ASAP7_75t_L g2293 ( 
.A(n_2229),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2236),
.Y(n_2294)
);

AOI21x1_ASAP7_75t_L g2295 ( 
.A1(n_2260),
.A2(n_89),
.B(n_90),
.Y(n_2295)
);

AND2x4_ASAP7_75t_L g2296 ( 
.A(n_2226),
.B(n_879),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2240),
.Y(n_2297)
);

AND2x4_ASAP7_75t_L g2298 ( 
.A(n_2220),
.B(n_880),
.Y(n_2298)
);

INVx2_ASAP7_75t_SL g2299 ( 
.A(n_2252),
.Y(n_2299)
);

INVxp67_ASAP7_75t_L g2300 ( 
.A(n_2244),
.Y(n_2300)
);

NAND3xp33_ASAP7_75t_L g2301 ( 
.A(n_2256),
.B(n_90),
.C(n_91),
.Y(n_2301)
);

AOI21x1_ASAP7_75t_L g2302 ( 
.A1(n_2227),
.A2(n_93),
.B(n_94),
.Y(n_2302)
);

INVx3_ASAP7_75t_L g2303 ( 
.A(n_2250),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2210),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2218),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2242),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2247),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2245),
.B(n_93),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2219),
.Y(n_2309)
);

AO31x2_ASAP7_75t_L g2310 ( 
.A1(n_2234),
.A2(n_97),
.A3(n_95),
.B(n_96),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2254),
.Y(n_2311)
);

AO21x2_ASAP7_75t_L g2312 ( 
.A1(n_2249),
.A2(n_2251),
.B(n_2255),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2217),
.Y(n_2313)
);

OR2x2_ASAP7_75t_L g2314 ( 
.A(n_2257),
.B(n_95),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2211),
.B(n_96),
.Y(n_2315)
);

AO21x2_ASAP7_75t_L g2316 ( 
.A1(n_2213),
.A2(n_98),
.B(n_99),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2222),
.Y(n_2317)
);

HB1xp67_ASAP7_75t_L g2318 ( 
.A(n_2211),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2211),
.B(n_98),
.Y(n_2319)
);

OA21x2_ASAP7_75t_L g2320 ( 
.A1(n_2213),
.A2(n_107),
.B(n_99),
.Y(n_2320)
);

AOI22xp33_ASAP7_75t_L g2321 ( 
.A1(n_2212),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_2321)
);

INVx3_ASAP7_75t_L g2322 ( 
.A(n_2250),
.Y(n_2322)
);

INVx1_ASAP7_75t_SL g2323 ( 
.A(n_2245),
.Y(n_2323)
);

HB1xp67_ASAP7_75t_L g2324 ( 
.A(n_2211),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_2230),
.Y(n_2325)
);

INVx3_ASAP7_75t_L g2326 ( 
.A(n_2250),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2222),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2211),
.B(n_100),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2222),
.Y(n_2329)
);

AOI21x1_ASAP7_75t_L g2330 ( 
.A1(n_2212),
.A2(n_101),
.B(n_103),
.Y(n_2330)
);

INVx3_ASAP7_75t_L g2331 ( 
.A(n_2250),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2211),
.B(n_103),
.Y(n_2332)
);

INVx3_ASAP7_75t_L g2333 ( 
.A(n_2250),
.Y(n_2333)
);

OA21x2_ASAP7_75t_L g2334 ( 
.A1(n_2213),
.A2(n_112),
.B(n_104),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_2233),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_2211),
.B(n_104),
.Y(n_2336)
);

OAI21xp5_ASAP7_75t_L g2337 ( 
.A1(n_2213),
.A2(n_105),
.B(n_106),
.Y(n_2337)
);

BUFx3_ASAP7_75t_L g2338 ( 
.A(n_2262),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2277),
.Y(n_2339)
);

OAI22xp33_ASAP7_75t_L g2340 ( 
.A1(n_2337),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2270),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2317),
.Y(n_2342)
);

OAI22xp5_ASAP7_75t_L g2343 ( 
.A1(n_2301),
.A2(n_2321),
.B1(n_2311),
.B2(n_2278),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2327),
.Y(n_2344)
);

BUFx2_ASAP7_75t_L g2345 ( 
.A(n_2268),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_2288),
.B(n_108),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2329),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2269),
.B(n_108),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2318),
.B(n_109),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2324),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2280),
.Y(n_2351)
);

BUFx3_ASAP7_75t_L g2352 ( 
.A(n_2290),
.Y(n_2352)
);

AOI21xp5_ASAP7_75t_L g2353 ( 
.A1(n_2312),
.A2(n_882),
.B(n_881),
.Y(n_2353)
);

AOI22xp33_ASAP7_75t_L g2354 ( 
.A1(n_2287),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_2354)
);

AOI21xp5_ASAP7_75t_L g2355 ( 
.A1(n_2284),
.A2(n_884),
.B(n_883),
.Y(n_2355)
);

OAI22xp33_ASAP7_75t_L g2356 ( 
.A1(n_2306),
.A2(n_113),
.B1(n_110),
.B2(n_111),
.Y(n_2356)
);

OA21x2_ASAP7_75t_L g2357 ( 
.A1(n_2304),
.A2(n_113),
.B(n_114),
.Y(n_2357)
);

OAI211xp5_ASAP7_75t_L g2358 ( 
.A1(n_2271),
.A2(n_2330),
.B(n_2320),
.C(n_2334),
.Y(n_2358)
);

AOI211xp5_ASAP7_75t_L g2359 ( 
.A1(n_2289),
.A2(n_116),
.B(n_114),
.C(n_115),
.Y(n_2359)
);

AOI221xp5_ASAP7_75t_L g2360 ( 
.A1(n_2297),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.C(n_118),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2283),
.B(n_117),
.Y(n_2361)
);

BUFx2_ASAP7_75t_L g2362 ( 
.A(n_2303),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2264),
.Y(n_2363)
);

INVx4_ASAP7_75t_L g2364 ( 
.A(n_2290),
.Y(n_2364)
);

AO31x2_ASAP7_75t_L g2365 ( 
.A1(n_2309),
.A2(n_121),
.A3(n_119),
.B(n_120),
.Y(n_2365)
);

AOI22xp33_ASAP7_75t_L g2366 ( 
.A1(n_2263),
.A2(n_122),
.B1(n_119),
.B2(n_121),
.Y(n_2366)
);

OAI211xp5_ASAP7_75t_L g2367 ( 
.A1(n_2302),
.A2(n_126),
.B(n_124),
.C(n_125),
.Y(n_2367)
);

INVx5_ASAP7_75t_L g2368 ( 
.A(n_2293),
.Y(n_2368)
);

OAI21x1_ASAP7_75t_L g2369 ( 
.A1(n_2285),
.A2(n_125),
.B(n_126),
.Y(n_2369)
);

AOI22xp33_ASAP7_75t_SL g2370 ( 
.A1(n_2316),
.A2(n_129),
.B1(n_130),
.B2(n_128),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2281),
.Y(n_2371)
);

AOI22xp33_ASAP7_75t_L g2372 ( 
.A1(n_2300),
.A2(n_131),
.B1(n_127),
.B2(n_130),
.Y(n_2372)
);

AOI22xp33_ASAP7_75t_L g2373 ( 
.A1(n_2314),
.A2(n_132),
.B1(n_127),
.B2(n_131),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2286),
.B(n_133),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_2274),
.B(n_133),
.Y(n_2375)
);

BUFx4f_ASAP7_75t_SL g2376 ( 
.A(n_2273),
.Y(n_2376)
);

AOI22xp33_ASAP7_75t_L g2377 ( 
.A1(n_2314),
.A2(n_2313),
.B1(n_2286),
.B2(n_2308),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2325),
.Y(n_2378)
);

AOI22xp33_ASAP7_75t_L g2379 ( 
.A1(n_2305),
.A2(n_137),
.B1(n_134),
.B2(n_136),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2266),
.Y(n_2380)
);

BUFx6f_ASAP7_75t_L g2381 ( 
.A(n_2338),
.Y(n_2381)
);

OAI221xp5_ASAP7_75t_L g2382 ( 
.A1(n_2315),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.C(n_139),
.Y(n_2382)
);

NOR3xp33_ASAP7_75t_L g2383 ( 
.A(n_2295),
.B(n_139),
.C(n_140),
.Y(n_2383)
);

NAND3xp33_ASAP7_75t_L g2384 ( 
.A(n_2294),
.B(n_140),
.C(n_141),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2272),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2282),
.Y(n_2386)
);

AOI22xp33_ASAP7_75t_SL g2387 ( 
.A1(n_2265),
.A2(n_144),
.B1(n_145),
.B2(n_143),
.Y(n_2387)
);

AOI22xp33_ASAP7_75t_L g2388 ( 
.A1(n_2296),
.A2(n_2326),
.B1(n_2331),
.B2(n_2322),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2276),
.Y(n_2389)
);

AOI22xp33_ASAP7_75t_L g2390 ( 
.A1(n_2333),
.A2(n_2307),
.B1(n_2291),
.B2(n_2299),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_L g2391 ( 
.A(n_2323),
.B(n_2335),
.Y(n_2391)
);

BUFx4f_ASAP7_75t_SL g2392 ( 
.A(n_2292),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2276),
.Y(n_2393)
);

AO21x2_ASAP7_75t_L g2394 ( 
.A1(n_2319),
.A2(n_142),
.B(n_143),
.Y(n_2394)
);

AOI22xp33_ASAP7_75t_SL g2395 ( 
.A1(n_2275),
.A2(n_147),
.B1(n_148),
.B2(n_146),
.Y(n_2395)
);

AOI221xp5_ASAP7_75t_L g2396 ( 
.A1(n_2328),
.A2(n_147),
.B1(n_142),
.B2(n_146),
.C(n_148),
.Y(n_2396)
);

OAI21x1_ASAP7_75t_SL g2397 ( 
.A1(n_2292),
.A2(n_149),
.B(n_150),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2332),
.Y(n_2398)
);

AOI221xp5_ASAP7_75t_L g2399 ( 
.A1(n_2336),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.C(n_152),
.Y(n_2399)
);

OAI22xp5_ASAP7_75t_L g2400 ( 
.A1(n_2298),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2310),
.Y(n_2401)
);

AOI22xp33_ASAP7_75t_L g2402 ( 
.A1(n_2279),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.Y(n_2402)
);

OAI21x1_ASAP7_75t_L g2403 ( 
.A1(n_2267),
.A2(n_2310),
.B(n_156),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2277),
.Y(n_2404)
);

BUFx8_ASAP7_75t_SL g2405 ( 
.A(n_2290),
.Y(n_2405)
);

OAI22xp5_ASAP7_75t_L g2406 ( 
.A1(n_2301),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_2406)
);

AOI22xp33_ASAP7_75t_L g2407 ( 
.A1(n_2337),
.A2(n_160),
.B1(n_157),
.B2(n_159),
.Y(n_2407)
);

INVx2_ASAP7_75t_SL g2408 ( 
.A(n_2299),
.Y(n_2408)
);

AOI21x1_ASAP7_75t_L g2409 ( 
.A1(n_2284),
.A2(n_159),
.B(n_161),
.Y(n_2409)
);

AOI22xp33_ASAP7_75t_L g2410 ( 
.A1(n_2337),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.Y(n_2410)
);

AOI22xp33_ASAP7_75t_L g2411 ( 
.A1(n_2337),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2270),
.Y(n_2412)
);

OAI22xp5_ASAP7_75t_L g2413 ( 
.A1(n_2301),
.A2(n_167),
.B1(n_164),
.B2(n_165),
.Y(n_2413)
);

OAI33xp33_ASAP7_75t_L g2414 ( 
.A1(n_2311),
.A2(n_169),
.A3(n_171),
.B1(n_165),
.B2(n_167),
.B3(n_170),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2270),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2268),
.B(n_169),
.Y(n_2416)
);

AOI221xp5_ASAP7_75t_L g2417 ( 
.A1(n_2311),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.C(n_174),
.Y(n_2417)
);

OAI22xp33_ASAP7_75t_L g2418 ( 
.A1(n_2337),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_2418)
);

AOI22xp33_ASAP7_75t_L g2419 ( 
.A1(n_2337),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2270),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2270),
.Y(n_2421)
);

OAI22xp5_ASAP7_75t_L g2422 ( 
.A1(n_2301),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_2422)
);

OAI22xp5_ASAP7_75t_L g2423 ( 
.A1(n_2301),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.Y(n_2423)
);

AOI21xp5_ASAP7_75t_L g2424 ( 
.A1(n_2337),
.A2(n_888),
.B(n_885),
.Y(n_2424)
);

INVx1_ASAP7_75t_SL g2425 ( 
.A(n_2323),
.Y(n_2425)
);

OAI22xp5_ASAP7_75t_L g2426 ( 
.A1(n_2301),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_2426)
);

AOI22xp33_ASAP7_75t_L g2427 ( 
.A1(n_2337),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_2427)
);

AOI21xp5_ASAP7_75t_L g2428 ( 
.A1(n_2337),
.A2(n_891),
.B(n_889),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2268),
.B(n_182),
.Y(n_2429)
);

OR2x2_ASAP7_75t_L g2430 ( 
.A(n_2283),
.B(n_184),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2277),
.Y(n_2431)
);

NAND3xp33_ASAP7_75t_L g2432 ( 
.A(n_2337),
.B(n_184),
.C(n_185),
.Y(n_2432)
);

AND2x2_ASAP7_75t_L g2433 ( 
.A(n_2268),
.B(n_185),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2270),
.Y(n_2434)
);

AOI21xp33_ASAP7_75t_L g2435 ( 
.A1(n_2312),
.A2(n_186),
.B(n_187),
.Y(n_2435)
);

AOI22xp33_ASAP7_75t_L g2436 ( 
.A1(n_2337),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2342),
.Y(n_2437)
);

NOR2xp33_ASAP7_75t_L g2438 ( 
.A(n_2368),
.B(n_188),
.Y(n_2438)
);

AOI22xp33_ASAP7_75t_L g2439 ( 
.A1(n_2432),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.Y(n_2439)
);

INVx3_ASAP7_75t_SL g2440 ( 
.A(n_2364),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2412),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2386),
.Y(n_2442)
);

BUFx2_ASAP7_75t_L g2443 ( 
.A(n_2345),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2350),
.B(n_189),
.Y(n_2444)
);

HB1xp67_ASAP7_75t_L g2445 ( 
.A(n_2389),
.Y(n_2445)
);

OR2x2_ASAP7_75t_L g2446 ( 
.A(n_2393),
.B(n_2385),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2415),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2420),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_2362),
.B(n_192),
.Y(n_2449)
);

OAI22xp5_ASAP7_75t_L g2450 ( 
.A1(n_2407),
.A2(n_194),
.B1(n_192),
.B2(n_193),
.Y(n_2450)
);

NOR2x1p5_ASAP7_75t_L g2451 ( 
.A(n_2352),
.B(n_2381),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_2421),
.B(n_193),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_2390),
.B(n_195),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2408),
.B(n_195),
.Y(n_2454)
);

NAND2x1p5_ASAP7_75t_SL g2455 ( 
.A(n_2416),
.B(n_196),
.Y(n_2455)
);

INVxp67_ASAP7_75t_SL g2456 ( 
.A(n_2341),
.Y(n_2456)
);

AND2x4_ASAP7_75t_L g2457 ( 
.A(n_2368),
.B(n_196),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2434),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2344),
.Y(n_2459)
);

AND2x2_ASAP7_75t_L g2460 ( 
.A(n_2398),
.B(n_197),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2339),
.B(n_197),
.Y(n_2461)
);

NOR2xp33_ASAP7_75t_L g2462 ( 
.A(n_2368),
.B(n_2376),
.Y(n_2462)
);

AND2x2_ASAP7_75t_L g2463 ( 
.A(n_2404),
.B(n_198),
.Y(n_2463)
);

AND2x2_ASAP7_75t_L g2464 ( 
.A(n_2431),
.B(n_199),
.Y(n_2464)
);

OR2x2_ASAP7_75t_L g2465 ( 
.A(n_2378),
.B(n_200),
.Y(n_2465)
);

NOR2xp33_ASAP7_75t_L g2466 ( 
.A(n_2405),
.B(n_200),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2347),
.B(n_201),
.Y(n_2467)
);

INVx5_ASAP7_75t_L g2468 ( 
.A(n_2381),
.Y(n_2468)
);

NOR2xp33_ASAP7_75t_L g2469 ( 
.A(n_2391),
.B(n_202),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2351),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2363),
.B(n_202),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2380),
.B(n_2374),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2371),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2430),
.Y(n_2474)
);

BUFx2_ASAP7_75t_L g2475 ( 
.A(n_2392),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2375),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2361),
.B(n_204),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2401),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2357),
.Y(n_2479)
);

OAI21xp5_ASAP7_75t_SL g2480 ( 
.A1(n_2410),
.A2(n_212),
.B(n_204),
.Y(n_2480)
);

HB1xp67_ASAP7_75t_L g2481 ( 
.A(n_2357),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2377),
.B(n_205),
.Y(n_2482)
);

AND2x2_ASAP7_75t_L g2483 ( 
.A(n_2388),
.B(n_205),
.Y(n_2483)
);

AND2x2_ASAP7_75t_L g2484 ( 
.A(n_2346),
.B(n_206),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2348),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2365),
.Y(n_2486)
);

OAI22xp5_ASAP7_75t_L g2487 ( 
.A1(n_2411),
.A2(n_208),
.B1(n_206),
.B2(n_207),
.Y(n_2487)
);

BUFx3_ASAP7_75t_L g2488 ( 
.A(n_2425),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2349),
.B(n_207),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2429),
.B(n_208),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2343),
.B(n_209),
.Y(n_2491)
);

AND2x2_ASAP7_75t_L g2492 ( 
.A(n_2433),
.B(n_209),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2394),
.B(n_210),
.Y(n_2493)
);

INVxp67_ASAP7_75t_L g2494 ( 
.A(n_2397),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2365),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2365),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2409),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2403),
.Y(n_2498)
);

NOR2xp33_ASAP7_75t_L g2499 ( 
.A(n_2382),
.B(n_211),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2435),
.B(n_212),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2369),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2384),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2400),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_L g2504 ( 
.A(n_2414),
.B(n_213),
.Y(n_2504)
);

OR2x2_ASAP7_75t_L g2505 ( 
.A(n_2358),
.B(n_213),
.Y(n_2505)
);

INVx1_ASAP7_75t_SL g2506 ( 
.A(n_2353),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2383),
.B(n_214),
.Y(n_2507)
);

INVx5_ASAP7_75t_L g2508 ( 
.A(n_2359),
.Y(n_2508)
);

NAND2x1_ASAP7_75t_L g2509 ( 
.A(n_2355),
.B(n_214),
.Y(n_2509)
);

BUFx6f_ASAP7_75t_L g2510 ( 
.A(n_2395),
.Y(n_2510)
);

AND2x2_ASAP7_75t_L g2511 ( 
.A(n_2387),
.B(n_215),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2370),
.B(n_2366),
.Y(n_2512)
);

AOI222xp33_ASAP7_75t_L g2513 ( 
.A1(n_2396),
.A2(n_217),
.B1(n_219),
.B2(n_215),
.C1(n_216),
.C2(n_218),
.Y(n_2513)
);

INVxp67_ASAP7_75t_L g2514 ( 
.A(n_2406),
.Y(n_2514)
);

OR2x2_ASAP7_75t_L g2515 ( 
.A(n_2356),
.B(n_2367),
.Y(n_2515)
);

AND2x4_ASAP7_75t_L g2516 ( 
.A(n_2424),
.B(n_216),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2413),
.Y(n_2517)
);

AND2x4_ASAP7_75t_L g2518 ( 
.A(n_2428),
.B(n_218),
.Y(n_2518)
);

INVx3_ASAP7_75t_L g2519 ( 
.A(n_2417),
.Y(n_2519)
);

BUFx2_ASAP7_75t_L g2520 ( 
.A(n_2399),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2422),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2423),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2426),
.Y(n_2523)
);

NOR2xp33_ASAP7_75t_L g2524 ( 
.A(n_2340),
.B(n_220),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_2418),
.B(n_2419),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2402),
.B(n_220),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2360),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2372),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2379),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2354),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2373),
.B(n_221),
.Y(n_2531)
);

BUFx3_ASAP7_75t_L g2532 ( 
.A(n_2427),
.Y(n_2532)
);

OR2x2_ASAP7_75t_L g2533 ( 
.A(n_2436),
.B(n_221),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2350),
.B(n_222),
.Y(n_2534)
);

NOR2xp33_ASAP7_75t_L g2535 ( 
.A(n_2368),
.B(n_222),
.Y(n_2535)
);

BUFx2_ASAP7_75t_L g2536 ( 
.A(n_2345),
.Y(n_2536)
);

AND2x2_ASAP7_75t_L g2537 ( 
.A(n_2345),
.B(n_223),
.Y(n_2537)
);

OR2x2_ASAP7_75t_L g2538 ( 
.A(n_2389),
.B(n_223),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2342),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2350),
.B(n_224),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2350),
.B(n_224),
.Y(n_2541)
);

AND2x2_ASAP7_75t_L g2542 ( 
.A(n_2345),
.B(n_225),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2342),
.Y(n_2543)
);

HB1xp67_ASAP7_75t_L g2544 ( 
.A(n_2389),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2342),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2350),
.B(n_225),
.Y(n_2546)
);

OR2x2_ASAP7_75t_L g2547 ( 
.A(n_2389),
.B(n_226),
.Y(n_2547)
);

AND2x4_ASAP7_75t_L g2548 ( 
.A(n_2345),
.B(n_226),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2345),
.B(n_227),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2345),
.B(n_227),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2342),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2345),
.B(n_228),
.Y(n_2552)
);

AND2x4_ASAP7_75t_L g2553 ( 
.A(n_2345),
.B(n_229),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2342),
.Y(n_2554)
);

BUFx3_ASAP7_75t_L g2555 ( 
.A(n_2405),
.Y(n_2555)
);

AND2x4_ASAP7_75t_L g2556 ( 
.A(n_2345),
.B(n_230),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2342),
.Y(n_2557)
);

AND2x4_ASAP7_75t_SL g2558 ( 
.A(n_2364),
.B(n_230),
.Y(n_2558)
);

AOI22xp5_ASAP7_75t_L g2559 ( 
.A1(n_2432),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2342),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2502),
.B(n_232),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2443),
.Y(n_2562)
);

INVx4_ASAP7_75t_L g2563 ( 
.A(n_2468),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_L g2564 ( 
.A(n_2501),
.B(n_2472),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2474),
.B(n_2498),
.Y(n_2565)
);

OR2x2_ASAP7_75t_L g2566 ( 
.A(n_2446),
.B(n_2536),
.Y(n_2566)
);

INVxp67_ASAP7_75t_SL g2567 ( 
.A(n_2494),
.Y(n_2567)
);

BUFx2_ASAP7_75t_SL g2568 ( 
.A(n_2555),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_2497),
.B(n_2471),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_SL g2570 ( 
.A(n_2506),
.B(n_233),
.Y(n_2570)
);

AND2x4_ASAP7_75t_L g2571 ( 
.A(n_2475),
.B(n_234),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2437),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2461),
.B(n_234),
.Y(n_2573)
);

NAND3xp33_ASAP7_75t_L g2574 ( 
.A(n_2508),
.B(n_235),
.C(n_236),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2441),
.Y(n_2575)
);

AND2x2_ASAP7_75t_L g2576 ( 
.A(n_2485),
.B(n_236),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2476),
.B(n_237),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2447),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2442),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2459),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2448),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2463),
.B(n_238),
.Y(n_2582)
);

INVx2_ASAP7_75t_SL g2583 ( 
.A(n_2468),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2464),
.B(n_239),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2458),
.Y(n_2585)
);

AND2x2_ASAP7_75t_L g2586 ( 
.A(n_2488),
.B(n_239),
.Y(n_2586)
);

NOR2xp33_ASAP7_75t_L g2587 ( 
.A(n_2440),
.B(n_240),
.Y(n_2587)
);

AOI22xp33_ASAP7_75t_L g2588 ( 
.A1(n_2520),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.Y(n_2588)
);

AND2x2_ASAP7_75t_L g2589 ( 
.A(n_2445),
.B(n_2544),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_2444),
.B(n_241),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2534),
.B(n_243),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2540),
.B(n_244),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2539),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2456),
.B(n_244),
.Y(n_2594)
);

AND2x2_ASAP7_75t_L g2595 ( 
.A(n_2451),
.B(n_245),
.Y(n_2595)
);

AND2x2_ASAP7_75t_L g2596 ( 
.A(n_2479),
.B(n_245),
.Y(n_2596)
);

AND2x2_ASAP7_75t_L g2597 ( 
.A(n_2462),
.B(n_246),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2543),
.Y(n_2598)
);

AOI221xp5_ASAP7_75t_L g2599 ( 
.A1(n_2519),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.C(n_249),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2545),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2551),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2554),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2557),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2560),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2481),
.B(n_247),
.Y(n_2605)
);

NOR2xp33_ASAP7_75t_L g2606 ( 
.A(n_2514),
.B(n_2491),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2541),
.B(n_250),
.Y(n_2607)
);

AND2x4_ASAP7_75t_L g2608 ( 
.A(n_2478),
.B(n_252),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2546),
.B(n_251),
.Y(n_2609)
);

OR2x2_ASAP7_75t_L g2610 ( 
.A(n_2486),
.B(n_251),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2470),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2473),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2452),
.B(n_252),
.Y(n_2613)
);

AND2x2_ASAP7_75t_L g2614 ( 
.A(n_2460),
.B(n_253),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2495),
.Y(n_2615)
);

INVx2_ASAP7_75t_SL g2616 ( 
.A(n_2548),
.Y(n_2616)
);

OR2x2_ASAP7_75t_L g2617 ( 
.A(n_2496),
.B(n_253),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2537),
.B(n_254),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2465),
.Y(n_2619)
);

AND2x2_ASAP7_75t_L g2620 ( 
.A(n_2542),
.B(n_2549),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2505),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2467),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2517),
.B(n_254),
.Y(n_2623)
);

AND2x2_ASAP7_75t_L g2624 ( 
.A(n_2550),
.B(n_255),
.Y(n_2624)
);

AND2x2_ASAP7_75t_L g2625 ( 
.A(n_2552),
.B(n_255),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2538),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2521),
.B(n_256),
.Y(n_2627)
);

HB1xp67_ASAP7_75t_L g2628 ( 
.A(n_2547),
.Y(n_2628)
);

NAND3xp33_ASAP7_75t_L g2629 ( 
.A(n_2508),
.B(n_2499),
.C(n_2527),
.Y(n_2629)
);

AND2x2_ASAP7_75t_L g2630 ( 
.A(n_2449),
.B(n_256),
.Y(n_2630)
);

INVxp67_ASAP7_75t_L g2631 ( 
.A(n_2438),
.Y(n_2631)
);

AND2x2_ASAP7_75t_L g2632 ( 
.A(n_2553),
.B(n_257),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2522),
.B(n_2523),
.Y(n_2633)
);

OAI221xp5_ASAP7_75t_SL g2634 ( 
.A1(n_2515),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.C(n_261),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2493),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2454),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2507),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_2556),
.B(n_2503),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2453),
.Y(n_2639)
);

AND2x2_ASAP7_75t_L g2640 ( 
.A(n_2483),
.B(n_2489),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2529),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2457),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2482),
.Y(n_2643)
);

HB1xp67_ASAP7_75t_L g2644 ( 
.A(n_2484),
.Y(n_2644)
);

NAND4xp25_ASAP7_75t_L g2645 ( 
.A(n_2513),
.B(n_260),
.C(n_258),
.D(n_259),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2528),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2477),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2455),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2532),
.B(n_261),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2490),
.Y(n_2650)
);

HB1xp67_ASAP7_75t_L g2651 ( 
.A(n_2492),
.Y(n_2651)
);

AND2x2_ASAP7_75t_L g2652 ( 
.A(n_2530),
.B(n_262),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2504),
.B(n_262),
.Y(n_2653)
);

INVx4_ASAP7_75t_L g2654 ( 
.A(n_2558),
.Y(n_2654)
);

OR2x2_ASAP7_75t_L g2655 ( 
.A(n_2525),
.B(n_263),
.Y(n_2655)
);

HB1xp67_ASAP7_75t_L g2656 ( 
.A(n_2535),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_SL g2657 ( 
.A(n_2510),
.B(n_264),
.Y(n_2657)
);

AOI22xp33_ASAP7_75t_L g2658 ( 
.A1(n_2510),
.A2(n_266),
.B1(n_264),
.B2(n_265),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2512),
.B(n_2469),
.Y(n_2659)
);

AND2x2_ASAP7_75t_L g2660 ( 
.A(n_2516),
.B(n_2518),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2466),
.B(n_2511),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2500),
.B(n_267),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2524),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2559),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2526),
.B(n_2439),
.Y(n_2665)
);

AND2x4_ASAP7_75t_L g2666 ( 
.A(n_2509),
.B(n_267),
.Y(n_2666)
);

AND2x2_ASAP7_75t_L g2667 ( 
.A(n_2531),
.B(n_268),
.Y(n_2667)
);

AND2x2_ASAP7_75t_L g2668 ( 
.A(n_2533),
.B(n_268),
.Y(n_2668)
);

INVx2_ASAP7_75t_L g2669 ( 
.A(n_2450),
.Y(n_2669)
);

NAND3xp33_ASAP7_75t_L g2670 ( 
.A(n_2480),
.B(n_269),
.C(n_270),
.Y(n_2670)
);

AND2x4_ASAP7_75t_SL g2671 ( 
.A(n_2487),
.B(n_269),
.Y(n_2671)
);

AND2x4_ASAP7_75t_L g2672 ( 
.A(n_2475),
.B(n_270),
.Y(n_2672)
);

OR2x2_ASAP7_75t_L g2673 ( 
.A(n_2472),
.B(n_271),
.Y(n_2673)
);

INVx3_ASAP7_75t_L g2674 ( 
.A(n_2468),
.Y(n_2674)
);

OR2x2_ASAP7_75t_L g2675 ( 
.A(n_2472),
.B(n_271),
.Y(n_2675)
);

BUFx2_ASAP7_75t_L g2676 ( 
.A(n_2443),
.Y(n_2676)
);

AND2x2_ASAP7_75t_L g2677 ( 
.A(n_2443),
.B(n_272),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2443),
.B(n_272),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2502),
.B(n_273),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2502),
.B(n_273),
.Y(n_2680)
);

AND2x4_ASAP7_75t_SL g2681 ( 
.A(n_2462),
.B(n_274),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2443),
.Y(n_2682)
);

AND2x4_ASAP7_75t_L g2683 ( 
.A(n_2475),
.B(n_274),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2437),
.Y(n_2684)
);

NOR2xp33_ASAP7_75t_L g2685 ( 
.A(n_2440),
.B(n_275),
.Y(n_2685)
);

AND2x2_ASAP7_75t_L g2686 ( 
.A(n_2443),
.B(n_276),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2502),
.B(n_277),
.Y(n_2687)
);

INVxp67_ASAP7_75t_SL g2688 ( 
.A(n_2443),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2437),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2437),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2502),
.B(n_278),
.Y(n_2691)
);

AND2x2_ASAP7_75t_L g2692 ( 
.A(n_2443),
.B(n_279),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2502),
.B(n_280),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2502),
.B(n_280),
.Y(n_2694)
);

OR2x2_ASAP7_75t_L g2695 ( 
.A(n_2472),
.B(n_281),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2437),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2443),
.B(n_281),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_2502),
.B(n_282),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2437),
.Y(n_2699)
);

NOR2xp33_ASAP7_75t_L g2700 ( 
.A(n_2440),
.B(n_282),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2443),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2502),
.B(n_283),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2443),
.Y(n_2703)
);

NAND3xp33_ASAP7_75t_L g2704 ( 
.A(n_2508),
.B(n_283),
.C(n_284),
.Y(n_2704)
);

AND2x2_ASAP7_75t_L g2705 ( 
.A(n_2443),
.B(n_284),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2437),
.Y(n_2706)
);

AND2x2_ASAP7_75t_L g2707 ( 
.A(n_2443),
.B(n_285),
.Y(n_2707)
);

AND2x2_ASAP7_75t_L g2708 ( 
.A(n_2443),
.B(n_286),
.Y(n_2708)
);

NOR2xp67_ASAP7_75t_SL g2709 ( 
.A(n_2508),
.B(n_286),
.Y(n_2709)
);

INVx2_ASAP7_75t_L g2710 ( 
.A(n_2443),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2502),
.B(n_287),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2437),
.Y(n_2712)
);

AND2x2_ASAP7_75t_L g2713 ( 
.A(n_2443),
.B(n_287),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2502),
.B(n_288),
.Y(n_2714)
);

AND2x2_ASAP7_75t_L g2715 ( 
.A(n_2443),
.B(n_289),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2437),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2443),
.B(n_289),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_2443),
.B(n_290),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2437),
.Y(n_2719)
);

INVx3_ASAP7_75t_L g2720 ( 
.A(n_2468),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2437),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2437),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2443),
.B(n_291),
.Y(n_2723)
);

AND2x2_ASAP7_75t_L g2724 ( 
.A(n_2443),
.B(n_291),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2443),
.Y(n_2725)
);

AND2x4_ASAP7_75t_L g2726 ( 
.A(n_2475),
.B(n_293),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2502),
.B(n_293),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2437),
.Y(n_2728)
);

OR2x2_ASAP7_75t_L g2729 ( 
.A(n_2472),
.B(n_294),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2443),
.B(n_294),
.Y(n_2730)
);

AOI22xp33_ASAP7_75t_L g2731 ( 
.A1(n_2629),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.Y(n_2731)
);

AOI22xp33_ASAP7_75t_SL g2732 ( 
.A1(n_2648),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.Y(n_2732)
);

BUFx2_ASAP7_75t_L g2733 ( 
.A(n_2563),
.Y(n_2733)
);

OAI31xp33_ASAP7_75t_L g2734 ( 
.A1(n_2574),
.A2(n_300),
.A3(n_298),
.B(n_299),
.Y(n_2734)
);

HB1xp67_ASAP7_75t_L g2735 ( 
.A(n_2676),
.Y(n_2735)
);

INVx1_ASAP7_75t_SL g2736 ( 
.A(n_2568),
.Y(n_2736)
);

AOI33xp33_ASAP7_75t_L g2737 ( 
.A1(n_2621),
.A2(n_300),
.A3(n_303),
.B1(n_298),
.B2(n_299),
.B3(n_302),
.Y(n_2737)
);

BUFx2_ASAP7_75t_L g2738 ( 
.A(n_2674),
.Y(n_2738)
);

NOR2xp33_ASAP7_75t_L g2739 ( 
.A(n_2583),
.B(n_302),
.Y(n_2739)
);

OAI221xp5_ASAP7_75t_SL g2740 ( 
.A1(n_2645),
.A2(n_2599),
.B1(n_2658),
.B2(n_2588),
.C(n_2670),
.Y(n_2740)
);

NAND4xp25_ASAP7_75t_L g2741 ( 
.A(n_2634),
.B(n_306),
.C(n_307),
.D(n_304),
.Y(n_2741)
);

AOI22xp33_ASAP7_75t_L g2742 ( 
.A1(n_2664),
.A2(n_307),
.B1(n_303),
.B2(n_304),
.Y(n_2742)
);

AND2x2_ASAP7_75t_L g2743 ( 
.A(n_2688),
.B(n_308),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2615),
.Y(n_2744)
);

NOR2x1p5_ASAP7_75t_L g2745 ( 
.A(n_2720),
.B(n_308),
.Y(n_2745)
);

AND2x2_ASAP7_75t_L g2746 ( 
.A(n_2637),
.B(n_309),
.Y(n_2746)
);

AOI22xp33_ASAP7_75t_L g2747 ( 
.A1(n_2606),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2676),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2572),
.Y(n_2749)
);

INVx2_ASAP7_75t_SL g2750 ( 
.A(n_2616),
.Y(n_2750)
);

OAI221xp5_ASAP7_75t_SL g2751 ( 
.A1(n_2704),
.A2(n_2653),
.B1(n_2659),
.B2(n_2665),
.C(n_2649),
.Y(n_2751)
);

INVx2_ASAP7_75t_SL g2752 ( 
.A(n_2654),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2575),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2562),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2682),
.Y(n_2755)
);

INVx2_ASAP7_75t_SL g2756 ( 
.A(n_2566),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2701),
.B(n_310),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2703),
.Y(n_2758)
);

AND2x2_ASAP7_75t_L g2759 ( 
.A(n_2710),
.B(n_311),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2656),
.B(n_2635),
.Y(n_2760)
);

AND2x2_ASAP7_75t_L g2761 ( 
.A(n_2725),
.B(n_312),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2641),
.B(n_312),
.Y(n_2762)
);

AOI22xp33_ASAP7_75t_L g2763 ( 
.A1(n_2663),
.A2(n_2669),
.B1(n_2646),
.B2(n_2643),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2578),
.Y(n_2764)
);

OR2x2_ASAP7_75t_L g2765 ( 
.A(n_2569),
.B(n_313),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2581),
.Y(n_2766)
);

OR2x2_ASAP7_75t_L g2767 ( 
.A(n_2564),
.B(n_313),
.Y(n_2767)
);

AOI221xp5_ASAP7_75t_L g2768 ( 
.A1(n_2709),
.A2(n_317),
.B1(n_314),
.B2(n_315),
.C(n_318),
.Y(n_2768)
);

OAI221xp5_ASAP7_75t_L g2769 ( 
.A1(n_2567),
.A2(n_320),
.B1(n_315),
.B2(n_319),
.C(n_321),
.Y(n_2769)
);

INVxp67_ASAP7_75t_SL g2770 ( 
.A(n_2651),
.Y(n_2770)
);

OAI221xp5_ASAP7_75t_L g2771 ( 
.A1(n_2657),
.A2(n_322),
.B1(n_319),
.B2(n_321),
.C(n_323),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2642),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2585),
.Y(n_2773)
);

AO21x2_ASAP7_75t_L g2774 ( 
.A1(n_2605),
.A2(n_323),
.B(n_324),
.Y(n_2774)
);

NOR2xp33_ASAP7_75t_L g2775 ( 
.A(n_2631),
.B(n_2647),
.Y(n_2775)
);

XNOR2x2_ASAP7_75t_L g2776 ( 
.A(n_2570),
.B(n_324),
.Y(n_2776)
);

HB1xp67_ASAP7_75t_L g2777 ( 
.A(n_2589),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2601),
.Y(n_2778)
);

OR2x2_ASAP7_75t_L g2779 ( 
.A(n_2633),
.B(n_325),
.Y(n_2779)
);

AND2x2_ASAP7_75t_L g2780 ( 
.A(n_2644),
.B(n_2628),
.Y(n_2780)
);

BUFx2_ASAP7_75t_L g2781 ( 
.A(n_2608),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2602),
.Y(n_2782)
);

AND2x2_ASAP7_75t_L g2783 ( 
.A(n_2660),
.B(n_325),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_SL g2784 ( 
.A(n_2666),
.B(n_326),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2650),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_2608),
.Y(n_2786)
);

OAI31xp33_ASAP7_75t_L g2787 ( 
.A1(n_2671),
.A2(n_328),
.A3(n_326),
.B(n_327),
.Y(n_2787)
);

OR2x2_ASAP7_75t_L g2788 ( 
.A(n_2639),
.B(n_327),
.Y(n_2788)
);

AOI22xp33_ASAP7_75t_L g2789 ( 
.A1(n_2655),
.A2(n_330),
.B1(n_328),
.B2(n_329),
.Y(n_2789)
);

OR2x2_ASAP7_75t_L g2790 ( 
.A(n_2619),
.B(n_329),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_2638),
.B(n_331),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2604),
.Y(n_2792)
);

HB1xp67_ASAP7_75t_L g2793 ( 
.A(n_2580),
.Y(n_2793)
);

NOR2xp33_ASAP7_75t_L g2794 ( 
.A(n_2561),
.B(n_332),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2626),
.B(n_332),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2579),
.Y(n_2796)
);

AND2x2_ASAP7_75t_L g2797 ( 
.A(n_2622),
.B(n_333),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2611),
.Y(n_2798)
);

AND2x2_ASAP7_75t_L g2799 ( 
.A(n_2636),
.B(n_333),
.Y(n_2799)
);

OAI22xp5_ASAP7_75t_L g2800 ( 
.A1(n_2623),
.A2(n_2627),
.B1(n_2610),
.B2(n_2617),
.Y(n_2800)
);

OAI221xp5_ASAP7_75t_L g2801 ( 
.A1(n_2679),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.C(n_337),
.Y(n_2801)
);

OAI22xp5_ASAP7_75t_L g2802 ( 
.A1(n_2673),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2612),
.Y(n_2803)
);

OAI31xp33_ASAP7_75t_L g2804 ( 
.A1(n_2587),
.A2(n_339),
.A3(n_337),
.B(n_338),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2620),
.B(n_338),
.Y(n_2805)
);

NOR2x1_ASAP7_75t_L g2806 ( 
.A(n_2675),
.B(n_339),
.Y(n_2806)
);

AND2x2_ASAP7_75t_L g2807 ( 
.A(n_2640),
.B(n_340),
.Y(n_2807)
);

INVx2_ASAP7_75t_SL g2808 ( 
.A(n_2595),
.Y(n_2808)
);

NOR2xp67_ASAP7_75t_L g2809 ( 
.A(n_2565),
.B(n_340),
.Y(n_2809)
);

OAI31xp33_ASAP7_75t_L g2810 ( 
.A1(n_2685),
.A2(n_343),
.A3(n_341),
.B(n_342),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2684),
.Y(n_2811)
);

AOI22xp33_ASAP7_75t_L g2812 ( 
.A1(n_2661),
.A2(n_344),
.B1(n_341),
.B2(n_342),
.Y(n_2812)
);

OAI31xp33_ASAP7_75t_L g2813 ( 
.A1(n_2700),
.A2(n_346),
.A3(n_344),
.B(n_345),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2689),
.Y(n_2814)
);

OR2x2_ASAP7_75t_L g2815 ( 
.A(n_2695),
.B(n_345),
.Y(n_2815)
);

AND2x2_ASAP7_75t_L g2816 ( 
.A(n_2677),
.B(n_346),
.Y(n_2816)
);

OAI22xp33_ASAP7_75t_L g2817 ( 
.A1(n_2729),
.A2(n_349),
.B1(n_347),
.B2(n_348),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2690),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2696),
.Y(n_2819)
);

OAI22xp33_ASAP7_75t_L g2820 ( 
.A1(n_2680),
.A2(n_351),
.B1(n_348),
.B2(n_350),
.Y(n_2820)
);

NAND4xp25_ASAP7_75t_L g2821 ( 
.A(n_2687),
.B(n_352),
.C(n_353),
.D(n_351),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2593),
.Y(n_2822)
);

OAI33xp33_ASAP7_75t_L g2823 ( 
.A1(n_2691),
.A2(n_354),
.A3(n_356),
.B1(n_350),
.B2(n_352),
.B3(n_355),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2699),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2706),
.Y(n_2825)
);

INVx3_ASAP7_75t_L g2826 ( 
.A(n_2571),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2596),
.B(n_354),
.Y(n_2827)
);

NOR2xp33_ASAP7_75t_SL g2828 ( 
.A(n_2672),
.B(n_355),
.Y(n_2828)
);

AND2x2_ASAP7_75t_L g2829 ( 
.A(n_2678),
.B(n_356),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2594),
.B(n_2686),
.Y(n_2830)
);

INVx1_ASAP7_75t_SL g2831 ( 
.A(n_2681),
.Y(n_2831)
);

OR2x2_ASAP7_75t_L g2832 ( 
.A(n_2598),
.B(n_357),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2600),
.Y(n_2833)
);

NAND4xp25_ASAP7_75t_L g2834 ( 
.A(n_2693),
.B(n_2698),
.C(n_2702),
.D(n_2694),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2603),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2692),
.B(n_357),
.Y(n_2836)
);

NAND3xp33_ASAP7_75t_L g2837 ( 
.A(n_2711),
.B(n_358),
.C(n_359),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2712),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2716),
.Y(n_2839)
);

OR2x2_ASAP7_75t_L g2840 ( 
.A(n_2719),
.B(n_358),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2697),
.B(n_359),
.Y(n_2841)
);

INVx3_ASAP7_75t_L g2842 ( 
.A(n_2683),
.Y(n_2842)
);

AOI22xp33_ASAP7_75t_L g2843 ( 
.A1(n_2714),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.Y(n_2843)
);

OAI33xp33_ASAP7_75t_L g2844 ( 
.A1(n_2727),
.A2(n_363),
.A3(n_365),
.B1(n_361),
.B2(n_362),
.B3(n_364),
.Y(n_2844)
);

OAI22xp33_ASAP7_75t_L g2845 ( 
.A1(n_2662),
.A2(n_365),
.B1(n_363),
.B2(n_364),
.Y(n_2845)
);

AND2x2_ASAP7_75t_L g2846 ( 
.A(n_2705),
.B(n_366),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2721),
.Y(n_2847)
);

OAI21xp33_ASAP7_75t_L g2848 ( 
.A1(n_2652),
.A2(n_366),
.B(n_367),
.Y(n_2848)
);

AOI31xp33_ASAP7_75t_L g2849 ( 
.A1(n_2730),
.A2(n_369),
.A3(n_367),
.B(n_368),
.Y(n_2849)
);

AOI22xp33_ASAP7_75t_L g2850 ( 
.A1(n_2668),
.A2(n_372),
.B1(n_369),
.B2(n_371),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2722),
.Y(n_2851)
);

NAND3xp33_ASAP7_75t_L g2852 ( 
.A(n_2590),
.B(n_372),
.C(n_373),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2707),
.B(n_373),
.Y(n_2853)
);

NOR2xp33_ASAP7_75t_L g2854 ( 
.A(n_2736),
.B(n_2726),
.Y(n_2854)
);

NOR2xp33_ASAP7_75t_L g2855 ( 
.A(n_2752),
.B(n_2613),
.Y(n_2855)
);

NAND3xp33_ASAP7_75t_L g2856 ( 
.A(n_2734),
.B(n_2592),
.C(n_2591),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2733),
.Y(n_2857)
);

INVxp67_ASAP7_75t_SL g2858 ( 
.A(n_2735),
.Y(n_2858)
);

OR2x2_ASAP7_75t_L g2859 ( 
.A(n_2770),
.B(n_2728),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2738),
.Y(n_2860)
);

AOI22xp5_ASAP7_75t_L g2861 ( 
.A1(n_2741),
.A2(n_2597),
.B1(n_2713),
.B2(n_2708),
.Y(n_2861)
);

AND2x2_ASAP7_75t_L g2862 ( 
.A(n_2842),
.B(n_2715),
.Y(n_2862)
);

AND2x2_ASAP7_75t_L g2863 ( 
.A(n_2842),
.B(n_2717),
.Y(n_2863)
);

HB1xp67_ASAP7_75t_L g2864 ( 
.A(n_2781),
.Y(n_2864)
);

HB1xp67_ASAP7_75t_L g2865 ( 
.A(n_2748),
.Y(n_2865)
);

INVx2_ASAP7_75t_L g2866 ( 
.A(n_2826),
.Y(n_2866)
);

INVxp67_ASAP7_75t_SL g2867 ( 
.A(n_2809),
.Y(n_2867)
);

HB1xp67_ASAP7_75t_L g2868 ( 
.A(n_2777),
.Y(n_2868)
);

OR2x2_ASAP7_75t_L g2869 ( 
.A(n_2760),
.B(n_2607),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2780),
.Y(n_2870)
);

NAND4xp75_ASAP7_75t_L g2871 ( 
.A(n_2806),
.B(n_2718),
.C(n_2724),
.D(n_2723),
.Y(n_2871)
);

AND2x2_ASAP7_75t_L g2872 ( 
.A(n_2808),
.B(n_2586),
.Y(n_2872)
);

INVxp67_ASAP7_75t_L g2873 ( 
.A(n_2776),
.Y(n_2873)
);

INVx1_ASAP7_75t_SL g2874 ( 
.A(n_2831),
.Y(n_2874)
);

INVx2_ASAP7_75t_SL g2875 ( 
.A(n_2745),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2744),
.Y(n_2876)
);

NAND2x1p5_ASAP7_75t_L g2877 ( 
.A(n_2750),
.B(n_2576),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2749),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2786),
.Y(n_2879)
);

AND2x2_ASAP7_75t_L g2880 ( 
.A(n_2772),
.B(n_2756),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2753),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2764),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2774),
.B(n_2667),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2763),
.B(n_2577),
.Y(n_2884)
);

NOR2xp33_ASAP7_75t_L g2885 ( 
.A(n_2751),
.B(n_2609),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2832),
.Y(n_2886)
);

BUFx2_ASAP7_75t_L g2887 ( 
.A(n_2793),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2775),
.B(n_2630),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2754),
.B(n_2618),
.Y(n_2889)
);

INVx4_ASAP7_75t_L g2890 ( 
.A(n_2783),
.Y(n_2890)
);

AND2x2_ASAP7_75t_L g2891 ( 
.A(n_2755),
.B(n_2624),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_2758),
.B(n_2625),
.Y(n_2892)
);

AND2x2_ASAP7_75t_L g2893 ( 
.A(n_2785),
.B(n_2614),
.Y(n_2893)
);

BUFx6f_ASAP7_75t_L g2894 ( 
.A(n_2743),
.Y(n_2894)
);

AND2x2_ASAP7_75t_L g2895 ( 
.A(n_2791),
.B(n_2632),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2766),
.Y(n_2896)
);

OR2x2_ASAP7_75t_L g2897 ( 
.A(n_2834),
.B(n_2573),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2773),
.Y(n_2898)
);

AND2x2_ASAP7_75t_L g2899 ( 
.A(n_2807),
.B(n_2746),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2800),
.B(n_2582),
.Y(n_2900)
);

AND2x2_ASAP7_75t_L g2901 ( 
.A(n_2805),
.B(n_2584),
.Y(n_2901)
);

AND2x2_ASAP7_75t_L g2902 ( 
.A(n_2799),
.B(n_2797),
.Y(n_2902)
);

BUFx3_ASAP7_75t_L g2903 ( 
.A(n_2757),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2778),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2796),
.Y(n_2905)
);

AND2x2_ASAP7_75t_L g2906 ( 
.A(n_2762),
.B(n_2759),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2761),
.B(n_374),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2830),
.B(n_374),
.Y(n_2908)
);

AND2x2_ASAP7_75t_L g2909 ( 
.A(n_2816),
.B(n_375),
.Y(n_2909)
);

OR2x2_ASAP7_75t_L g2910 ( 
.A(n_2765),
.B(n_375),
.Y(n_2910)
);

AND2x2_ASAP7_75t_L g2911 ( 
.A(n_2829),
.B(n_376),
.Y(n_2911)
);

OR2x2_ASAP7_75t_L g2912 ( 
.A(n_2767),
.B(n_376),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2782),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2874),
.B(n_2849),
.Y(n_2914)
);

OR2x2_ASAP7_75t_L g2915 ( 
.A(n_2864),
.B(n_2779),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2887),
.Y(n_2916)
);

INVx1_ASAP7_75t_SL g2917 ( 
.A(n_2887),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2867),
.B(n_2739),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2873),
.B(n_2794),
.Y(n_2919)
);

AND2x2_ASAP7_75t_L g2920 ( 
.A(n_2875),
.B(n_2822),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2894),
.B(n_2795),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2868),
.Y(n_2922)
);

AND2x2_ASAP7_75t_L g2923 ( 
.A(n_2862),
.B(n_2863),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2877),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2858),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2859),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2894),
.B(n_2817),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2860),
.B(n_2845),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2857),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_L g2930 ( 
.A(n_2899),
.B(n_2906),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2865),
.Y(n_2931)
);

AND2x2_ASAP7_75t_L g2932 ( 
.A(n_2854),
.B(n_2833),
.Y(n_2932)
);

AND2x2_ASAP7_75t_L g2933 ( 
.A(n_2890),
.B(n_2835),
.Y(n_2933)
);

AND2x2_ASAP7_75t_L g2934 ( 
.A(n_2902),
.B(n_2836),
.Y(n_2934)
);

OR2x2_ASAP7_75t_L g2935 ( 
.A(n_2883),
.B(n_2788),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2903),
.Y(n_2936)
);

OR4x1_ASAP7_75t_L g2937 ( 
.A(n_2870),
.B(n_2740),
.C(n_2798),
.D(n_2792),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2901),
.B(n_2820),
.Y(n_2938)
);

AND2x2_ASAP7_75t_L g2939 ( 
.A(n_2872),
.B(n_2846),
.Y(n_2939)
);

AND2x2_ASAP7_75t_L g2940 ( 
.A(n_2866),
.B(n_2803),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2895),
.Y(n_2941)
);

OR2x2_ASAP7_75t_L g2942 ( 
.A(n_2897),
.B(n_2790),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2871),
.B(n_2891),
.Y(n_2943)
);

NAND2x1p5_ASAP7_75t_L g2944 ( 
.A(n_2880),
.B(n_2784),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2876),
.Y(n_2945)
);

INVxp67_ASAP7_75t_SL g2946 ( 
.A(n_2944),
.Y(n_2946)
);

AND2x4_ASAP7_75t_L g2947 ( 
.A(n_2923),
.B(n_2892),
.Y(n_2947)
);

OAI211xp5_ASAP7_75t_L g2948 ( 
.A1(n_2919),
.A2(n_2943),
.B(n_2928),
.C(n_2885),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2916),
.Y(n_2949)
);

INVxp67_ASAP7_75t_L g2950 ( 
.A(n_2914),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2917),
.Y(n_2951)
);

AND2x2_ASAP7_75t_L g2952 ( 
.A(n_2934),
.B(n_2893),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2925),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2922),
.Y(n_2954)
);

AO221x1_ASAP7_75t_L g2955 ( 
.A1(n_2931),
.A2(n_2879),
.B1(n_2802),
.B2(n_2881),
.C(n_2878),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2926),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2930),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2915),
.Y(n_2958)
);

AND2x2_ASAP7_75t_L g2959 ( 
.A(n_2939),
.B(n_2855),
.Y(n_2959)
);

AOI22xp33_ASAP7_75t_L g2960 ( 
.A1(n_2924),
.A2(n_2900),
.B1(n_2886),
.B2(n_2856),
.Y(n_2960)
);

AND2x2_ASAP7_75t_L g2961 ( 
.A(n_2920),
.B(n_2889),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_2936),
.B(n_2861),
.Y(n_2962)
);

AND2x2_ASAP7_75t_L g2963 ( 
.A(n_2932),
.B(n_2888),
.Y(n_2963)
);

AOI22xp5_ASAP7_75t_L g2964 ( 
.A1(n_2929),
.A2(n_2884),
.B1(n_2844),
.B2(n_2823),
.Y(n_2964)
);

INVx2_ASAP7_75t_L g2965 ( 
.A(n_2941),
.Y(n_2965)
);

OR2x2_ASAP7_75t_L g2966 ( 
.A(n_2951),
.B(n_2942),
.Y(n_2966)
);

OAI21xp33_ASAP7_75t_L g2967 ( 
.A1(n_2948),
.A2(n_2918),
.B(n_2927),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2958),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2949),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2947),
.B(n_2933),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2952),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2965),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2956),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2946),
.B(n_2940),
.Y(n_2974)
);

OAI32xp33_ASAP7_75t_L g2975 ( 
.A1(n_2950),
.A2(n_2937),
.A3(n_2935),
.B1(n_2938),
.B2(n_2821),
.Y(n_2975)
);

OR2x2_ASAP7_75t_L g2976 ( 
.A(n_2966),
.B(n_2921),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2971),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2968),
.Y(n_2978)
);

OAI221xp5_ASAP7_75t_L g2979 ( 
.A1(n_2967),
.A2(n_2964),
.B1(n_2960),
.B2(n_2962),
.C(n_2954),
.Y(n_2979)
);

AND2x2_ASAP7_75t_L g2980 ( 
.A(n_2970),
.B(n_2959),
.Y(n_2980)
);

A2O1A1Ixp33_ASAP7_75t_L g2981 ( 
.A1(n_2975),
.A2(n_2737),
.B(n_2810),
.C(n_2804),
.Y(n_2981)
);

OR2x2_ASAP7_75t_L g2982 ( 
.A(n_2974),
.B(n_2869),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2972),
.Y(n_2983)
);

NOR4xp25_ASAP7_75t_L g2984 ( 
.A(n_2969),
.B(n_2953),
.C(n_2957),
.D(n_2945),
.Y(n_2984)
);

A2O1A1Ixp33_ASAP7_75t_L g2985 ( 
.A1(n_2981),
.A2(n_2813),
.B(n_2852),
.C(n_2837),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_SL g2986 ( 
.A(n_2980),
.B(n_2963),
.Y(n_2986)
);

NOR2xp33_ASAP7_75t_L g2987 ( 
.A(n_2979),
.B(n_2976),
.Y(n_2987)
);

AOI211xp5_ASAP7_75t_L g2988 ( 
.A1(n_2984),
.A2(n_2801),
.B(n_2769),
.C(n_2973),
.Y(n_2988)
);

OAI211xp5_ASAP7_75t_L g2989 ( 
.A1(n_2977),
.A2(n_2732),
.B(n_2731),
.C(n_2789),
.Y(n_2989)
);

AOI22xp5_ASAP7_75t_L g2990 ( 
.A1(n_2982),
.A2(n_2955),
.B1(n_2961),
.B2(n_2983),
.Y(n_2990)
);

AOI21xp33_ASAP7_75t_L g2991 ( 
.A1(n_2978),
.A2(n_2945),
.B(n_2905),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2980),
.B(n_2882),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_SL g2993 ( 
.A(n_2980),
.B(n_2828),
.Y(n_2993)
);

AOI322xp5_ASAP7_75t_L g2994 ( 
.A1(n_2981),
.A2(n_2848),
.A3(n_2812),
.B1(n_2747),
.B2(n_2850),
.C1(n_2768),
.C2(n_2896),
.Y(n_2994)
);

OR3x1_ASAP7_75t_L g2995 ( 
.A(n_2977),
.B(n_2904),
.C(n_2898),
.Y(n_2995)
);

NAND3xp33_ASAP7_75t_SL g2996 ( 
.A(n_2981),
.B(n_2787),
.C(n_2742),
.Y(n_2996)
);

OAI211xp5_ASAP7_75t_L g2997 ( 
.A1(n_2979),
.A2(n_2843),
.B(n_2771),
.C(n_2908),
.Y(n_2997)
);

AOI211x1_ASAP7_75t_L g2998 ( 
.A1(n_2979),
.A2(n_2913),
.B(n_2814),
.C(n_2818),
.Y(n_2998)
);

AOI221x1_ASAP7_75t_L g2999 ( 
.A1(n_2977),
.A2(n_2827),
.B1(n_2853),
.B2(n_2841),
.C(n_2907),
.Y(n_2999)
);

O2A1O1Ixp5_ASAP7_75t_SL g3000 ( 
.A1(n_2977),
.A2(n_2819),
.B(n_2824),
.C(n_2811),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2980),
.B(n_2909),
.Y(n_3001)
);

NAND4xp25_ASAP7_75t_L g3002 ( 
.A(n_2979),
.B(n_2912),
.C(n_2910),
.D(n_2911),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2988),
.B(n_2985),
.Y(n_3003)
);

AOI211xp5_ASAP7_75t_L g3004 ( 
.A1(n_2996),
.A2(n_2815),
.B(n_2840),
.C(n_2838),
.Y(n_3004)
);

NOR2x1_ASAP7_75t_L g3005 ( 
.A(n_2995),
.B(n_2825),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_3001),
.Y(n_3006)
);

AOI21xp5_ASAP7_75t_L g3007 ( 
.A1(n_2986),
.A2(n_2847),
.B(n_2839),
.Y(n_3007)
);

INVx2_ASAP7_75t_SL g3008 ( 
.A(n_2993),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2994),
.B(n_2987),
.Y(n_3009)
);

NAND4xp25_ASAP7_75t_L g3010 ( 
.A(n_2990),
.B(n_2851),
.C(n_379),
.D(n_377),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2992),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2999),
.B(n_378),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2998),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2991),
.Y(n_3014)
);

AND2x2_ASAP7_75t_L g3015 ( 
.A(n_2989),
.B(n_2997),
.Y(n_3015)
);

AOI22xp5_ASAP7_75t_L g3016 ( 
.A1(n_3002),
.A2(n_381),
.B1(n_378),
.B2(n_380),
.Y(n_3016)
);

OAI21xp5_ASAP7_75t_L g3017 ( 
.A1(n_3000),
.A2(n_380),
.B(n_381),
.Y(n_3017)
);

AOI211xp5_ASAP7_75t_L g3018 ( 
.A1(n_2996),
.A2(n_384),
.B(n_382),
.C(n_383),
.Y(n_3018)
);

INVx2_ASAP7_75t_L g3019 ( 
.A(n_2995),
.Y(n_3019)
);

OAI22xp33_ASAP7_75t_L g3020 ( 
.A1(n_2990),
.A2(n_385),
.B1(n_382),
.B2(n_384),
.Y(n_3020)
);

OAI31xp33_ASAP7_75t_SL g3021 ( 
.A1(n_2996),
.A2(n_387),
.A3(n_385),
.B(n_386),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_2993),
.B(n_386),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_3005),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_SL g3024 ( 
.A(n_3020),
.B(n_388),
.Y(n_3024)
);

AOI22xp5_ASAP7_75t_L g3025 ( 
.A1(n_3008),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_3021),
.B(n_390),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_3022),
.Y(n_3027)
);

OAI21xp5_ASAP7_75t_L g3028 ( 
.A1(n_3009),
.A2(n_391),
.B(n_392),
.Y(n_3028)
);

INVxp67_ASAP7_75t_L g3029 ( 
.A(n_3012),
.Y(n_3029)
);

O2A1O1Ixp33_ASAP7_75t_SL g3030 ( 
.A1(n_3017),
.A2(n_393),
.B(n_391),
.C(n_392),
.Y(n_3030)
);

AOI21xp5_ASAP7_75t_L g3031 ( 
.A1(n_3003),
.A2(n_393),
.B(n_394),
.Y(n_3031)
);

AOI22xp33_ASAP7_75t_L g3032 ( 
.A1(n_3010),
.A2(n_3015),
.B1(n_3006),
.B2(n_3014),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_3019),
.Y(n_3033)
);

OR2x2_ASAP7_75t_L g3034 ( 
.A(n_3013),
.B(n_394),
.Y(n_3034)
);

NOR3xp33_ASAP7_75t_L g3035 ( 
.A(n_3011),
.B(n_395),
.C(n_396),
.Y(n_3035)
);

OAI211xp5_ASAP7_75t_SL g3036 ( 
.A1(n_3018),
.A2(n_397),
.B(n_395),
.C(n_396),
.Y(n_3036)
);

OAI22xp5_ASAP7_75t_L g3037 ( 
.A1(n_3016),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_3004),
.Y(n_3038)
);

CKINVDCx16_ASAP7_75t_R g3039 ( 
.A(n_3007),
.Y(n_3039)
);

AOI21xp33_ASAP7_75t_L g3040 ( 
.A1(n_3008),
.A2(n_398),
.B(n_399),
.Y(n_3040)
);

HB1xp67_ASAP7_75t_L g3041 ( 
.A(n_3005),
.Y(n_3041)
);

O2A1O1Ixp33_ASAP7_75t_L g3042 ( 
.A1(n_3017),
.A2(n_402),
.B(n_400),
.C(n_401),
.Y(n_3042)
);

A2O1A1Ixp33_ASAP7_75t_L g3043 ( 
.A1(n_3017),
.A2(n_402),
.B(n_400),
.C(n_401),
.Y(n_3043)
);

AOI22xp5_ASAP7_75t_L g3044 ( 
.A1(n_3008),
.A2(n_405),
.B1(n_403),
.B2(n_404),
.Y(n_3044)
);

OAI21xp33_ASAP7_75t_L g3045 ( 
.A1(n_3032),
.A2(n_403),
.B(n_404),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_3039),
.B(n_405),
.Y(n_3046)
);

NOR4xp25_ASAP7_75t_L g3047 ( 
.A(n_3023),
.B(n_408),
.C(n_406),
.D(n_407),
.Y(n_3047)
);

INVxp67_ASAP7_75t_SL g3048 ( 
.A(n_3041),
.Y(n_3048)
);

AOI221xp5_ASAP7_75t_L g3049 ( 
.A1(n_3030),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.C(n_410),
.Y(n_3049)
);

A2O1A1Ixp33_ASAP7_75t_L g3050 ( 
.A1(n_3042),
.A2(n_412),
.B(n_410),
.C(n_411),
.Y(n_3050)
);

AOI221xp5_ASAP7_75t_L g3051 ( 
.A1(n_3028),
.A2(n_414),
.B1(n_411),
.B2(n_413),
.C(n_415),
.Y(n_3051)
);

AND2x2_ASAP7_75t_L g3052 ( 
.A(n_3029),
.B(n_413),
.Y(n_3052)
);

XNOR2xp5_ASAP7_75t_L g3053 ( 
.A(n_3025),
.B(n_414),
.Y(n_3053)
);

INVxp67_ASAP7_75t_L g3054 ( 
.A(n_3026),
.Y(n_3054)
);

O2A1O1Ixp33_ASAP7_75t_L g3055 ( 
.A1(n_3043),
.A2(n_418),
.B(n_416),
.C(n_417),
.Y(n_3055)
);

HB1xp67_ASAP7_75t_L g3056 ( 
.A(n_3034),
.Y(n_3056)
);

AOI22xp5_ASAP7_75t_L g3057 ( 
.A1(n_3033),
.A2(n_418),
.B1(n_416),
.B2(n_417),
.Y(n_3057)
);

NOR2x1_ASAP7_75t_L g3058 ( 
.A(n_3036),
.B(n_419),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_3044),
.Y(n_3059)
);

NOR4xp25_ASAP7_75t_L g3060 ( 
.A(n_3038),
.B(n_421),
.C(n_419),
.D(n_420),
.Y(n_3060)
);

AOI21xp5_ASAP7_75t_L g3061 ( 
.A1(n_3024),
.A2(n_3031),
.B(n_3040),
.Y(n_3061)
);

AOI321xp33_ASAP7_75t_L g3062 ( 
.A1(n_3027),
.A2(n_423),
.A3(n_425),
.B1(n_421),
.B2(n_422),
.C(n_424),
.Y(n_3062)
);

NAND2xp33_ASAP7_75t_SL g3063 ( 
.A(n_3037),
.B(n_422),
.Y(n_3063)
);

OAI221xp5_ASAP7_75t_L g3064 ( 
.A1(n_3035),
.A2(n_427),
.B1(n_424),
.B2(n_425),
.C(n_428),
.Y(n_3064)
);

O2A1O1Ixp33_ASAP7_75t_L g3065 ( 
.A1(n_3041),
.A2(n_429),
.B(n_427),
.C(n_428),
.Y(n_3065)
);

NAND4xp25_ASAP7_75t_L g3066 ( 
.A(n_3032),
.B(n_432),
.C(n_430),
.D(n_431),
.Y(n_3066)
);

OAI22xp33_ASAP7_75t_L g3067 ( 
.A1(n_3039),
.A2(n_432),
.B1(n_430),
.B2(n_431),
.Y(n_3067)
);

AOI221xp5_ASAP7_75t_L g3068 ( 
.A1(n_3030),
.A2(n_435),
.B1(n_433),
.B2(n_434),
.C(n_436),
.Y(n_3068)
);

INVx2_ASAP7_75t_SL g3069 ( 
.A(n_3041),
.Y(n_3069)
);

XNOR2x1_ASAP7_75t_L g3070 ( 
.A(n_3028),
.B(n_433),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_3041),
.Y(n_3071)
);

INVx2_ASAP7_75t_L g3072 ( 
.A(n_3023),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_3041),
.Y(n_3073)
);

AOI211xp5_ASAP7_75t_SL g3074 ( 
.A1(n_3030),
.A2(n_437),
.B(n_434),
.C(n_435),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_3039),
.B(n_437),
.Y(n_3075)
);

AOI321xp33_ASAP7_75t_L g3076 ( 
.A1(n_3032),
.A2(n_440),
.A3(n_442),
.B1(n_438),
.B2(n_439),
.C(n_441),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_3041),
.Y(n_3077)
);

AOI221x1_ASAP7_75t_L g3078 ( 
.A1(n_3040),
.A2(n_441),
.B1(n_439),
.B2(n_440),
.C(n_443),
.Y(n_3078)
);

NOR2x1_ASAP7_75t_L g3079 ( 
.A(n_3023),
.B(n_443),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_3041),
.Y(n_3080)
);

NAND4xp75_ASAP7_75t_L g3081 ( 
.A(n_3028),
.B(n_446),
.C(n_444),
.D(n_445),
.Y(n_3081)
);

A2O1A1Ixp33_ASAP7_75t_L g3082 ( 
.A1(n_3042),
.A2(n_446),
.B(n_444),
.C(n_445),
.Y(n_3082)
);

AOI22xp5_ASAP7_75t_L g3083 ( 
.A1(n_3033),
.A2(n_450),
.B1(n_447),
.B2(n_448),
.Y(n_3083)
);

NOR2x1_ASAP7_75t_L g3084 ( 
.A(n_3079),
.B(n_447),
.Y(n_3084)
);

NOR2x1_ASAP7_75t_L g3085 ( 
.A(n_3066),
.B(n_448),
.Y(n_3085)
);

NOR2x1p5_ASAP7_75t_L g3086 ( 
.A(n_3081),
.B(n_451),
.Y(n_3086)
);

NOR2xp67_ASAP7_75t_L g3087 ( 
.A(n_3069),
.B(n_451),
.Y(n_3087)
);

OR2x2_ASAP7_75t_L g3088 ( 
.A(n_3060),
.B(n_452),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_3046),
.Y(n_3089)
);

AND2x2_ASAP7_75t_L g3090 ( 
.A(n_3058),
.B(n_452),
.Y(n_3090)
);

NOR2xp67_ASAP7_75t_L g3091 ( 
.A(n_3056),
.B(n_453),
.Y(n_3091)
);

AOI22xp5_ASAP7_75t_L g3092 ( 
.A1(n_3045),
.A2(n_3048),
.B1(n_3059),
.B2(n_3071),
.Y(n_3092)
);

AND2x2_ASAP7_75t_L g3093 ( 
.A(n_3052),
.B(n_454),
.Y(n_3093)
);

NOR2x1_ASAP7_75t_L g3094 ( 
.A(n_3067),
.B(n_454),
.Y(n_3094)
);

AND2x2_ASAP7_75t_L g3095 ( 
.A(n_3074),
.B(n_455),
.Y(n_3095)
);

OA22x2_ASAP7_75t_L g3096 ( 
.A1(n_3073),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.Y(n_3096)
);

AND2x4_ASAP7_75t_L g3097 ( 
.A(n_3077),
.B(n_457),
.Y(n_3097)
);

INVx1_ASAP7_75t_SL g3098 ( 
.A(n_3075),
.Y(n_3098)
);

AND2x2_ASAP7_75t_L g3099 ( 
.A(n_3054),
.B(n_458),
.Y(n_3099)
);

INVxp67_ASAP7_75t_SL g3100 ( 
.A(n_3065),
.Y(n_3100)
);

AOI22xp5_ASAP7_75t_L g3101 ( 
.A1(n_3080),
.A2(n_460),
.B1(n_458),
.B2(n_459),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_3072),
.Y(n_3102)
);

AND2x4_ASAP7_75t_L g3103 ( 
.A(n_3078),
.B(n_459),
.Y(n_3103)
);

NOR2x1_ASAP7_75t_L g3104 ( 
.A(n_3070),
.B(n_461),
.Y(n_3104)
);

NOR2xp67_ASAP7_75t_L g3105 ( 
.A(n_3064),
.B(n_462),
.Y(n_3105)
);

AO22x2_ASAP7_75t_L g3106 ( 
.A1(n_3061),
.A2(n_464),
.B1(n_462),
.B2(n_463),
.Y(n_3106)
);

NOR2x1_ASAP7_75t_L g3107 ( 
.A(n_3050),
.B(n_464),
.Y(n_3107)
);

NOR2xp33_ASAP7_75t_L g3108 ( 
.A(n_3082),
.B(n_465),
.Y(n_3108)
);

HB1xp67_ASAP7_75t_L g3109 ( 
.A(n_3047),
.Y(n_3109)
);

AOI22xp5_ASAP7_75t_L g3110 ( 
.A1(n_3063),
.A2(n_467),
.B1(n_465),
.B2(n_466),
.Y(n_3110)
);

AND2x2_ASAP7_75t_L g3111 ( 
.A(n_3049),
.B(n_467),
.Y(n_3111)
);

AND2x2_ASAP7_75t_L g3112 ( 
.A(n_3068),
.B(n_468),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_3053),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_3076),
.Y(n_3114)
);

INVx2_ASAP7_75t_L g3115 ( 
.A(n_3057),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_3062),
.Y(n_3116)
);

NOR2x1_ASAP7_75t_L g3117 ( 
.A(n_3055),
.B(n_468),
.Y(n_3117)
);

NOR2x1_ASAP7_75t_L g3118 ( 
.A(n_3051),
.B(n_469),
.Y(n_3118)
);

AND2x4_ASAP7_75t_L g3119 ( 
.A(n_3083),
.B(n_469),
.Y(n_3119)
);

INVxp33_ASAP7_75t_SL g3120 ( 
.A(n_3056),
.Y(n_3120)
);

NOR2x1_ASAP7_75t_L g3121 ( 
.A(n_3079),
.B(n_470),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_3046),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_3046),
.Y(n_3123)
);

AOI22xp5_ASAP7_75t_L g3124 ( 
.A1(n_3069),
.A2(n_472),
.B1(n_470),
.B2(n_471),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_3046),
.Y(n_3125)
);

INVxp33_ASAP7_75t_SL g3126 ( 
.A(n_3056),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_3046),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_3046),
.Y(n_3128)
);

NAND2x1_ASAP7_75t_L g3129 ( 
.A(n_3079),
.B(n_471),
.Y(n_3129)
);

OAI211xp5_ASAP7_75t_SL g3130 ( 
.A1(n_3054),
.A2(n_474),
.B(n_472),
.C(n_473),
.Y(n_3130)
);

INVxp67_ASAP7_75t_SL g3131 ( 
.A(n_3079),
.Y(n_3131)
);

AND3x2_ASAP7_75t_L g3132 ( 
.A(n_3109),
.B(n_473),
.C(n_475),
.Y(n_3132)
);

AND2x4_ASAP7_75t_L g3133 ( 
.A(n_3087),
.B(n_475),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_3096),
.Y(n_3134)
);

AO22x2_ASAP7_75t_L g3135 ( 
.A1(n_3131),
.A2(n_478),
.B1(n_476),
.B2(n_477),
.Y(n_3135)
);

HB1xp67_ASAP7_75t_L g3136 ( 
.A(n_3091),
.Y(n_3136)
);

NOR2x1_ASAP7_75t_L g3137 ( 
.A(n_3084),
.B(n_476),
.Y(n_3137)
);

XNOR2x1_ASAP7_75t_L g3138 ( 
.A(n_3086),
.B(n_477),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_3106),
.Y(n_3139)
);

AND2x4_ASAP7_75t_L g3140 ( 
.A(n_3102),
.B(n_479),
.Y(n_3140)
);

NOR3xp33_ASAP7_75t_L g3141 ( 
.A(n_3100),
.B(n_480),
.C(n_481),
.Y(n_3141)
);

AND3x2_ASAP7_75t_L g3142 ( 
.A(n_3095),
.B(n_480),
.C(n_481),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_3097),
.B(n_482),
.Y(n_3143)
);

NAND4xp75_ASAP7_75t_L g3144 ( 
.A(n_3121),
.B(n_484),
.C(n_482),
.D(n_483),
.Y(n_3144)
);

NOR2x1_ASAP7_75t_L g3145 ( 
.A(n_3129),
.B(n_3104),
.Y(n_3145)
);

XNOR2xp5_ASAP7_75t_L g3146 ( 
.A(n_3092),
.B(n_483),
.Y(n_3146)
);

AND2x2_ASAP7_75t_L g3147 ( 
.A(n_3090),
.B(n_485),
.Y(n_3147)
);

NOR2x1_ASAP7_75t_L g3148 ( 
.A(n_3103),
.B(n_486),
.Y(n_3148)
);

OAI21xp33_ASAP7_75t_L g3149 ( 
.A1(n_3120),
.A2(n_487),
.B(n_488),
.Y(n_3149)
);

OR2x2_ASAP7_75t_L g3150 ( 
.A(n_3088),
.B(n_488),
.Y(n_3150)
);

INVxp67_ASAP7_75t_SL g3151 ( 
.A(n_3094),
.Y(n_3151)
);

AOI22xp5_ASAP7_75t_L g3152 ( 
.A1(n_3126),
.A2(n_491),
.B1(n_489),
.B2(n_490),
.Y(n_3152)
);

INVx2_ASAP7_75t_L g3153 ( 
.A(n_3106),
.Y(n_3153)
);

AOI22xp5_ASAP7_75t_L g3154 ( 
.A1(n_3116),
.A2(n_491),
.B1(n_489),
.B2(n_490),
.Y(n_3154)
);

OR2x2_ASAP7_75t_L g3155 ( 
.A(n_3114),
.B(n_492),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3093),
.Y(n_3156)
);

OAI322xp33_ASAP7_75t_L g3157 ( 
.A1(n_3113),
.A2(n_497),
.A3(n_496),
.B1(n_494),
.B2(n_492),
.C1(n_493),
.C2(n_495),
.Y(n_3157)
);

AOI22xp5_ASAP7_75t_L g3158 ( 
.A1(n_3085),
.A2(n_496),
.B1(n_493),
.B2(n_494),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_3099),
.Y(n_3159)
);

INVx3_ASAP7_75t_L g3160 ( 
.A(n_3119),
.Y(n_3160)
);

AND2x4_ASAP7_75t_L g3161 ( 
.A(n_3089),
.B(n_497),
.Y(n_3161)
);

INVx2_ASAP7_75t_SL g3162 ( 
.A(n_3107),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_3111),
.Y(n_3163)
);

NAND4xp75_ASAP7_75t_L g3164 ( 
.A(n_3117),
.B(n_500),
.C(n_498),
.D(n_499),
.Y(n_3164)
);

XNOR2xp5_ASAP7_75t_L g3165 ( 
.A(n_3110),
.B(n_3124),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_3112),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_3115),
.Y(n_3167)
);

NOR2xp33_ASAP7_75t_L g3168 ( 
.A(n_3130),
.B(n_498),
.Y(n_3168)
);

NOR3xp33_ASAP7_75t_SL g3169 ( 
.A(n_3108),
.B(n_500),
.C(n_501),
.Y(n_3169)
);

NAND4xp25_ASAP7_75t_L g3170 ( 
.A(n_3105),
.B(n_503),
.C(n_501),
.D(n_502),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_3101),
.B(n_502),
.Y(n_3171)
);

NAND4xp75_ASAP7_75t_L g3172 ( 
.A(n_3118),
.B(n_505),
.C(n_503),
.D(n_504),
.Y(n_3172)
);

OAI21xp5_ASAP7_75t_L g3173 ( 
.A1(n_3098),
.A2(n_505),
.B(n_506),
.Y(n_3173)
);

NOR2xp33_ASAP7_75t_SL g3174 ( 
.A(n_3122),
.B(n_506),
.Y(n_3174)
);

OAI221xp5_ASAP7_75t_L g3175 ( 
.A1(n_3123),
.A2(n_509),
.B1(n_507),
.B2(n_508),
.C(n_510),
.Y(n_3175)
);

NOR2x1_ASAP7_75t_L g3176 ( 
.A(n_3125),
.B(n_508),
.Y(n_3176)
);

NAND4xp75_ASAP7_75t_L g3177 ( 
.A(n_3127),
.B(n_512),
.C(n_510),
.D(n_511),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_3128),
.Y(n_3178)
);

INVxp67_ASAP7_75t_L g3179 ( 
.A(n_3084),
.Y(n_3179)
);

AND2x4_ASAP7_75t_L g3180 ( 
.A(n_3087),
.B(n_512),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_3096),
.Y(n_3181)
);

OAI22xp5_ASAP7_75t_L g3182 ( 
.A1(n_3092),
.A2(n_515),
.B1(n_513),
.B2(n_514),
.Y(n_3182)
);

BUFx2_ASAP7_75t_L g3183 ( 
.A(n_3084),
.Y(n_3183)
);

NOR2x1_ASAP7_75t_L g3184 ( 
.A(n_3084),
.B(n_513),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_3096),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_3106),
.Y(n_3186)
);

OR2x2_ASAP7_75t_L g3187 ( 
.A(n_3088),
.B(n_514),
.Y(n_3187)
);

NAND4xp75_ASAP7_75t_L g3188 ( 
.A(n_3084),
.B(n_518),
.C(n_516),
.D(n_517),
.Y(n_3188)
);

AOI22xp5_ASAP7_75t_L g3189 ( 
.A1(n_3120),
.A2(n_518),
.B1(n_516),
.B2(n_517),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_3096),
.Y(n_3190)
);

AND4x1_ASAP7_75t_L g3191 ( 
.A(n_3092),
.B(n_521),
.C(n_519),
.D(n_520),
.Y(n_3191)
);

AND2x4_ASAP7_75t_L g3192 ( 
.A(n_3087),
.B(n_519),
.Y(n_3192)
);

AOI321xp33_ASAP7_75t_L g3193 ( 
.A1(n_3151),
.A2(n_522),
.A3(n_524),
.B1(n_520),
.B2(n_521),
.C(n_523),
.Y(n_3193)
);

INVxp67_ASAP7_75t_SL g3194 ( 
.A(n_3137),
.Y(n_3194)
);

NAND5xp2_ASAP7_75t_L g3195 ( 
.A(n_3134),
.B(n_525),
.C(n_522),
.D(n_523),
.E(n_526),
.Y(n_3195)
);

AOI211xp5_ASAP7_75t_L g3196 ( 
.A1(n_3170),
.A2(n_528),
.B(n_526),
.C(n_527),
.Y(n_3196)
);

OAI21xp5_ASAP7_75t_L g3197 ( 
.A1(n_3148),
.A2(n_3179),
.B(n_3146),
.Y(n_3197)
);

A2O1A1Ixp33_ASAP7_75t_L g3198 ( 
.A1(n_3168),
.A2(n_529),
.B(n_527),
.C(n_528),
.Y(n_3198)
);

HB1xp67_ASAP7_75t_L g3199 ( 
.A(n_3135),
.Y(n_3199)
);

OAI211xp5_ASAP7_75t_SL g3200 ( 
.A1(n_3145),
.A2(n_531),
.B(n_529),
.C(n_530),
.Y(n_3200)
);

AO22x2_ASAP7_75t_L g3201 ( 
.A1(n_3139),
.A2(n_533),
.B1(n_531),
.B2(n_532),
.Y(n_3201)
);

AOI211xp5_ASAP7_75t_L g3202 ( 
.A1(n_3182),
.A2(n_535),
.B(n_532),
.C(n_534),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_3133),
.Y(n_3203)
);

AOI221x1_ASAP7_75t_L g3204 ( 
.A1(n_3141),
.A2(n_3186),
.B1(n_3153),
.B2(n_3185),
.C(n_3181),
.Y(n_3204)
);

OAI311xp33_ASAP7_75t_L g3205 ( 
.A1(n_3190),
.A2(n_537),
.A3(n_534),
.B1(n_536),
.C1(n_539),
.Y(n_3205)
);

OAI211xp5_ASAP7_75t_L g3206 ( 
.A1(n_3158),
.A2(n_539),
.B(n_536),
.C(n_537),
.Y(n_3206)
);

AOI22xp5_ASAP7_75t_L g3207 ( 
.A1(n_3167),
.A2(n_542),
.B1(n_540),
.B2(n_541),
.Y(n_3207)
);

OAI221xp5_ASAP7_75t_L g3208 ( 
.A1(n_3162),
.A2(n_3183),
.B1(n_3184),
.B2(n_3155),
.C(n_3136),
.Y(n_3208)
);

AOI22xp5_ASAP7_75t_L g3209 ( 
.A1(n_3156),
.A2(n_542),
.B1(n_540),
.B2(n_541),
.Y(n_3209)
);

NOR2xp33_ASAP7_75t_L g3210 ( 
.A(n_3191),
.B(n_3149),
.Y(n_3210)
);

AOI221xp5_ASAP7_75t_L g3211 ( 
.A1(n_3178),
.A2(n_3163),
.B1(n_3166),
.B2(n_3160),
.C(n_3147),
.Y(n_3211)
);

AOI21xp5_ASAP7_75t_L g3212 ( 
.A1(n_3138),
.A2(n_543),
.B(n_544),
.Y(n_3212)
);

OAI211xp5_ASAP7_75t_SL g3213 ( 
.A1(n_3169),
.A2(n_545),
.B(n_543),
.C(n_544),
.Y(n_3213)
);

OAI211xp5_ASAP7_75t_L g3214 ( 
.A1(n_3176),
.A2(n_547),
.B(n_545),
.C(n_546),
.Y(n_3214)
);

CKINVDCx20_ASAP7_75t_R g3215 ( 
.A(n_3165),
.Y(n_3215)
);

OAI211xp5_ASAP7_75t_L g3216 ( 
.A1(n_3171),
.A2(n_548),
.B(n_546),
.C(n_547),
.Y(n_3216)
);

OAI211xp5_ASAP7_75t_SL g3217 ( 
.A1(n_3159),
.A2(n_552),
.B(n_549),
.C(n_551),
.Y(n_3217)
);

NOR2xp67_ASAP7_75t_L g3218 ( 
.A(n_3180),
.B(n_549),
.Y(n_3218)
);

NOR2x1_ASAP7_75t_L g3219 ( 
.A(n_3144),
.B(n_3188),
.Y(n_3219)
);

NAND4xp75_ASAP7_75t_L g3220 ( 
.A(n_3173),
.B(n_554),
.C(n_551),
.D(n_553),
.Y(n_3220)
);

AND2x4_ASAP7_75t_L g3221 ( 
.A(n_3192),
.B(n_553),
.Y(n_3221)
);

AOI222xp33_ASAP7_75t_L g3222 ( 
.A1(n_3143),
.A2(n_556),
.B1(n_558),
.B2(n_554),
.C1(n_555),
.C2(n_557),
.Y(n_3222)
);

OAI221xp5_ASAP7_75t_L g3223 ( 
.A1(n_3150),
.A2(n_558),
.B1(n_555),
.B2(n_557),
.C(n_559),
.Y(n_3223)
);

NOR2xp67_ASAP7_75t_L g3224 ( 
.A(n_3154),
.B(n_559),
.Y(n_3224)
);

OAI21xp33_ASAP7_75t_SL g3225 ( 
.A1(n_3172),
.A2(n_3164),
.B(n_3187),
.Y(n_3225)
);

AOI22x1_ASAP7_75t_L g3226 ( 
.A1(n_3135),
.A2(n_562),
.B1(n_560),
.B2(n_561),
.Y(n_3226)
);

OAI221xp5_ASAP7_75t_L g3227 ( 
.A1(n_3174),
.A2(n_562),
.B1(n_560),
.B2(n_561),
.C(n_563),
.Y(n_3227)
);

OAI22x1_ASAP7_75t_L g3228 ( 
.A1(n_3152),
.A2(n_565),
.B1(n_563),
.B2(n_564),
.Y(n_3228)
);

OAI211xp5_ASAP7_75t_L g3229 ( 
.A1(n_3189),
.A2(n_566),
.B(n_564),
.C(n_565),
.Y(n_3229)
);

INVx1_ASAP7_75t_SL g3230 ( 
.A(n_3132),
.Y(n_3230)
);

AO22x2_ASAP7_75t_L g3231 ( 
.A1(n_3177),
.A2(n_568),
.B1(n_566),
.B2(n_567),
.Y(n_3231)
);

AO22x2_ASAP7_75t_L g3232 ( 
.A1(n_3140),
.A2(n_569),
.B1(n_567),
.B2(n_568),
.Y(n_3232)
);

OA22x2_ASAP7_75t_L g3233 ( 
.A1(n_3142),
.A2(n_571),
.B1(n_569),
.B2(n_570),
.Y(n_3233)
);

AOI221xp5_ASAP7_75t_L g3234 ( 
.A1(n_3157),
.A2(n_572),
.B1(n_570),
.B2(n_571),
.C(n_573),
.Y(n_3234)
);

AND4x1_ASAP7_75t_L g3235 ( 
.A(n_3175),
.B(n_576),
.C(n_572),
.D(n_575),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_L g3236 ( 
.A(n_3161),
.B(n_575),
.Y(n_3236)
);

XNOR2xp5_ASAP7_75t_L g3237 ( 
.A(n_3191),
.B(n_576),
.Y(n_3237)
);

AOI211xp5_ASAP7_75t_L g3238 ( 
.A1(n_3170),
.A2(n_579),
.B(n_577),
.C(n_578),
.Y(n_3238)
);

OAI211xp5_ASAP7_75t_SL g3239 ( 
.A1(n_3179),
.A2(n_579),
.B(n_577),
.C(n_578),
.Y(n_3239)
);

AOI22xp5_ASAP7_75t_L g3240 ( 
.A1(n_3134),
.A2(n_582),
.B1(n_580),
.B2(n_581),
.Y(n_3240)
);

A2O1A1Ixp33_ASAP7_75t_L g3241 ( 
.A1(n_3168),
.A2(n_584),
.B(n_580),
.C(n_583),
.Y(n_3241)
);

AOI22xp5_ASAP7_75t_L g3242 ( 
.A1(n_3134),
.A2(n_585),
.B1(n_583),
.B2(n_584),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_3132),
.B(n_585),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_3133),
.Y(n_3244)
);

AOI21xp33_ASAP7_75t_SL g3245 ( 
.A1(n_3139),
.A2(n_586),
.B(n_587),
.Y(n_3245)
);

NOR2x1_ASAP7_75t_L g3246 ( 
.A(n_3148),
.B(n_586),
.Y(n_3246)
);

NAND5xp2_ASAP7_75t_L g3247 ( 
.A(n_3134),
.B(n_589),
.C(n_587),
.D(n_588),
.E(n_590),
.Y(n_3247)
);

AND2x4_ASAP7_75t_L g3248 ( 
.A(n_3218),
.B(n_588),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_3199),
.B(n_589),
.Y(n_3249)
);

AND2x2_ASAP7_75t_L g3250 ( 
.A(n_3219),
.B(n_590),
.Y(n_3250)
);

OAI22xp5_ASAP7_75t_L g3251 ( 
.A1(n_3215),
.A2(n_593),
.B1(n_591),
.B2(n_592),
.Y(n_3251)
);

XOR2x2_ASAP7_75t_L g3252 ( 
.A(n_3237),
.B(n_592),
.Y(n_3252)
);

AOI21xp5_ASAP7_75t_L g3253 ( 
.A1(n_3194),
.A2(n_594),
.B(n_595),
.Y(n_3253)
);

AND3x1_ASAP7_75t_L g3254 ( 
.A(n_3196),
.B(n_594),
.C(n_596),
.Y(n_3254)
);

AND3x2_ASAP7_75t_L g3255 ( 
.A(n_3221),
.B(n_596),
.C(n_597),
.Y(n_3255)
);

HB1xp67_ASAP7_75t_L g3256 ( 
.A(n_3201),
.Y(n_3256)
);

INVx2_ASAP7_75t_SL g3257 ( 
.A(n_3246),
.Y(n_3257)
);

AO22x2_ASAP7_75t_L g3258 ( 
.A1(n_3230),
.A2(n_599),
.B1(n_597),
.B2(n_598),
.Y(n_3258)
);

INVx4_ASAP7_75t_L g3259 ( 
.A(n_3203),
.Y(n_3259)
);

AND2x2_ASAP7_75t_L g3260 ( 
.A(n_3244),
.B(n_598),
.Y(n_3260)
);

OAI22xp5_ASAP7_75t_SL g3261 ( 
.A1(n_3208),
.A2(n_603),
.B1(n_599),
.B2(n_601),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3233),
.Y(n_3262)
);

NOR2x1_ASAP7_75t_L g3263 ( 
.A(n_3243),
.B(n_601),
.Y(n_3263)
);

OR2x2_ASAP7_75t_L g3264 ( 
.A(n_3195),
.B(n_603),
.Y(n_3264)
);

CKINVDCx5p33_ASAP7_75t_R g3265 ( 
.A(n_3197),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_SL g3266 ( 
.A(n_3193),
.B(n_3245),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_3226),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_3240),
.B(n_604),
.Y(n_3268)
);

AOI22x1_ASAP7_75t_L g3269 ( 
.A1(n_3231),
.A2(n_606),
.B1(n_604),
.B2(n_605),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_3242),
.B(n_605),
.Y(n_3270)
);

XNOR2xp5_ASAP7_75t_L g3271 ( 
.A(n_3235),
.B(n_606),
.Y(n_3271)
);

CKINVDCx5p33_ASAP7_75t_R g3272 ( 
.A(n_3210),
.Y(n_3272)
);

INVx2_ASAP7_75t_SL g3273 ( 
.A(n_3231),
.Y(n_3273)
);

XOR2x2_ASAP7_75t_L g3274 ( 
.A(n_3220),
.B(n_607),
.Y(n_3274)
);

AND2x4_ASAP7_75t_L g3275 ( 
.A(n_3204),
.B(n_607),
.Y(n_3275)
);

HB1xp67_ASAP7_75t_L g3276 ( 
.A(n_3201),
.Y(n_3276)
);

INVx3_ASAP7_75t_L g3277 ( 
.A(n_3232),
.Y(n_3277)
);

AND4x1_ASAP7_75t_L g3278 ( 
.A(n_3211),
.B(n_610),
.C(n_608),
.D(n_609),
.Y(n_3278)
);

AND2x2_ASAP7_75t_L g3279 ( 
.A(n_3238),
.B(n_608),
.Y(n_3279)
);

NOR2xp33_ASAP7_75t_L g3280 ( 
.A(n_3247),
.B(n_610),
.Y(n_3280)
);

OR2x2_ASAP7_75t_L g3281 ( 
.A(n_3236),
.B(n_611),
.Y(n_3281)
);

OAI22xp5_ASAP7_75t_SL g3282 ( 
.A1(n_3227),
.A2(n_613),
.B1(n_611),
.B2(n_612),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_3232),
.B(n_612),
.Y(n_3283)
);

OR2x2_ASAP7_75t_L g3284 ( 
.A(n_3198),
.B(n_3241),
.Y(n_3284)
);

NOR3xp33_ASAP7_75t_SL g3285 ( 
.A(n_3225),
.B(n_613),
.C(n_614),
.Y(n_3285)
);

NOR3xp33_ASAP7_75t_L g3286 ( 
.A(n_3216),
.B(n_614),
.C(n_615),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_3214),
.Y(n_3287)
);

XNOR2xp5_ASAP7_75t_L g3288 ( 
.A(n_3228),
.B(n_3202),
.Y(n_3288)
);

HB1xp67_ASAP7_75t_L g3289 ( 
.A(n_3256),
.Y(n_3289)
);

AOI22xp5_ASAP7_75t_L g3290 ( 
.A1(n_3280),
.A2(n_3213),
.B1(n_3200),
.B2(n_3217),
.Y(n_3290)
);

OR2x2_ASAP7_75t_L g3291 ( 
.A(n_3264),
.B(n_3229),
.Y(n_3291)
);

NAND2x1_ASAP7_75t_L g3292 ( 
.A(n_3248),
.B(n_3224),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_3255),
.B(n_3234),
.Y(n_3293)
);

INVx2_ASAP7_75t_L g3294 ( 
.A(n_3258),
.Y(n_3294)
);

INVx2_ASAP7_75t_L g3295 ( 
.A(n_3258),
.Y(n_3295)
);

INVx2_ASAP7_75t_L g3296 ( 
.A(n_3269),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3276),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3283),
.Y(n_3298)
);

AND2x4_ASAP7_75t_L g3299 ( 
.A(n_3259),
.B(n_3250),
.Y(n_3299)
);

AOI31xp33_ASAP7_75t_L g3300 ( 
.A1(n_3267),
.A2(n_3212),
.A3(n_3206),
.B(n_3222),
.Y(n_3300)
);

INVx3_ASAP7_75t_L g3301 ( 
.A(n_3257),
.Y(n_3301)
);

OAI21xp5_ASAP7_75t_L g3302 ( 
.A1(n_3271),
.A2(n_3275),
.B(n_3266),
.Y(n_3302)
);

OR2x6_ASAP7_75t_L g3303 ( 
.A(n_3273),
.B(n_3205),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_3260),
.Y(n_3304)
);

AO21x2_ASAP7_75t_L g3305 ( 
.A1(n_3249),
.A2(n_3239),
.B(n_3207),
.Y(n_3305)
);

OA22x2_ASAP7_75t_L g3306 ( 
.A1(n_3261),
.A2(n_3209),
.B1(n_3223),
.B2(n_618),
.Y(n_3306)
);

BUFx2_ASAP7_75t_L g3307 ( 
.A(n_3277),
.Y(n_3307)
);

HB1xp67_ASAP7_75t_L g3308 ( 
.A(n_3278),
.Y(n_3308)
);

AND3x2_ASAP7_75t_L g3309 ( 
.A(n_3286),
.B(n_615),
.C(n_616),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3274),
.Y(n_3310)
);

XNOR2x1_ASAP7_75t_L g3311 ( 
.A(n_3252),
.B(n_616),
.Y(n_3311)
);

AND2x4_ASAP7_75t_L g3312 ( 
.A(n_3262),
.B(n_618),
.Y(n_3312)
);

INVx2_ASAP7_75t_L g3313 ( 
.A(n_3281),
.Y(n_3313)
);

AND2x4_ASAP7_75t_L g3314 ( 
.A(n_3285),
.B(n_619),
.Y(n_3314)
);

NAND3xp33_ASAP7_75t_SL g3315 ( 
.A(n_3265),
.B(n_619),
.C(n_620),
.Y(n_3315)
);

XOR2x1_ASAP7_75t_L g3316 ( 
.A(n_3251),
.B(n_621),
.Y(n_3316)
);

OR2x2_ASAP7_75t_L g3317 ( 
.A(n_3268),
.B(n_621),
.Y(n_3317)
);

XNOR2x1_ASAP7_75t_L g3318 ( 
.A(n_3288),
.B(n_622),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3263),
.Y(n_3319)
);

AND3x2_ASAP7_75t_L g3320 ( 
.A(n_3287),
.B(n_622),
.C(n_623),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_3312),
.B(n_3253),
.Y(n_3321)
);

XNOR2xp5_ASAP7_75t_L g3322 ( 
.A(n_3311),
.B(n_3254),
.Y(n_3322)
);

INVx2_ASAP7_75t_L g3323 ( 
.A(n_3320),
.Y(n_3323)
);

OR5x1_ASAP7_75t_L g3324 ( 
.A(n_3315),
.B(n_3272),
.C(n_3284),
.D(n_3282),
.E(n_3270),
.Y(n_3324)
);

AOI21x1_ASAP7_75t_L g3325 ( 
.A1(n_3294),
.A2(n_3279),
.B(n_623),
.Y(n_3325)
);

AOI22xp33_ASAP7_75t_L g3326 ( 
.A1(n_3307),
.A2(n_626),
.B1(n_624),
.B2(n_625),
.Y(n_3326)
);

XNOR2xp5_ASAP7_75t_L g3327 ( 
.A(n_3318),
.B(n_3290),
.Y(n_3327)
);

AOI22xp5_ASAP7_75t_L g3328 ( 
.A1(n_3297),
.A2(n_627),
.B1(n_624),
.B2(n_626),
.Y(n_3328)
);

AOI22xp5_ASAP7_75t_L g3329 ( 
.A1(n_3301),
.A2(n_629),
.B1(n_627),
.B2(n_628),
.Y(n_3329)
);

INVxp67_ASAP7_75t_SL g3330 ( 
.A(n_3295),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3289),
.Y(n_3331)
);

NOR2xp33_ASAP7_75t_R g3332 ( 
.A(n_3319),
.B(n_628),
.Y(n_3332)
);

AOI22xp5_ASAP7_75t_L g3333 ( 
.A1(n_3299),
.A2(n_631),
.B1(n_629),
.B2(n_630),
.Y(n_3333)
);

AO21x2_ASAP7_75t_L g3334 ( 
.A1(n_3302),
.A2(n_3298),
.B(n_3310),
.Y(n_3334)
);

NAND4xp25_ASAP7_75t_L g3335 ( 
.A(n_3293),
.B(n_632),
.C(n_630),
.D(n_631),
.Y(n_3335)
);

NOR3xp33_ASAP7_75t_L g3336 ( 
.A(n_3292),
.B(n_3300),
.C(n_3296),
.Y(n_3336)
);

AOI22xp5_ASAP7_75t_L g3337 ( 
.A1(n_3303),
.A2(n_635),
.B1(n_633),
.B2(n_634),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_3337),
.B(n_3309),
.Y(n_3338)
);

OAI22xp5_ASAP7_75t_L g3339 ( 
.A1(n_3331),
.A2(n_3303),
.B1(n_3291),
.B2(n_3317),
.Y(n_3339)
);

OAI22xp5_ASAP7_75t_L g3340 ( 
.A1(n_3330),
.A2(n_3308),
.B1(n_3314),
.B2(n_3304),
.Y(n_3340)
);

AOI21xp5_ASAP7_75t_L g3341 ( 
.A1(n_3321),
.A2(n_3306),
.B(n_3305),
.Y(n_3341)
);

OAI21xp5_ASAP7_75t_SL g3342 ( 
.A1(n_3322),
.A2(n_3313),
.B(n_3316),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_L g3343 ( 
.A(n_3323),
.B(n_634),
.Y(n_3343)
);

AOI22xp5_ASAP7_75t_L g3344 ( 
.A1(n_3336),
.A2(n_637),
.B1(n_635),
.B2(n_636),
.Y(n_3344)
);

INVxp67_ASAP7_75t_SL g3345 ( 
.A(n_3328),
.Y(n_3345)
);

XNOR2xp5_ASAP7_75t_L g3346 ( 
.A(n_3327),
.B(n_636),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3325),
.Y(n_3347)
);

AOI21xp5_ASAP7_75t_L g3348 ( 
.A1(n_3334),
.A2(n_637),
.B(n_638),
.Y(n_3348)
);

AND3x4_ASAP7_75t_L g3349 ( 
.A(n_3324),
.B(n_638),
.C(n_639),
.Y(n_3349)
);

OAI22xp5_ASAP7_75t_L g3350 ( 
.A1(n_3326),
.A2(n_641),
.B1(n_639),
.B2(n_640),
.Y(n_3350)
);

XNOR2xp5_ASAP7_75t_L g3351 ( 
.A(n_3349),
.B(n_3335),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3343),
.Y(n_3352)
);

OAI22x1_ASAP7_75t_SL g3353 ( 
.A1(n_3347),
.A2(n_3332),
.B1(n_3329),
.B2(n_3333),
.Y(n_3353)
);

OAI22xp5_ASAP7_75t_L g3354 ( 
.A1(n_3344),
.A2(n_642),
.B1(n_640),
.B2(n_641),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_3346),
.Y(n_3355)
);

OAI22xp5_ASAP7_75t_L g3356 ( 
.A1(n_3338),
.A2(n_644),
.B1(n_642),
.B2(n_643),
.Y(n_3356)
);

OAI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_3348),
.A2(n_644),
.B(n_645),
.Y(n_3357)
);

CKINVDCx20_ASAP7_75t_R g3358 ( 
.A(n_3339),
.Y(n_3358)
);

INVx1_ASAP7_75t_SL g3359 ( 
.A(n_3350),
.Y(n_3359)
);

OAI22xp5_ASAP7_75t_L g3360 ( 
.A1(n_3345),
.A2(n_648),
.B1(n_646),
.B2(n_647),
.Y(n_3360)
);

INVx2_ASAP7_75t_L g3361 ( 
.A(n_3340),
.Y(n_3361)
);

NAND3xp33_ASAP7_75t_L g3362 ( 
.A(n_3361),
.B(n_3342),
.C(n_3341),
.Y(n_3362)
);

AO22x2_ASAP7_75t_L g3363 ( 
.A1(n_3359),
.A2(n_649),
.B1(n_647),
.B2(n_648),
.Y(n_3363)
);

OAI21xp5_ASAP7_75t_L g3364 ( 
.A1(n_3351),
.A2(n_650),
.B(n_651),
.Y(n_3364)
);

BUFx2_ASAP7_75t_L g3365 ( 
.A(n_3357),
.Y(n_3365)
);

AOI22xp5_ASAP7_75t_L g3366 ( 
.A1(n_3358),
.A2(n_654),
.B1(n_652),
.B2(n_653),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3353),
.Y(n_3367)
);

AOI22xp5_ASAP7_75t_L g3368 ( 
.A1(n_3354),
.A2(n_655),
.B1(n_652),
.B2(n_654),
.Y(n_3368)
);

AOI22xp5_ASAP7_75t_L g3369 ( 
.A1(n_3355),
.A2(n_658),
.B1(n_656),
.B2(n_657),
.Y(n_3369)
);

OAI21xp5_ASAP7_75t_L g3370 ( 
.A1(n_3352),
.A2(n_656),
.B(n_657),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3356),
.B(n_658),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3363),
.Y(n_3372)
);

NOR2xp33_ASAP7_75t_L g3373 ( 
.A(n_3367),
.B(n_3360),
.Y(n_3373)
);

OAI22xp5_ASAP7_75t_L g3374 ( 
.A1(n_3362),
.A2(n_661),
.B1(n_659),
.B2(n_660),
.Y(n_3374)
);

OAI22xp5_ASAP7_75t_L g3375 ( 
.A1(n_3368),
.A2(n_3371),
.B1(n_3365),
.B2(n_3366),
.Y(n_3375)
);

AOI21xp5_ASAP7_75t_L g3376 ( 
.A1(n_3364),
.A2(n_660),
.B(n_661),
.Y(n_3376)
);

AOI221xp5_ASAP7_75t_L g3377 ( 
.A1(n_3363),
.A2(n_664),
.B1(n_662),
.B2(n_663),
.C(n_665),
.Y(n_3377)
);

AOI21xp5_ASAP7_75t_L g3378 ( 
.A1(n_3370),
.A2(n_662),
.B(n_663),
.Y(n_3378)
);

AOI22xp33_ASAP7_75t_L g3379 ( 
.A1(n_3373),
.A2(n_3372),
.B1(n_3376),
.B2(n_3378),
.Y(n_3379)
);

AOI22xp5_ASAP7_75t_L g3380 ( 
.A1(n_3374),
.A2(n_3369),
.B1(n_667),
.B2(n_664),
.Y(n_3380)
);

OA22x2_ASAP7_75t_L g3381 ( 
.A1(n_3375),
.A2(n_668),
.B1(n_666),
.B2(n_667),
.Y(n_3381)
);

OAI21xp5_ASAP7_75t_L g3382 ( 
.A1(n_3377),
.A2(n_666),
.B(n_668),
.Y(n_3382)
);

XNOR2xp5_ASAP7_75t_L g3383 ( 
.A(n_3375),
.B(n_669),
.Y(n_3383)
);

AOI22xp5_ASAP7_75t_L g3384 ( 
.A1(n_3380),
.A2(n_671),
.B1(n_669),
.B2(n_670),
.Y(n_3384)
);

NAND2xp33_ASAP7_75t_SL g3385 ( 
.A(n_3383),
.B(n_670),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_L g3386 ( 
.A(n_3384),
.B(n_3382),
.Y(n_3386)
);

OAI21xp5_ASAP7_75t_SL g3387 ( 
.A1(n_3385),
.A2(n_3379),
.B(n_3381),
.Y(n_3387)
);

AOI21xp5_ASAP7_75t_L g3388 ( 
.A1(n_3387),
.A2(n_671),
.B(n_672),
.Y(n_3388)
);

AOI211xp5_ASAP7_75t_L g3389 ( 
.A1(n_3388),
.A2(n_3386),
.B(n_674),
.C(n_673),
.Y(n_3389)
);


endmodule