module real_aes_7239_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g174 ( .A1(n_0), .A2(n_175), .B(n_178), .C(n_182), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_1), .B(n_166), .Y(n_185) );
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_2), .B(n_105), .C(n_106), .Y(n_104) );
INVx1_ASAP7_75t_L g122 ( .A(n_2), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_3), .B(n_176), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_4), .A2(n_135), .B(n_487), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_5), .A2(n_140), .B(n_143), .C(n_514), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_6), .A2(n_135), .B(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_7), .B(n_166), .Y(n_493) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_8), .A2(n_168), .B(n_243), .Y(n_242) );
AND2x6_ASAP7_75t_L g140 ( .A(n_9), .B(n_141), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_10), .A2(n_140), .B(n_143), .C(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g527 ( .A(n_11), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_12), .B(n_41), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_13), .B(n_181), .Y(n_516) );
INVx1_ASAP7_75t_L g161 ( .A(n_14), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_15), .B(n_176), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_16), .A2(n_177), .B(n_547), .C(n_549), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_17), .B(n_166), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_18), .B(n_155), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g142 ( .A1(n_19), .A2(n_143), .B(n_146), .C(n_154), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_20), .A2(n_180), .B(n_236), .C(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_21), .B(n_181), .Y(n_465) );
AOI222xp33_ASAP7_75t_L g444 ( .A1(n_22), .A2(n_23), .B1(n_445), .B2(n_711), .C1(n_716), .C2(n_717), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_22), .Y(n_716) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_24), .B(n_181), .Y(n_501) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_25), .Y(n_461) );
INVx1_ASAP7_75t_L g500 ( .A(n_26), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_27), .A2(n_143), .B(n_154), .C(n_246), .Y(n_245) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_28), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_29), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_30), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g478 ( .A(n_31), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_32), .A2(n_135), .B(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g138 ( .A(n_33), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_34), .A2(n_194), .B(n_195), .C(n_199), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_35), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_36), .A2(n_180), .B(n_490), .C(n_492), .Y(n_489) );
INVxp67_ASAP7_75t_L g479 ( .A(n_37), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_38), .B(n_248), .Y(n_247) );
CKINVDCx14_ASAP7_75t_R g488 ( .A(n_39), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_40), .A2(n_143), .B(n_154), .C(n_499), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_42), .A2(n_182), .B(n_525), .C(n_526), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_43), .B(n_134), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_44), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_45), .B(n_176), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_46), .B(n_135), .Y(n_244) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_47), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_48), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_49), .A2(n_194), .B(n_199), .C(n_221), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_50), .A2(n_100), .B1(n_111), .B2(n_722), .Y(n_99) );
INVx1_ASAP7_75t_L g179 ( .A(n_51), .Y(n_179) );
INVx1_ASAP7_75t_L g222 ( .A(n_52), .Y(n_222) );
INVx1_ASAP7_75t_L g533 ( .A(n_53), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_54), .B(n_135), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_55), .Y(n_163) );
CKINVDCx14_ASAP7_75t_R g523 ( .A(n_56), .Y(n_523) );
INVx1_ASAP7_75t_L g141 ( .A(n_57), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_58), .B(n_135), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_59), .B(n_166), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_60), .A2(n_153), .B(n_209), .C(n_211), .Y(n_208) );
INVx1_ASAP7_75t_L g160 ( .A(n_61), .Y(n_160) );
INVx1_ASAP7_75t_SL g491 ( .A(n_62), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_63), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_64), .B(n_176), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_65), .B(n_166), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_66), .B(n_177), .Y(n_233) );
INVx1_ASAP7_75t_L g464 ( .A(n_67), .Y(n_464) );
CKINVDCx16_ASAP7_75t_R g172 ( .A(n_68), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_69), .B(n_148), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_70), .A2(n_143), .B(n_199), .C(n_262), .Y(n_261) );
CKINVDCx16_ASAP7_75t_R g207 ( .A(n_71), .Y(n_207) );
INVx1_ASAP7_75t_L g108 ( .A(n_72), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_73), .A2(n_135), .B(n_522), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_74), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_75), .A2(n_135), .B(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_76), .A2(n_124), .B1(n_125), .B2(n_439), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_76), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_77), .A2(n_134), .B(n_474), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g497 ( .A(n_78), .Y(n_497) );
INVx1_ASAP7_75t_L g545 ( .A(n_79), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_80), .B(n_151), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_81), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_82), .A2(n_135), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g548 ( .A(n_83), .Y(n_548) );
INVx2_ASAP7_75t_L g158 ( .A(n_84), .Y(n_158) );
INVx1_ASAP7_75t_L g515 ( .A(n_85), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_86), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_87), .B(n_181), .Y(n_234) );
INVx2_ASAP7_75t_L g105 ( .A(n_88), .Y(n_105) );
OR2x2_ASAP7_75t_L g119 ( .A(n_88), .B(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g448 ( .A(n_88), .B(n_121), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_L g462 ( .A1(n_89), .A2(n_143), .B(n_199), .C(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_90), .B(n_135), .Y(n_192) );
INVx1_ASAP7_75t_L g196 ( .A(n_91), .Y(n_196) );
INVxp67_ASAP7_75t_L g212 ( .A(n_92), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_93), .B(n_168), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_94), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g229 ( .A(n_95), .Y(n_229) );
INVx1_ASAP7_75t_L g263 ( .A(n_96), .Y(n_263) );
INVx2_ASAP7_75t_L g536 ( .A(n_97), .Y(n_536) );
AND2x2_ASAP7_75t_L g224 ( .A(n_98), .B(n_157), .Y(n_224) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_102), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
OR2x2_ASAP7_75t_SL g103 ( .A(n_104), .B(n_109), .Y(n_103) );
OR2x2_ASAP7_75t_L g449 ( .A(n_105), .B(n_121), .Y(n_449) );
NOR2x2_ASAP7_75t_L g719 ( .A(n_105), .B(n_120), .Y(n_719) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g121 ( .A(n_110), .B(n_122), .Y(n_121) );
OA21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_117), .B(n_443), .Y(n_111) );
BUFx2_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_SL g721 ( .A(n_115), .Y(n_721) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OAI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_123), .B(n_440), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_119), .Y(n_442) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_125), .A2(n_446), .B1(n_449), .B2(n_450), .Y(n_445) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_SL g711 ( .A1(n_126), .A2(n_712), .B1(n_713), .B2(n_714), .Y(n_711) );
AND2x2_ASAP7_75t_SL g126 ( .A(n_127), .B(n_375), .Y(n_126) );
NOR5xp2_ASAP7_75t_L g127 ( .A(n_128), .B(n_306), .C(n_335), .D(n_355), .E(n_362), .Y(n_127) );
OAI211xp5_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_186), .B(n_250), .C(n_293), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_130), .A2(n_378), .B1(n_380), .B2(n_381), .Y(n_377) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_165), .Y(n_130) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_131), .Y(n_253) );
AND2x4_ASAP7_75t_L g286 ( .A(n_131), .B(n_287), .Y(n_286) );
INVx5_ASAP7_75t_L g304 ( .A(n_131), .Y(n_304) );
AND2x2_ASAP7_75t_L g313 ( .A(n_131), .B(n_305), .Y(n_313) );
AND2x2_ASAP7_75t_L g325 ( .A(n_131), .B(n_190), .Y(n_325) );
AND2x2_ASAP7_75t_L g421 ( .A(n_131), .B(n_289), .Y(n_421) );
OR2x6_ASAP7_75t_L g131 ( .A(n_132), .B(n_162), .Y(n_131) );
AOI21xp5_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_142), .B(n_155), .Y(n_132) );
BUFx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
NAND2x1p5_ASAP7_75t_L g230 ( .A(n_136), .B(n_140), .Y(n_230) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g153 ( .A(n_137), .Y(n_153) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g144 ( .A(n_138), .Y(n_144) );
INVx1_ASAP7_75t_L g237 ( .A(n_138), .Y(n_237) );
INVx1_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_139), .Y(n_149) );
INVx3_ASAP7_75t_L g177 ( .A(n_139), .Y(n_177) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
INVx1_ASAP7_75t_L g248 ( .A(n_139), .Y(n_248) );
BUFx3_ASAP7_75t_L g154 ( .A(n_140), .Y(n_154) );
INVx4_ASAP7_75t_SL g184 ( .A(n_140), .Y(n_184) );
INVx5_ASAP7_75t_L g173 ( .A(n_143), .Y(n_173) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx3_ASAP7_75t_L g183 ( .A(n_144), .Y(n_183) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_144), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_150), .B(n_152), .Y(n_146) );
INVx2_ASAP7_75t_L g151 ( .A(n_148), .Y(n_151) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx4_ASAP7_75t_L g210 ( .A(n_149), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_151), .A2(n_196), .B(n_197), .C(n_198), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_151), .A2(n_198), .B(n_222), .C(n_223), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_151), .A2(n_464), .B(n_465), .C(n_466), .Y(n_463) );
O2A1O1Ixp5_ASAP7_75t_L g514 ( .A1(n_151), .A2(n_466), .B(n_515), .C(n_516), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_152), .A2(n_176), .B(n_500), .C(n_501), .Y(n_499) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_153), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_156), .B(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g164 ( .A(n_157), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_157), .A2(n_192), .B(n_193), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_157), .A2(n_219), .B(n_220), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_157), .A2(n_230), .B(n_497), .C(n_498), .Y(n_496) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_157), .A2(n_521), .B(n_528), .Y(n_520) );
AND2x2_ASAP7_75t_SL g157 ( .A(n_158), .B(n_159), .Y(n_157) );
AND2x2_ASAP7_75t_L g169 ( .A(n_158), .B(n_159), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_164), .A2(n_511), .B(n_517), .Y(n_510) );
INVx2_ASAP7_75t_L g287 ( .A(n_165), .Y(n_287) );
AND2x2_ASAP7_75t_L g305 ( .A(n_165), .B(n_259), .Y(n_305) );
AND2x2_ASAP7_75t_L g324 ( .A(n_165), .B(n_258), .Y(n_324) );
AND2x2_ASAP7_75t_L g364 ( .A(n_165), .B(n_304), .Y(n_364) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_170), .B(n_185), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_167), .B(n_201), .Y(n_200) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_167), .A2(n_228), .B(n_238), .Y(n_227) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_167), .A2(n_260), .B(n_268), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_167), .B(n_269), .Y(n_268) );
AO21x2_ASAP7_75t_L g459 ( .A1(n_167), .A2(n_460), .B(n_467), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_167), .B(n_503), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_167), .B(n_518), .Y(n_517) );
INVx4_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_168), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_168), .A2(n_244), .B(n_245), .Y(n_243) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g240 ( .A(n_169), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_SL g171 ( .A1(n_172), .A2(n_173), .B(n_174), .C(n_184), .Y(n_171) );
INVx2_ASAP7_75t_L g194 ( .A(n_173), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g206 ( .A1(n_173), .A2(n_184), .B(n_207), .C(n_208), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_SL g474 ( .A1(n_173), .A2(n_184), .B(n_475), .C(n_476), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_173), .A2(n_184), .B(n_488), .C(n_489), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_SL g522 ( .A1(n_173), .A2(n_184), .B(n_523), .C(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_SL g532 ( .A1(n_173), .A2(n_184), .B(n_533), .C(n_534), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_SL g544 ( .A1(n_173), .A2(n_184), .B(n_545), .C(n_546), .Y(n_544) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_176), .B(n_212), .Y(n_211) );
OAI22xp33_ASAP7_75t_L g477 ( .A1(n_176), .A2(n_210), .B1(n_478), .B2(n_479), .Y(n_477) );
INVx5_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_177), .B(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_180), .B(n_491), .Y(n_490) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g525 ( .A(n_181), .Y(n_525) );
INVx2_ASAP7_75t_L g466 ( .A(n_182), .Y(n_466) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_183), .Y(n_198) );
INVx1_ASAP7_75t_L g549 ( .A(n_183), .Y(n_549) );
INVx1_ASAP7_75t_L g199 ( .A(n_184), .Y(n_199) );
INVxp67_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_188), .B(n_214), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AOI322xp5_ASAP7_75t_L g423 ( .A1(n_189), .A2(n_225), .A3(n_278), .B1(n_286), .B2(n_340), .C1(n_424), .C2(n_427), .Y(n_423) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_202), .Y(n_189) );
INVx5_ASAP7_75t_L g255 ( .A(n_190), .Y(n_255) );
AND2x2_ASAP7_75t_L g272 ( .A(n_190), .B(n_257), .Y(n_272) );
BUFx2_ASAP7_75t_L g350 ( .A(n_190), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_190), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g427 ( .A(n_190), .B(n_334), .Y(n_427) );
OR2x6_ASAP7_75t_L g190 ( .A(n_191), .B(n_200), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_202), .B(n_216), .Y(n_281) );
INVx1_ASAP7_75t_L g308 ( .A(n_202), .Y(n_308) );
AND2x2_ASAP7_75t_L g321 ( .A(n_202), .B(n_241), .Y(n_321) );
AND2x2_ASAP7_75t_L g422 ( .A(n_202), .B(n_340), .Y(n_422) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
OR2x2_ASAP7_75t_L g276 ( .A(n_203), .B(n_216), .Y(n_276) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_203), .Y(n_284) );
OR2x2_ASAP7_75t_L g291 ( .A(n_203), .B(n_241), .Y(n_291) );
AND2x2_ASAP7_75t_L g301 ( .A(n_203), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_203), .B(n_227), .Y(n_330) );
INVxp67_ASAP7_75t_L g354 ( .A(n_203), .Y(n_354) );
AND2x2_ASAP7_75t_L g361 ( .A(n_203), .B(n_225), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_203), .B(n_241), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_203), .B(n_226), .Y(n_387) );
OA21x2_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_213), .Y(n_203) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_204), .A2(n_486), .B(n_493), .Y(n_485) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_204), .A2(n_531), .B(n_537), .Y(n_530) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_204), .A2(n_543), .B(n_550), .Y(n_542) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_209), .A2(n_263), .B(n_264), .C(n_265), .Y(n_262) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_210), .B(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_210), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_225), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_216), .B(n_242), .Y(n_331) );
OR2x2_ASAP7_75t_L g353 ( .A(n_216), .B(n_226), .Y(n_353) );
AND2x2_ASAP7_75t_L g366 ( .A(n_216), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_216), .B(n_321), .Y(n_372) );
OAI211xp5_ASAP7_75t_SL g376 ( .A1(n_216), .A2(n_377), .B(n_382), .C(n_391), .Y(n_376) );
AND2x2_ASAP7_75t_L g437 ( .A(n_216), .B(n_241), .Y(n_437) );
INVx5_ASAP7_75t_SL g216 ( .A(n_217), .Y(n_216) );
OR2x2_ASAP7_75t_L g290 ( .A(n_217), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_217), .B(n_296), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_217), .B(n_285), .Y(n_297) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_217), .Y(n_299) );
OR2x2_ASAP7_75t_L g310 ( .A(n_217), .B(n_226), .Y(n_310) );
AND2x2_ASAP7_75t_SL g315 ( .A(n_217), .B(n_301), .Y(n_315) );
AND2x2_ASAP7_75t_L g340 ( .A(n_217), .B(n_226), .Y(n_340) );
AND2x2_ASAP7_75t_L g360 ( .A(n_217), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g398 ( .A(n_217), .B(n_225), .Y(n_398) );
OR2x2_ASAP7_75t_L g401 ( .A(n_217), .B(n_387), .Y(n_401) );
OR2x6_ASAP7_75t_L g217 ( .A(n_218), .B(n_224), .Y(n_217) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_241), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g344 ( .A1(n_226), .A2(n_345), .B(n_348), .C(n_354), .Y(n_344) );
INVx5_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_227), .B(n_241), .Y(n_275) );
AND2x2_ASAP7_75t_L g279 ( .A(n_227), .B(n_242), .Y(n_279) );
OR2x2_ASAP7_75t_L g285 ( .A(n_227), .B(n_241), .Y(n_285) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_231), .Y(n_228) );
OAI21xp5_ASAP7_75t_L g460 ( .A1(n_230), .A2(n_461), .B(n_462), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g511 ( .A1(n_230), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_235), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_235), .A2(n_247), .B(n_249), .Y(n_246) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
INVx2_ASAP7_75t_L g471 ( .A(n_240), .Y(n_471) );
INVx1_ASAP7_75t_SL g302 ( .A(n_241), .Y(n_302) );
OR2x2_ASAP7_75t_L g430 ( .A(n_241), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_270), .B(n_273), .C(n_282), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AOI31xp33_ASAP7_75t_L g355 ( .A1(n_252), .A2(n_356), .A3(n_358), .B(n_359), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_253), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_254), .B(n_286), .Y(n_292) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_255), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g312 ( .A(n_255), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g317 ( .A(n_255), .B(n_287), .Y(n_317) );
AND2x2_ASAP7_75t_L g327 ( .A(n_255), .B(n_286), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_255), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g347 ( .A(n_255), .B(n_304), .Y(n_347) );
AND2x2_ASAP7_75t_L g352 ( .A(n_255), .B(n_324), .Y(n_352) );
OR2x2_ASAP7_75t_L g371 ( .A(n_255), .B(n_257), .Y(n_371) );
OR2x2_ASAP7_75t_L g373 ( .A(n_255), .B(n_374), .Y(n_373) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_255), .Y(n_420) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g320 ( .A(n_257), .B(n_287), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_257), .B(n_304), .Y(n_343) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
BUFx2_ASAP7_75t_L g289 ( .A(n_259), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_267), .Y(n_260) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx3_ASAP7_75t_L g492 ( .A(n_266), .Y(n_492) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g380 ( .A(n_272), .B(n_304), .Y(n_380) );
AOI322xp5_ASAP7_75t_L g382 ( .A1(n_272), .A2(n_286), .A3(n_324), .B1(n_383), .B2(n_384), .C1(n_385), .C2(n_388), .Y(n_382) );
INVx1_ASAP7_75t_L g390 ( .A(n_272), .Y(n_390) );
NAND2xp33_ASAP7_75t_L g273 ( .A(n_274), .B(n_277), .Y(n_273) );
INVx1_ASAP7_75t_SL g384 ( .A(n_274), .Y(n_384) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
OR2x2_ASAP7_75t_L g336 ( .A(n_275), .B(n_281), .Y(n_336) );
INVx1_ASAP7_75t_L g367 ( .A(n_275), .Y(n_367) );
INVx2_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OAI32xp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_286), .A3(n_288), .B1(n_290), .B2(n_292), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AOI21xp33_ASAP7_75t_SL g322 ( .A1(n_285), .A2(n_300), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g337 ( .A(n_286), .Y(n_337) );
AND2x4_ASAP7_75t_L g334 ( .A(n_287), .B(n_304), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_287), .B(n_370), .Y(n_369) );
AOI322xp5_ASAP7_75t_L g399 ( .A1(n_288), .A2(n_315), .A3(n_334), .B1(n_367), .B2(n_400), .C1(n_402), .C2(n_403), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g428 ( .A1(n_288), .A2(n_365), .B1(n_429), .B2(n_430), .C(n_432), .Y(n_428) );
AND2x2_ASAP7_75t_L g316 ( .A(n_289), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_SL g296 ( .A(n_291), .Y(n_296) );
OR2x2_ASAP7_75t_L g368 ( .A(n_291), .B(n_353), .Y(n_368) );
OAI31xp33_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_297), .A3(n_298), .B(n_303), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_294), .A2(n_327), .B1(n_328), .B2(n_332), .Y(n_326) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g339 ( .A(n_296), .B(n_340), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_298), .A2(n_339), .B1(n_392), .B2(n_395), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g381 ( .A(n_301), .B(n_350), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_301), .B(n_340), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_302), .B(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g415 ( .A(n_302), .B(n_353), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_303), .A2(n_398), .B1(n_411), .B2(n_414), .Y(n_410) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx2_ASAP7_75t_L g319 ( .A(n_304), .Y(n_319) );
AND2x2_ASAP7_75t_L g402 ( .A(n_304), .B(n_324), .Y(n_402) );
OR2x2_ASAP7_75t_L g404 ( .A(n_304), .B(n_371), .Y(n_404) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_304), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_305), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_305), .B(n_350), .Y(n_358) );
OAI211xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_311), .B(n_314), .C(n_326), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AOI221xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_316), .B1(n_318), .B2(n_321), .C(n_322), .Y(n_314) );
INVxp67_ASAP7_75t_L g426 ( .A(n_317), .Y(n_426) );
INVx1_ASAP7_75t_L g393 ( .A(n_318), .Y(n_393) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g357 ( .A(n_319), .B(n_324), .Y(n_357) );
INVx1_ASAP7_75t_L g374 ( .A(n_320), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_320), .B(n_347), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g389 ( .A(n_324), .Y(n_389) );
AND2x2_ASAP7_75t_L g395 ( .A(n_324), .B(n_350), .Y(n_395) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_SL g383 ( .A(n_331), .Y(n_383) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_334), .B(n_370), .Y(n_394) );
OAI221xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_337), .B1(n_338), .B2(n_341), .C(n_344), .Y(n_335) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g431 ( .A(n_340), .Y(n_431) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g349 ( .A(n_343), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_347), .B(n_406), .Y(n_405) );
AOI21xp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_351), .B(n_353), .Y(n_348) );
OAI211xp5_ASAP7_75t_SL g396 ( .A1(n_351), .A2(n_397), .B(n_399), .C(n_405), .Y(n_396) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g408 ( .A(n_353), .Y(n_408) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OAI222xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_365), .B1(n_368), .B2(n_369), .C1(n_372), .C2(n_373), .Y(n_362) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g438 ( .A(n_369), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_370), .B(n_413), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_370), .A2(n_417), .B1(n_419), .B2(n_422), .Y(n_416) );
INVx2_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
NOR4xp25_ASAP7_75t_L g375 ( .A(n_376), .B(n_396), .C(n_409), .D(n_428), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_378), .B(n_408), .Y(n_418) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g385 ( .A(n_383), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_386), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND3xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_416), .C(n_423), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx2_ASAP7_75t_L g425 ( .A(n_421), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
OAI21xp5_ASAP7_75t_SL g432 ( .A1(n_433), .A2(n_435), .B(n_438), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND3xp33_ASAP7_75t_L g443 ( .A(n_440), .B(n_444), .C(n_720), .Y(n_443) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g712 ( .A(n_447), .Y(n_712) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g715 ( .A(n_449), .Y(n_715) );
INVx2_ASAP7_75t_L g713 ( .A(n_450), .Y(n_713) );
OR2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_645), .Y(n_450) );
NAND5xp2_ASAP7_75t_L g451 ( .A(n_452), .B(n_574), .C(n_604), .D(n_625), .E(n_631), .Y(n_451) );
AOI221xp5_ASAP7_75t_SL g452 ( .A1(n_453), .A2(n_507), .B1(n_538), .B2(n_540), .C(n_551), .Y(n_452) );
INVxp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_455), .B(n_504), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_482), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_SL g625 ( .A1(n_457), .A2(n_494), .B(n_626), .C(n_629), .Y(n_625) );
AND2x2_ASAP7_75t_L g695 ( .A(n_457), .B(n_495), .Y(n_695) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_469), .Y(n_457) );
AND2x2_ASAP7_75t_L g553 ( .A(n_458), .B(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g557 ( .A(n_458), .B(n_554), .Y(n_557) );
OR2x2_ASAP7_75t_L g583 ( .A(n_458), .B(n_495), .Y(n_583) );
AND2x2_ASAP7_75t_L g585 ( .A(n_458), .B(n_485), .Y(n_585) );
AND2x2_ASAP7_75t_L g603 ( .A(n_458), .B(n_484), .Y(n_603) );
INVx1_ASAP7_75t_L g636 ( .A(n_458), .Y(n_636) );
INVx2_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
BUFx2_ASAP7_75t_L g506 ( .A(n_459), .Y(n_506) );
AND2x2_ASAP7_75t_L g539 ( .A(n_459), .B(n_485), .Y(n_539) );
AND2x2_ASAP7_75t_L g692 ( .A(n_459), .B(n_495), .Y(n_692) );
AND2x2_ASAP7_75t_L g573 ( .A(n_469), .B(n_483), .Y(n_573) );
OR2x2_ASAP7_75t_L g577 ( .A(n_469), .B(n_495), .Y(n_577) );
AND2x2_ASAP7_75t_L g602 ( .A(n_469), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_SL g649 ( .A(n_469), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_469), .B(n_611), .Y(n_697) );
AO21x2_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_472), .B(n_480), .Y(n_469) );
INVx1_ASAP7_75t_L g555 ( .A(n_470), .Y(n_555) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OA21x2_ASAP7_75t_L g554 ( .A1(n_473), .A2(n_481), .B(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OAI322xp33_ASAP7_75t_L g698 ( .A1(n_482), .A2(n_634), .A3(n_657), .B1(n_678), .B2(n_699), .C1(n_701), .C2(n_702), .Y(n_698) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_483), .B(n_554), .Y(n_701) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_494), .Y(n_483) );
AND2x2_ASAP7_75t_L g505 ( .A(n_484), .B(n_506), .Y(n_505) );
AND2x4_ASAP7_75t_L g570 ( .A(n_484), .B(n_495), .Y(n_570) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g611 ( .A(n_485), .B(n_495), .Y(n_611) );
AND2x2_ASAP7_75t_L g655 ( .A(n_485), .B(n_494), .Y(n_655) );
AND2x2_ASAP7_75t_L g538 ( .A(n_494), .B(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g556 ( .A(n_494), .B(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_494), .B(n_585), .Y(n_709) );
INVx3_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g504 ( .A(n_495), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_495), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g623 ( .A(n_495), .B(n_554), .Y(n_623) );
AND2x2_ASAP7_75t_L g650 ( .A(n_495), .B(n_585), .Y(n_650) );
OR2x2_ASAP7_75t_L g706 ( .A(n_495), .B(n_557), .Y(n_706) );
OR2x6_ASAP7_75t_L g495 ( .A(n_496), .B(n_502), .Y(n_495) );
INVx1_ASAP7_75t_SL g592 ( .A(n_504), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_505), .B(n_623), .Y(n_624) );
AND2x2_ASAP7_75t_L g658 ( .A(n_505), .B(n_648), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_505), .B(n_581), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_505), .B(n_703), .Y(n_702) );
OAI31xp33_ASAP7_75t_L g676 ( .A1(n_507), .A2(n_538), .A3(n_677), .B(n_679), .Y(n_676) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_519), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_508), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g659 ( .A(n_508), .B(n_594), .Y(n_659) );
OR2x2_ASAP7_75t_L g666 ( .A(n_508), .B(n_667), .Y(n_666) );
OR2x2_ASAP7_75t_L g678 ( .A(n_508), .B(n_567), .Y(n_678) );
CKINVDCx16_ASAP7_75t_R g508 ( .A(n_509), .Y(n_508) );
OR2x2_ASAP7_75t_L g612 ( .A(n_509), .B(n_613), .Y(n_612) );
BUFx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g540 ( .A(n_510), .B(n_541), .Y(n_540) );
INVx4_ASAP7_75t_L g561 ( .A(n_510), .Y(n_561) );
AND2x2_ASAP7_75t_L g598 ( .A(n_510), .B(n_542), .Y(n_598) );
AND2x2_ASAP7_75t_L g597 ( .A(n_519), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_SL g667 ( .A(n_519), .Y(n_667) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_529), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_520), .B(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g567 ( .A(n_520), .B(n_530), .Y(n_567) );
INVx2_ASAP7_75t_L g587 ( .A(n_520), .Y(n_587) );
AND2x2_ASAP7_75t_L g601 ( .A(n_520), .B(n_530), .Y(n_601) );
AND2x2_ASAP7_75t_L g608 ( .A(n_520), .B(n_564), .Y(n_608) );
BUFx3_ASAP7_75t_L g618 ( .A(n_520), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_520), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g563 ( .A(n_529), .Y(n_563) );
AND2x2_ASAP7_75t_L g571 ( .A(n_529), .B(n_561), .Y(n_571) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g541 ( .A(n_530), .B(n_542), .Y(n_541) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_530), .Y(n_595) );
INVx2_ASAP7_75t_SL g578 ( .A(n_539), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_539), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_539), .B(n_648), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_540), .B(n_618), .Y(n_671) );
INVx1_ASAP7_75t_SL g705 ( .A(n_540), .Y(n_705) );
INVx1_ASAP7_75t_SL g613 ( .A(n_541), .Y(n_613) );
INVx1_ASAP7_75t_SL g564 ( .A(n_542), .Y(n_564) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_542), .Y(n_575) );
OR2x2_ASAP7_75t_L g586 ( .A(n_542), .B(n_561), .Y(n_586) );
AND2x2_ASAP7_75t_L g600 ( .A(n_542), .B(n_561), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_542), .B(n_590), .Y(n_652) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_556), .B(n_558), .C(n_569), .Y(n_551) );
AOI31xp33_ASAP7_75t_L g668 ( .A1(n_552), .A2(n_669), .A3(n_670), .B(n_671), .Y(n_668) );
AND2x2_ASAP7_75t_L g641 ( .A(n_553), .B(n_570), .Y(n_641) );
BUFx3_ASAP7_75t_L g581 ( .A(n_554), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_554), .B(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g617 ( .A(n_554), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_554), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_SL g572 ( .A(n_557), .Y(n_572) );
OAI222xp33_ASAP7_75t_L g681 ( .A1(n_557), .A2(n_682), .B1(n_685), .B2(n_686), .C1(n_687), .C2(n_688), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_565), .Y(n_558) );
INVx1_ASAP7_75t_L g687 ( .A(n_559), .Y(n_687) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_561), .B(n_564), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_561), .B(n_587), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_561), .B(n_562), .Y(n_657) );
INVx1_ASAP7_75t_L g708 ( .A(n_561), .Y(n_708) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_562), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g710 ( .A(n_562), .Y(n_710) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx2_ASAP7_75t_L g590 ( .A(n_563), .Y(n_590) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_564), .Y(n_633) );
AOI32xp33_ASAP7_75t_L g569 ( .A1(n_565), .A2(n_570), .A3(n_571), .B1(n_572), .B2(n_573), .Y(n_569) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_567), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g644 ( .A(n_567), .Y(n_644) );
OR2x2_ASAP7_75t_L g685 ( .A(n_567), .B(n_586), .Y(n_685) );
INVx1_ASAP7_75t_L g621 ( .A(n_568), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_570), .B(n_581), .Y(n_606) );
INVx3_ASAP7_75t_L g615 ( .A(n_570), .Y(n_615) );
AOI322xp5_ASAP7_75t_L g631 ( .A1(n_570), .A2(n_615), .A3(n_632), .B1(n_634), .B2(n_637), .C1(n_641), .C2(n_642), .Y(n_631) );
AND2x2_ASAP7_75t_L g607 ( .A(n_571), .B(n_608), .Y(n_607) );
INVxp67_ASAP7_75t_L g684 ( .A(n_571), .Y(n_684) );
A2O1A1O1Ixp25_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B(n_579), .C(n_587), .D(n_588), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_575), .B(n_618), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
OAI221xp5_ASAP7_75t_L g588 ( .A1(n_577), .A2(n_589), .B1(n_592), .B2(n_593), .C(n_596), .Y(n_588) );
INVx1_ASAP7_75t_SL g703 ( .A(n_577), .Y(n_703) );
AOI21xp33_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_584), .B(n_586), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_581), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OAI221xp5_ASAP7_75t_SL g673 ( .A1(n_583), .A2(n_667), .B1(n_674), .B2(n_675), .C(n_676), .Y(n_673) );
OAI222xp33_ASAP7_75t_L g704 ( .A1(n_584), .A2(n_705), .B1(n_706), .B2(n_707), .C1(n_709), .C2(n_710), .Y(n_704) );
AND2x2_ASAP7_75t_L g662 ( .A(n_585), .B(n_648), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_585), .A2(n_600), .B(n_647), .Y(n_674) );
INVx1_ASAP7_75t_L g688 ( .A(n_585), .Y(n_688) );
INVx2_ASAP7_75t_SL g591 ( .A(n_586), .Y(n_591) );
AND2x2_ASAP7_75t_L g594 ( .A(n_587), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx1_ASAP7_75t_SL g628 ( .A(n_590), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_590), .B(n_600), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_591), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_591), .B(n_601), .Y(n_630) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OAI21xp5_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_599), .B(n_602), .Y(n_596) );
INVx1_ASAP7_75t_SL g614 ( .A(n_598), .Y(n_614) );
AND2x2_ASAP7_75t_L g661 ( .A(n_598), .B(n_644), .Y(n_661) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
AND2x2_ASAP7_75t_L g700 ( .A(n_600), .B(n_618), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_601), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g686 ( .A(n_602), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_607), .B1(n_609), .B2(n_616), .C(n_619), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_612), .B1(n_614), .B2(n_615), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_613), .A2(n_620), .B1(n_622), .B2(n_624), .Y(n_619) );
OR2x2_ASAP7_75t_L g690 ( .A(n_614), .B(n_618), .Y(n_690) );
OR2x2_ASAP7_75t_L g693 ( .A(n_614), .B(n_628), .Y(n_693) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI221xp5_ASAP7_75t_L g689 ( .A1(n_635), .A2(n_690), .B1(n_691), .B2(n_693), .C(n_694), .Y(n_689) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVxp67_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND3xp33_ASAP7_75t_SL g645 ( .A(n_646), .B(n_660), .C(n_672), .Y(n_645) );
AOI222xp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_651), .B1(n_653), .B2(n_656), .C1(n_658), .C2(n_659), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_648), .B(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g670 ( .A(n_650), .Y(n_670) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .B1(n_663), .B2(n_665), .C(n_668), .Y(n_660) );
INVx1_ASAP7_75t_L g675 ( .A(n_661), .Y(n_675) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OAI21xp33_ASAP7_75t_L g694 ( .A1(n_665), .A2(n_695), .B(n_696), .Y(n_694) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
NOR5xp2_ASAP7_75t_L g672 ( .A(n_673), .B(n_681), .C(n_689), .D(n_698), .E(n_704), .Y(n_672) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVxp67_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx3_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
endmodule