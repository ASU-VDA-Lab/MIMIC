module fake_jpeg_11066_n_134 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_30),
.Y(n_61)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_12),
.B(n_0),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_45),
.Y(n_52)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_40),
.Y(n_66)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_42),
.Y(n_71)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_1),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_1),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_13),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_23),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_31),
.A2(n_15),
.B1(n_23),
.B2(n_16),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_58),
.B1(n_67),
.B2(n_32),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_15),
.B1(n_11),
.B2(n_14),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_11),
.B1(n_26),
.B2(n_13),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_60),
.A2(n_68),
.B1(n_67),
.B2(n_50),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_62),
.B(n_65),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_28),
.B(n_26),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_69),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_30),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_37),
.A2(n_24),
.B1(n_22),
.B2(n_21),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_38),
.A2(n_24),
.B1(n_22),
.B2(n_21),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_17),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_52),
.Y(n_85)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_65),
.B(n_10),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_76),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_82),
.B1(n_55),
.B2(n_56),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_2),
.Y(n_76)
);

AOI32xp33_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_2),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_77),
.B(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_81),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_61),
.A2(n_4),
.B1(n_6),
.B2(n_71),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_56),
.B1(n_53),
.B2(n_64),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_64),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_59),
.C(n_78),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_50),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_48),
.B(n_51),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_89),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_95),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_96),
.B(n_100),
.Y(n_109)
);

CKINVDCx12_ASAP7_75t_R g95 ( 
.A(n_83),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_97),
.A2(n_73),
.B1(n_86),
.B2(n_75),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_72),
.A2(n_51),
.B(n_59),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_59),
.B(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_85),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_81),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_107),
.Y(n_116)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_110),
.B1(n_96),
.B2(n_98),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_82),
.B1(n_85),
.B2(n_78),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_73),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_111),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_97),
.A2(n_101),
.B1(n_92),
.B2(n_102),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_99),
.B(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_93),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_113),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_117),
.B(n_120),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_118),
.A2(n_116),
.B1(n_104),
.B2(n_107),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_103),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_110),
.B(n_106),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_111),
.C(n_103),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_122),
.A2(n_124),
.B(n_109),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_123),
.A2(n_109),
.B1(n_95),
.B2(n_116),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_128),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_125),
.C(n_114),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_114),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_130),
.B(n_125),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_90),
.A3(n_98),
.B1(n_128),
.B2(n_131),
.C1(n_125),
.C2(n_132),
.Y(n_134)
);


endmodule