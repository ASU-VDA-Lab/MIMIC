module fake_jpeg_6608_n_125 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_125);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx2_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx2_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_27),
.A2(n_10),
.B1(n_11),
.B2(n_30),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_13),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_9),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_39),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

OR2x2_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_1),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_18),
.B1(n_23),
.B2(n_10),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_30),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_13),
.B(n_4),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_25),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_6),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_24),
.B1(n_22),
.B2(n_14),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_27),
.B1(n_38),
.B2(n_30),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_16),
.B1(n_5),
.B2(n_4),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_45),
.B1(n_51),
.B2(n_57),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_16),
.B1(n_5),
.B2(n_4),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_25),
.B1(n_17),
.B2(n_21),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_40),
.B1(n_27),
.B2(n_38),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_21),
.C(n_18),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_52),
.Y(n_64)
);

OAI22x1_ASAP7_75t_L g51 ( 
.A1(n_31),
.A2(n_16),
.B1(n_23),
.B2(n_5),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_45),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_55),
.B(n_56),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_61),
.Y(n_68)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_77),
.B1(n_47),
.B2(n_48),
.Y(n_87)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_59),
.B1(n_71),
.B2(n_62),
.Y(n_91)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_76),
.Y(n_85)
);

NAND3xp33_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_78),
.C(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_51),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_43),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_90),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_49),
.C(n_43),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_73),
.C(n_64),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_56),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_87),
.B(n_74),
.Y(n_97)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_41),
.Y(n_88)
);

AOI21x1_ASAP7_75t_SL g90 ( 
.A1(n_70),
.A2(n_41),
.B(n_54),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_91),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_97),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_86),
.B(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_96),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_66),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_80),
.C(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_99),
.B(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_63),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_106),
.C(n_101),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_88),
.C(n_85),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_92),
.B1(n_90),
.B2(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_96),
.A2(n_92),
.B(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_100),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_111),
.C(n_113),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_105),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_94),
.B1(n_89),
.B2(n_83),
.Y(n_114)
);

OAI21x1_ASAP7_75t_SL g117 ( 
.A1(n_114),
.A2(n_102),
.B(n_105),
.Y(n_117)
);

AOI21x1_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_102),
.B(n_101),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_SL g120 ( 
.A1(n_116),
.A2(n_117),
.B(n_118),
.C(n_69),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_115),
.A2(n_110),
.B(n_104),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_119),
.B(n_82),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_120),
.A2(n_72),
.B(n_76),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_122),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_67),
.Y(n_125)
);


endmodule