module fake_jpeg_22689_n_317 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

HAxp5_ASAP7_75t_SL g58 ( 
.A(n_31),
.B(n_33),
.CON(n_58),
.SN(n_58)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_36),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_42),
.Y(n_60)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_43),
.Y(n_71)
);

OR2x2_ASAP7_75t_SL g44 ( 
.A(n_29),
.B(n_33),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_31),
.A2(n_28),
.B1(n_14),
.B2(n_16),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_28),
.B1(n_14),
.B2(n_26),
.Y(n_61)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_16),
.Y(n_68)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_52),
.B1(n_42),
.B2(n_34),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_28),
.B1(n_14),
.B2(n_16),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_76),
.B1(n_27),
.B2(n_21),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_58),
.A2(n_28),
.B1(n_16),
.B2(n_26),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_66),
.B(n_47),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_26),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_70),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_37),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_75),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_40),
.A2(n_26),
.B1(n_38),
.B2(n_20),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_48),
.B1(n_40),
.B2(n_57),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_36),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_18),
.B1(n_24),
.B2(n_25),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_37),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_56),
.Y(n_87)
);

AND2x4_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_96),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_102),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_93),
.B1(n_76),
.B2(n_70),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_41),
.C(n_45),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_98),
.C(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_18),
.Y(n_90)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_97),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_59),
.A2(n_24),
.B1(n_18),
.B2(n_15),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_23),
.B1(n_25),
.B2(n_24),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_21),
.Y(n_94)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_59),
.A2(n_19),
.B1(n_21),
.B2(n_15),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_66),
.A2(n_20),
.B1(n_23),
.B2(n_25),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_66),
.B(n_34),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_99),
.A2(n_77),
.B1(n_79),
.B2(n_72),
.Y(n_115)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_20),
.B1(n_25),
.B2(n_23),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_103),
.B1(n_34),
.B2(n_30),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_64),
.B(n_27),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_75),
.B1(n_61),
.B2(n_62),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_75),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_67),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_105),
.A2(n_106),
.B1(n_101),
.B2(n_97),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_59),
.B1(n_67),
.B2(n_75),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_107),
.A2(n_81),
.B1(n_79),
.B2(n_77),
.Y(n_151)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_109),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_92),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_113),
.A2(n_117),
.B(n_123),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_115),
.Y(n_145)
);

XNOR2x1_ASAP7_75t_SL g132 ( 
.A(n_116),
.B(n_127),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_13),
.Y(n_117)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_120),
.Y(n_140)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_85),
.A2(n_72),
.B1(n_79),
.B2(n_60),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_84),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_122),
.Y(n_137)
);

AND2x6_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_13),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_128),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_126),
.A2(n_85),
.B1(n_84),
.B2(n_83),
.Y(n_130)
);

NOR2x1p5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_30),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_71),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_106),
.B1(n_119),
.B2(n_126),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_98),
.B(n_83),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_32),
.B(n_30),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_89),
.Y(n_135)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_136),
.B(n_139),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_122),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_138),
.Y(n_156)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_102),
.B(n_98),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_141),
.A2(n_150),
.B(n_117),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_114),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_143),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_103),
.B1(n_91),
.B2(n_99),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_116),
.A2(n_99),
.B1(n_89),
.B2(n_96),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_105),
.A2(n_104),
.B1(n_93),
.B2(n_95),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_112),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_111),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_113),
.B(n_127),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_151),
.Y(n_171)
);

OA21x2_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_109),
.B(n_121),
.Y(n_152)
);

AO22x1_ASAP7_75t_L g155 ( 
.A1(n_152),
.A2(n_132),
.B1(n_119),
.B2(n_129),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_94),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_90),
.Y(n_154)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_152),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_125),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_135),
.C(n_134),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_177),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_140),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_172),
.Y(n_190)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_170),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_110),
.C(n_123),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_173),
.A2(n_174),
.B1(n_178),
.B2(n_132),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_150),
.A2(n_110),
.B(n_71),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_148),
.A2(n_120),
.B1(n_118),
.B2(n_114),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_175),
.A2(n_176),
.B1(n_147),
.B2(n_145),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_148),
.A2(n_77),
.B1(n_63),
.B2(n_65),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_114),
.B1(n_63),
.B2(n_65),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_136),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_143),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_180),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_17),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_181),
.B(n_150),
.Y(n_205)
);

NOR4xp25_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_131),
.C(n_138),
.D(n_132),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_183),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_186),
.A2(n_160),
.B1(n_144),
.B2(n_152),
.Y(n_222)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_188),
.A2(n_195),
.B1(n_196),
.B2(n_180),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_156),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_189),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_168),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_192),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_199),
.Y(n_213)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_197),
.A2(n_164),
.B1(n_179),
.B2(n_170),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_159),
.C(n_158),
.Y(n_211)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_204),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_145),
.B1(n_148),
.B2(n_130),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_155),
.Y(n_207)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_206),
.A2(n_191),
.B(n_187),
.Y(n_210)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_196),
.B(n_146),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_217),
.Y(n_236)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_214),
.C(n_218),
.Y(n_234)
);

NOR2x1_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_166),
.Y(n_212)
);

O2A1O1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_212),
.A2(n_27),
.B(n_19),
.C(n_25),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_158),
.C(n_134),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_215),
.A2(n_216),
.B1(n_165),
.B2(n_152),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_188),
.A2(n_164),
.B1(n_173),
.B2(n_171),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_146),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_177),
.C(n_174),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_222),
.A2(n_223),
.B1(n_227),
.B2(n_219),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_185),
.B1(n_199),
.B2(n_194),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_161),
.C(n_141),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_225),
.C(n_165),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_161),
.C(n_141),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_130),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_149),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_222),
.A2(n_197),
.B1(n_201),
.B2(n_190),
.Y(n_229)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_153),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_233),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_231),
.A2(n_240),
.B1(n_218),
.B2(n_219),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_152),
.Y(n_233)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_243),
.C(n_246),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_220),
.A2(n_182),
.B1(n_185),
.B2(n_168),
.Y(n_238)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_239),
.B(n_245),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_216),
.A2(n_191),
.B1(n_195),
.B2(n_193),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_151),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_223),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_17),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_242),
.B(n_248),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_56),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_19),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_212),
.B(n_20),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_78),
.C(n_23),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_226),
.B(n_13),
.Y(n_248)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_250),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_213),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_261),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_254),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_257),
.A2(n_233),
.B1(n_78),
.B2(n_2),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_245),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_258),
.A2(n_263),
.B(n_230),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_213),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_225),
.C(n_224),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_265),
.C(n_237),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_210),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_246),
.B(n_208),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_256),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_78),
.C(n_23),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_270),
.C(n_280),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_243),
.C(n_236),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_276),
.C(n_254),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_269),
.A2(n_277),
.B(n_261),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_236),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_271),
.B(n_273),
.Y(n_288)
);

INVxp33_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

INVx11_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_260),
.B(n_239),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_275),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_263),
.B(n_0),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_32),
.C(n_1),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_265),
.A2(n_0),
.B(n_1),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_270),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_17),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_257),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_289),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_282),
.A2(n_2),
.B(n_3),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_283),
.A2(n_286),
.B1(n_3),
.B2(n_4),
.Y(n_297)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_279),
.Y(n_284)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_284),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_276),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_1),
.C(n_2),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_268),
.A2(n_1),
.B(n_2),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_290),
.A2(n_272),
.B(n_3),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_280),
.Y(n_295)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_294),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_297),
.Y(n_304)
);

MAJx2_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_298),
.C(n_5),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_17),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_281),
.A2(n_4),
.B(n_5),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_299),
.B(n_6),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_17),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_287),
.A3(n_291),
.B1(n_285),
.B2(n_32),
.C1(n_9),
.C2(n_10),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_303),
.Y(n_308)
);

AOI322xp5_ASAP7_75t_L g305 ( 
.A1(n_293),
.A2(n_291),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_5),
.C2(n_11),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_306),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_299),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_310),
.C(n_11),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_L g311 ( 
.A1(n_308),
.A2(n_307),
.A3(n_300),
.B1(n_8),
.B2(n_10),
.C1(n_6),
.C2(n_12),
.Y(n_311)
);

NAND3xp33_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_312),
.C(n_7),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_309),
.B(n_11),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_314),
.B(n_7),
.Y(n_315)
);

NAND4xp25_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_7),
.C(n_11),
.D(n_12),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_12),
.C(n_17),
.Y(n_317)
);


endmodule