module fake_jpeg_2599_n_195 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_195);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_1),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_25),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

BUFx4f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

BUFx24_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_61),
.Y(n_92)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_48),
.C(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_58),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_69),
.B1(n_48),
.B2(n_55),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_69),
.B1(n_55),
.B2(n_87),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_58),
.B1(n_50),
.B2(n_59),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_87),
.B1(n_58),
.B2(n_91),
.Y(n_99)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_91),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_54),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_97),
.B(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_66),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_107),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_108),
.B1(n_68),
.B2(n_65),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_64),
.B(n_56),
.C(n_62),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_102),
.B(n_81),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_61),
.B(n_49),
.C(n_68),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_0),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_24),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_21),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_83),
.A2(n_88),
.B1(n_78),
.B2(n_68),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_23),
.Y(n_109)
);

MAJx2_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_88),
.C(n_49),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_4),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_116),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_0),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_126),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_65),
.B(n_2),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_1),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_127),
.B(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_109),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_129),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_3),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_145),
.Y(n_157)
);

AO22x1_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_95),
.B1(n_18),
.B2(n_26),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_148),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_3),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_137),
.B(n_139),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_4),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_144),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_45),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_147),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_44),
.B1(n_42),
.B2(n_39),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_146),
.Y(n_169)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_117),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_38),
.Y(n_147)
);

AOI21x1_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_34),
.B(n_33),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_5),
.Y(n_149)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_6),
.Y(n_150)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_163),
.Y(n_175)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_111),
.A3(n_124),
.B1(n_123),
.B2(n_118),
.C1(n_31),
.C2(n_30),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_158),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_118),
.A3(n_29),
.B1(n_28),
.B2(n_27),
.C1(n_10),
.C2(n_11),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_138),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_166),
.B1(n_13),
.B2(n_14),
.Y(n_178)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_151),
.A2(n_146),
.B1(n_142),
.B2(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_143),
.Y(n_173)
);

OAI32xp33_ASAP7_75t_L g168 ( 
.A1(n_143),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_168),
.A2(n_9),
.B(n_12),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_166),
.A2(n_148),
.B(n_133),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_174),
.Y(n_183)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_154),
.C(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_178),
.Y(n_184)
);

OAI321xp33_ASAP7_75t_L g179 ( 
.A1(n_174),
.A2(n_177),
.A3(n_175),
.B1(n_169),
.B2(n_152),
.C(n_171),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_153),
.Y(n_185)
);

AOI322xp5_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_152),
.A3(n_162),
.B1(n_160),
.B2(n_168),
.C1(n_164),
.C2(n_156),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_181),
.A2(n_159),
.B(n_153),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_186),
.Y(n_190)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_180),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_188),
.C(n_184),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_182),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_191),
.A2(n_190),
.B(n_181),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_172),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_193),
.A2(n_14),
.B(n_15),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_16),
.Y(n_195)
);


endmodule