module fake_jpeg_28422_n_98 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_98);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_98;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_29),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_22),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_44),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_47),
.Y(n_51)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_0),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_59),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_40),
.B1(n_35),
.B2(n_34),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_54),
.B1(n_60),
.B2(n_3),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_38),
.B1(n_36),
.B2(n_33),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_56),
.Y(n_69)
);

OR2x2_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_31),
.Y(n_57)
);

AO21x1_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_3),
.B(n_4),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_41),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_58),
.B(n_2),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_1),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_15),
.B1(n_26),
.B2(n_24),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_1),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_68),
.B(n_75),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_70),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_2),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_72),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_73),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_61),
.A2(n_14),
.B1(n_21),
.B2(n_17),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_52),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_71),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_53),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_4),
.B(n_5),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_51),
.B(n_5),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_49),
.B(n_12),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_85),
.A2(n_69),
.B1(n_68),
.B2(n_78),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_88),
.B1(n_89),
.B2(n_85),
.Y(n_91)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_80),
.A2(n_71),
.B1(n_63),
.B2(n_16),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_82),
.B(n_84),
.Y(n_90)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_91),
.C(n_86),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_83),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_78),
.C(n_81),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

BUFx24_ASAP7_75t_SL g97 ( 
.A(n_96),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_13),
.Y(n_98)
);


endmodule