module fake_ariane_2045_n_108 (n_8, n_3, n_2, n_11, n_7, n_16, n_5, n_14, n_1, n_0, n_12, n_15, n_6, n_13, n_9, n_4, n_10, n_108);

input n_8;
input n_3;
input n_2;
input n_11;
input n_7;
input n_16;
input n_5;
input n_14;
input n_1;
input n_0;
input n_12;
input n_15;
input n_6;
input n_13;
input n_9;
input n_4;
input n_10;

output n_108;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_18;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_19;
wire n_40;
wire n_106;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_17;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_42;
wire n_31;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_102;
wire n_22;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

INVxp33_ASAP7_75t_SL g17 ( 
.A(n_11),
.Y(n_17)
);

INVxp67_ASAP7_75t_SL g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVxp67_ASAP7_75t_SL g22 ( 
.A(n_15),
.Y(n_22)
);

INVxp67_ASAP7_75t_SL g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVxp67_ASAP7_75t_SL g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVxp33_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVxp67_ASAP7_75t_SL g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_R g35 ( 
.A(n_24),
.B(n_8),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_29),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_27),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

AND2x4_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_19),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_27),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_18),
.B1(n_30),
.B2(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_34),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

AOI22x1_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_30),
.B1(n_25),
.B2(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_R g59 ( 
.A(n_47),
.B(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_49),
.B(n_48),
.Y(n_62)
);

AND2x4_ASAP7_75t_SL g63 ( 
.A(n_59),
.B(n_53),
.Y(n_63)
);

OAI21x1_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_46),
.B(n_34),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2x1_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_33),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_SL g67 ( 
.A(n_62),
.B(n_57),
.C(n_26),
.Y(n_67)
);

NAND2xp33_ASAP7_75t_SL g68 ( 
.A(n_65),
.B(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_65),
.B(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_63),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_50),
.C(n_58),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

NOR3xp33_ASAP7_75t_SL g79 ( 
.A(n_75),
.B(n_68),
.C(n_61),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_63),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_66),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_76),
.C(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_82),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_76),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_83),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_84),
.Y(n_95)
);

AOI211xp5_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_95),
.B(n_92),
.C(n_94),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_93),
.A2(n_40),
.B1(n_51),
.B2(n_61),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_SL g100 ( 
.A(n_96),
.B(n_40),
.C(n_61),
.Y(n_100)
);

OAI221xp5_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_23),
.B1(n_22),
.B2(n_33),
.C(n_6),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_R g102 ( 
.A(n_100),
.B(n_2),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_101),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_103),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_99),
.Y(n_105)
);

AOI221xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_102),
.B1(n_97),
.B2(n_6),
.C(n_3),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_64),
.B1(n_33),
.B2(n_4),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_64),
.B(n_4),
.Y(n_108)
);


endmodule