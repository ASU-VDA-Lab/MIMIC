module fake_netlist_6_3899_n_2060 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2060);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2060;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1888;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_76),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_58),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_1),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_131),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_13),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_106),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_150),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_148),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_32),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_193),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_166),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_182),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_6),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_171),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_135),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_138),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_102),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_31),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_67),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_90),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_58),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_80),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_205),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_61),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_86),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_139),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_96),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_179),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_130),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_198),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_177),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_202),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_126),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_137),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_120),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_93),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_4),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_85),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_29),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_64),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_95),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_161),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_178),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_51),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_114),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_208),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_71),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_105),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_65),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_40),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_197),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_123),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_6),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_49),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_206),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_209),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_162),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_68),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_133),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_169),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_207),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_192),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_10),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_187),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_170),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_203),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_11),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_20),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_183),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_60),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_160),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_62),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_10),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_77),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_136),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_60),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_36),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_180),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_176),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_154),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_204),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_13),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_22),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_144),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_8),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_153),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_103),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_63),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_88),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_84),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_155),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_5),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_132),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_212),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_181),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_141),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_16),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_56),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_189),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_89),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_140),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_17),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_149),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_185),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_73),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_4),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_104),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_2),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_2),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_54),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_81),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_75),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_83),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_33),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_79),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_23),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_53),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_151),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_36),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_30),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_74),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_158),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_175),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_51),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_1),
.Y(n_340)
);

BUFx10_ASAP7_75t_L g341 ( 
.A(n_116),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_72),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_19),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_112),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_184),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_124),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_32),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_15),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_47),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_127),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_118),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_8),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_35),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_62),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_115),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_74),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_39),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_55),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_34),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_99),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_72),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_61),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_71),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_23),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_167),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_98),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_164),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_91),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_199),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_0),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_125),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_11),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_172),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_196),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_174),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_188),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_128),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_100),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_195),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_20),
.Y(n_380)
);

BUFx10_ASAP7_75t_L g381 ( 
.A(n_18),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_146),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_38),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_194),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_77),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_50),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_190),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_92),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_65),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_121),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_75),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_82),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_54),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_24),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_59),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_14),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_107),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_69),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_0),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_40),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_83),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_200),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_68),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_41),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_108),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_17),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_152),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_101),
.Y(n_408)
);

BUFx10_ASAP7_75t_L g409 ( 
.A(n_97),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_191),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_43),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_57),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_186),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_119),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_214),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_266),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_214),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_267),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_214),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_214),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_214),
.B(n_3),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_214),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_244),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_247),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_327),
.B(n_3),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_315),
.B(n_5),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_224),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_272),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_214),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_285),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_275),
.Y(n_431)
);

NOR2xp67_ASAP7_75t_L g432 ( 
.A(n_245),
.B(n_7),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_276),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_279),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_280),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_402),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_270),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_214),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_273),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_284),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_286),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_229),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_290),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_273),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_293),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_273),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_258),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_295),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_258),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_304),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_271),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_281),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_273),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_377),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_239),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_378),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_239),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_292),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_292),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_310),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_370),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_370),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_273),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_314),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_406),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_406),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_406),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_406),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_406),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_278),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_404),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_278),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_312),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_316),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_322),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_333),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_338),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_344),
.Y(n_478)
);

CKINVDCx14_ASAP7_75t_R g479 ( 
.A(n_381),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_345),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_346),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_313),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_313),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_349),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_350),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_349),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_357),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_414),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_357),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_217),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_287),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_217),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_358),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_381),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_358),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_215),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_222),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_265),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_236),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_237),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_264),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_298),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_309),
.B(n_7),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_219),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_245),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_317),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_268),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_219),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_320),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_321),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_325),
.Y(n_511)
);

NOR2xp67_ASAP7_75t_L g512 ( 
.A(n_245),
.B(n_9),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_381),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_269),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_226),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_282),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_309),
.B(n_9),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_283),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_336),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_342),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_235),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_288),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_343),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_220),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_347),
.Y(n_525)
);

INVxp67_ASAP7_75t_SL g526 ( 
.A(n_216),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_354),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_226),
.B(n_12),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_359),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_361),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_416),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_423),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_418),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_427),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_428),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_431),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_439),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_439),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_434),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_505),
.B(n_220),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_435),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_444),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_446),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_415),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_427),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_446),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_427),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_415),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_526),
.B(n_221),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_453),
.Y(n_550)
);

CKINVDCx6p67_ASAP7_75t_R g551 ( 
.A(n_437),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_447),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_463),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_429),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_465),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_440),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_429),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_449),
.B(n_352),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_465),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_441),
.Y(n_560)
);

OA21x2_ASAP7_75t_L g561 ( 
.A1(n_421),
.A2(n_393),
.B(n_391),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_466),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_427),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_430),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_417),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_443),
.Y(n_566)
);

BUFx8_ASAP7_75t_L g567 ( 
.A(n_425),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_471),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_466),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_467),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_467),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_468),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_468),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_445),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_432),
.B(n_263),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_417),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_447),
.Y(n_577)
);

AND3x1_ASAP7_75t_L g578 ( 
.A(n_426),
.B(n_352),
.C(n_396),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_469),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_448),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_469),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_517),
.B(n_221),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_450),
.Y(n_583)
);

OA21x2_ASAP7_75t_L g584 ( 
.A1(n_419),
.A2(n_411),
.B(n_398),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_419),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_470),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_491),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_460),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_498),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_474),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_470),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_507),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_424),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_475),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_476),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_420),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_477),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_478),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_433),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_422),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_422),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_436),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_515),
.Y(n_603)
);

INVx5_ASAP7_75t_L g604 ( 
.A(n_515),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_438),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_438),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_515),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_480),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_472),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_500),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_514),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_512),
.B(n_263),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_516),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_425),
.A2(n_323),
.B1(n_326),
.B2(n_305),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_485),
.Y(n_615)
);

CKINVDCx11_ASAP7_75t_R g616 ( 
.A(n_568),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_552),
.B(n_496),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_544),
.Y(n_618)
);

AND2x6_ASAP7_75t_L g619 ( 
.A(n_575),
.B(n_294),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_561),
.A2(n_442),
.B1(n_528),
.B2(n_503),
.Y(n_620)
);

BUFx10_ASAP7_75t_L g621 ( 
.A(n_531),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_540),
.B(n_518),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_568),
.B(n_294),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_575),
.B(n_318),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_540),
.B(n_522),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_582),
.B(n_464),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_575),
.B(n_318),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_596),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_561),
.A2(n_412),
.B1(n_369),
.B2(n_525),
.Y(n_629)
);

AND2x6_ASAP7_75t_L g630 ( 
.A(n_575),
.B(n_369),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_582),
.B(n_481),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_544),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_552),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_578),
.A2(n_488),
.B1(n_492),
.B2(n_490),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_561),
.A2(n_612),
.B1(n_558),
.B2(n_584),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_577),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_577),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_596),
.B(n_521),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_600),
.B(n_521),
.Y(n_639)
);

OAI22xp33_ASAP7_75t_L g640 ( 
.A1(n_614),
.A2(n_291),
.B1(n_297),
.B2(n_289),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_544),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_600),
.B(n_360),
.Y(n_642)
);

INVxp67_ASAP7_75t_SL g643 ( 
.A(n_552),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_612),
.B(n_224),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_601),
.Y(n_645)
);

NAND2xp33_ASAP7_75t_L g646 ( 
.A(n_601),
.B(n_224),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_601),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_532),
.Y(n_648)
);

NAND3xp33_ASAP7_75t_SL g649 ( 
.A(n_614),
.B(n_508),
.C(n_504),
.Y(n_649)
);

OAI22xp33_ASAP7_75t_L g650 ( 
.A1(n_549),
.A2(n_303),
.B1(n_307),
.B2(n_300),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_558),
.B(n_366),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_612),
.B(n_455),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_601),
.Y(n_653)
);

BUFx10_ASAP7_75t_L g654 ( 
.A(n_533),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_612),
.B(n_530),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_578),
.B(n_224),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_561),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_548),
.Y(n_658)
);

INVx4_ASAP7_75t_L g659 ( 
.A(n_601),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_592),
.B(n_479),
.Y(n_660)
);

AOI22x1_ASAP7_75t_L g661 ( 
.A1(n_603),
.A2(n_458),
.B1(n_459),
.B2(n_457),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_549),
.B(n_494),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_610),
.B(n_461),
.Y(n_663)
);

AND2x2_ASAP7_75t_SL g664 ( 
.A(n_561),
.B(n_224),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_565),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_535),
.A2(n_524),
.B1(n_452),
.B2(n_454),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_567),
.B(n_231),
.Y(n_667)
);

INVxp33_ASAP7_75t_L g668 ( 
.A(n_587),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_601),
.Y(n_669)
);

BUFx10_ASAP7_75t_L g670 ( 
.A(n_536),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_610),
.B(n_462),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_576),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_584),
.A2(n_231),
.B1(n_246),
.B2(n_240),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_576),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_539),
.B(n_451),
.Y(n_675)
);

OR2x6_ASAP7_75t_L g676 ( 
.A(n_592),
.B(n_513),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_567),
.B(n_231),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_SL g678 ( 
.A(n_541),
.B(n_456),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_556),
.B(n_223),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_576),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_548),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_585),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_548),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_560),
.B(n_225),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_554),
.Y(n_685)
);

AND3x4_ASAP7_75t_L g686 ( 
.A(n_564),
.B(n_340),
.C(n_332),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_585),
.B(n_232),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_567),
.B(n_231),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_564),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_587),
.B(n_497),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_605),
.B(n_241),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_584),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_605),
.Y(n_693)
);

AND3x2_ASAP7_75t_L g694 ( 
.A(n_611),
.B(n_243),
.C(n_242),
.Y(n_694)
);

AO22x2_ASAP7_75t_L g695 ( 
.A1(n_605),
.A2(n_274),
.B1(n_277),
.B2(n_251),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_554),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_554),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_551),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_586),
.B(n_473),
.Y(n_699)
);

AND2x2_ASAP7_75t_SL g700 ( 
.A(n_584),
.B(n_231),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_606),
.B(n_299),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_584),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_557),
.Y(n_703)
);

AND2x6_ASAP7_75t_L g704 ( 
.A(n_606),
.B(n_240),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_611),
.Y(n_705)
);

BUFx10_ASAP7_75t_L g706 ( 
.A(n_566),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_534),
.B(n_301),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_534),
.Y(n_708)
);

BUFx4f_ASAP7_75t_L g709 ( 
.A(n_570),
.Y(n_709)
);

NAND2xp33_ASAP7_75t_L g710 ( 
.A(n_537),
.B(n_240),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_567),
.A2(n_410),
.B1(n_240),
.B2(n_246),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_593),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_537),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_574),
.B(n_225),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_580),
.B(n_240),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_570),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_583),
.B(n_246),
.Y(n_717)
);

INVx4_ASAP7_75t_SL g718 ( 
.A(n_571),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_557),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_538),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_SL g721 ( 
.A(n_588),
.B(n_362),
.Y(n_721)
);

INVx5_ASAP7_75t_L g722 ( 
.A(n_571),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_542),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_590),
.A2(n_261),
.B1(n_413),
.B2(n_253),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_594),
.B(n_228),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_542),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_571),
.Y(n_727)
);

INVxp67_ASAP7_75t_SL g728 ( 
.A(n_534),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_595),
.B(n_246),
.Y(n_729)
);

INVx6_ASAP7_75t_L g730 ( 
.A(n_571),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_572),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_543),
.Y(n_732)
);

AND2x2_ASAP7_75t_SL g733 ( 
.A(n_589),
.B(n_246),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_543),
.B(n_410),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_599),
.Y(n_735)
);

OAI22xp33_ASAP7_75t_SL g736 ( 
.A1(n_589),
.A2(n_262),
.B1(n_252),
.B2(n_234),
.Y(n_736)
);

AND2x6_ASAP7_75t_L g737 ( 
.A(n_546),
.B(n_410),
.Y(n_737)
);

BUFx10_ASAP7_75t_L g738 ( 
.A(n_597),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_572),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_572),
.Y(n_740)
);

BUFx8_ASAP7_75t_SL g741 ( 
.A(n_602),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_546),
.Y(n_742)
);

BUFx10_ASAP7_75t_L g743 ( 
.A(n_598),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_608),
.B(n_410),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_550),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_615),
.B(n_410),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_572),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_591),
.B(n_482),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_625),
.B(n_613),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_733),
.B(n_613),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_690),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_692),
.A2(n_392),
.B1(n_364),
.B2(n_306),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_626),
.A2(n_631),
.B1(n_733),
.B2(n_622),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_662),
.B(n_228),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_732),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_708),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_628),
.B(n_553),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_651),
.A2(n_238),
.B1(n_248),
.B2(n_230),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_636),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_705),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_692),
.A2(n_308),
.B1(n_311),
.B2(n_302),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_636),
.B(n_230),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_629),
.B(n_553),
.Y(n_763)
);

AO221x1_ASAP7_75t_L g764 ( 
.A1(n_640),
.A2(n_319),
.B1(n_376),
.B2(n_382),
.C(n_374),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_663),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_700),
.B(n_555),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_637),
.B(n_238),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_637),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_700),
.B(n_555),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_635),
.B(n_559),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_655),
.B(n_248),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_708),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_679),
.B(n_249),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_673),
.B(n_559),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_620),
.B(n_562),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_663),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_671),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_655),
.B(n_249),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_671),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_713),
.B(n_569),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_617),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_720),
.B(n_569),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_684),
.B(n_250),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_714),
.B(n_250),
.Y(n_784)
);

NOR2xp67_ASAP7_75t_L g785 ( 
.A(n_666),
.B(n_573),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_723),
.B(n_579),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_728),
.A2(n_604),
.B(n_607),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_618),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_726),
.B(n_534),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_617),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_725),
.B(n_256),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_617),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_742),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_745),
.Y(n_794)
);

INVx8_ASAP7_75t_L g795 ( 
.A(n_676),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_643),
.B(n_257),
.Y(n_796)
);

INVx8_ASAP7_75t_L g797 ( 
.A(n_676),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_745),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_656),
.B(n_715),
.Y(n_799)
);

OR2x6_ASAP7_75t_L g800 ( 
.A(n_676),
.B(n_497),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_664),
.B(n_545),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_642),
.B(n_547),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_702),
.A2(n_387),
.B(n_337),
.C(n_365),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_633),
.B(n_499),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_711),
.A2(n_384),
.B1(n_379),
.B2(n_405),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_702),
.A2(n_407),
.B1(n_356),
.B2(n_353),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_633),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_638),
.B(n_547),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_618),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_660),
.B(n_257),
.Y(n_810)
);

AND2x6_ASAP7_75t_SL g811 ( 
.A(n_676),
.B(n_499),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_667),
.A2(n_373),
.B1(n_260),
.B2(n_261),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_639),
.B(n_652),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_632),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_667),
.A2(n_375),
.B1(n_260),
.B2(n_351),
.Y(n_815)
);

OR2x6_ASAP7_75t_L g816 ( 
.A(n_677),
.B(n_501),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_689),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_652),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_715),
.B(n_351),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_699),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_621),
.Y(n_821)
);

NOR2x1p5_ASAP7_75t_L g822 ( 
.A(n_649),
.B(n_551),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_632),
.Y(n_823)
);

AND2x6_ASAP7_75t_L g824 ( 
.A(n_657),
.B(n_641),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_641),
.Y(n_825)
);

AND2x4_ASAP7_75t_SL g826 ( 
.A(n_621),
.B(n_551),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_657),
.A2(n_695),
.B1(n_630),
.B2(n_619),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_699),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_695),
.A2(n_630),
.B1(n_619),
.B2(n_627),
.Y(n_829)
);

BUFx6f_ASAP7_75t_SL g830 ( 
.A(n_621),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_650),
.B(n_355),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_630),
.B(n_563),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_741),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_630),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_658),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_717),
.B(n_355),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_681),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_717),
.B(n_729),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_729),
.B(n_367),
.Y(n_839)
);

BUFx8_ASAP7_75t_L g840 ( 
.A(n_741),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_681),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_748),
.Y(n_842)
);

INVx1_ASAP7_75t_SL g843 ( 
.A(n_616),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_661),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_683),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_683),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_744),
.B(n_367),
.Y(n_847)
);

BUFx4_ASAP7_75t_L g848 ( 
.A(n_616),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_685),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_695),
.A2(n_233),
.B1(n_213),
.B2(n_218),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_654),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_724),
.B(n_368),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_677),
.A2(n_373),
.B1(n_368),
.B2(n_371),
.Y(n_853)
);

INVxp67_ASAP7_75t_L g854 ( 
.A(n_721),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_685),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_744),
.B(n_371),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_696),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_746),
.B(n_375),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_746),
.B(n_388),
.Y(n_859)
);

AND2x2_ASAP7_75t_SL g860 ( 
.A(n_634),
.B(n_501),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_665),
.B(n_572),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_668),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_672),
.B(n_581),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_668),
.B(n_388),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_696),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_623),
.B(n_390),
.Y(n_866)
);

INVx5_ASAP7_75t_L g867 ( 
.A(n_704),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_697),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_674),
.B(n_581),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_624),
.A2(n_383),
.B1(n_218),
.B2(n_227),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_627),
.A2(n_385),
.B1(n_227),
.B2(n_233),
.Y(n_871)
);

O2A1O1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_644),
.A2(n_506),
.B(n_529),
.C(n_527),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_623),
.B(n_736),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_688),
.B(n_390),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_697),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_680),
.B(n_581),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_703),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_703),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_682),
.B(n_581),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_644),
.A2(n_385),
.B1(n_234),
.B2(n_252),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_688),
.B(n_397),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_799),
.B(n_654),
.Y(n_882)
);

INVx4_ASAP7_75t_L g883 ( 
.A(n_807),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_770),
.A2(n_709),
.B(n_653),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_775),
.A2(n_653),
.B(n_645),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_799),
.A2(n_675),
.B(n_687),
.C(n_691),
.Y(n_886)
);

A2O1A1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_838),
.A2(n_701),
.B(n_510),
.C(n_511),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_756),
.Y(n_888)
);

BUFx10_ASAP7_75t_L g889 ( 
.A(n_830),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_813),
.B(n_693),
.Y(n_890)
);

AO21x1_ASAP7_75t_L g891 ( 
.A1(n_838),
.A2(n_707),
.B(n_646),
.Y(n_891)
);

INVx3_ASAP7_75t_SL g892 ( 
.A(n_826),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_773),
.B(n_719),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_756),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_755),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_773),
.B(n_719),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_783),
.B(n_716),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_SL g898 ( 
.A(n_830),
.B(n_654),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_784),
.B(n_727),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_766),
.A2(n_659),
.B(n_645),
.Y(n_900)
);

A2O1A1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_752),
.A2(n_502),
.B(n_506),
.C(n_509),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_749),
.B(n_751),
.Y(n_902)
);

NOR3xp33_ASAP7_75t_L g903 ( 
.A(n_750),
.B(n_712),
.C(n_648),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_755),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_L g905 ( 
.A1(n_761),
.A2(n_686),
.B1(n_659),
.B2(n_669),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_818),
.B(n_694),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_862),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_808),
.A2(n_659),
.B(n_647),
.Y(n_908)
);

INVx1_ASAP7_75t_SL g909 ( 
.A(n_760),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_802),
.A2(n_669),
.B(n_647),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_817),
.Y(n_911)
);

O2A1O1Ixp33_ASAP7_75t_SL g912 ( 
.A1(n_803),
.A2(n_502),
.B(n_527),
.C(n_523),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_806),
.A2(n_646),
.B(n_710),
.C(n_734),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_840),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_759),
.Y(n_915)
);

OAI21xp33_ASAP7_75t_L g916 ( 
.A1(n_754),
.A2(n_678),
.B(n_254),
.Y(n_916)
);

OAI21xp33_ASAP7_75t_L g917 ( 
.A1(n_754),
.A2(n_254),
.B(n_213),
.Y(n_917)
);

OAI21xp5_ASAP7_75t_L g918 ( 
.A1(n_769),
.A2(n_761),
.B(n_763),
.Y(n_918)
);

INVx11_ASAP7_75t_L g919 ( 
.A(n_840),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_874),
.A2(n_731),
.B(n_740),
.C(n_413),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_806),
.A2(n_710),
.B(n_734),
.C(n_519),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_873),
.A2(n_791),
.B1(n_881),
.B2(n_874),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_881),
.A2(n_731),
.B(n_740),
.C(n_408),
.Y(n_923)
);

AOI21x1_ASAP7_75t_L g924 ( 
.A1(n_787),
.A2(n_609),
.B(n_483),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_768),
.Y(n_925)
);

AOI21x1_ASAP7_75t_L g926 ( 
.A1(n_789),
.A2(n_609),
.B(n_483),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_752),
.A2(n_686),
.B1(n_408),
.B2(n_397),
.Y(n_927)
);

OR2x6_ASAP7_75t_L g928 ( 
.A(n_795),
.B(n_670),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_873),
.A2(n_670),
.B1(n_743),
.B2(n_706),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_764),
.A2(n_400),
.B1(n_255),
.B2(n_259),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_831),
.A2(n_805),
.B(n_776),
.C(n_777),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_793),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_794),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_834),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_762),
.B(n_670),
.Y(n_935)
);

AOI21xp33_ASAP7_75t_L g936 ( 
.A1(n_819),
.A2(n_735),
.B(n_698),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_765),
.A2(n_523),
.B(n_520),
.C(n_519),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_779),
.A2(n_520),
.B(n_511),
.C(n_510),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_820),
.B(n_828),
.Y(n_939)
);

AO32x2_ASAP7_75t_L g940 ( 
.A1(n_827),
.A2(n_737),
.A3(n_383),
.B1(n_380),
.B2(n_372),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_832),
.A2(n_747),
.B(n_739),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_772),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_798),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_774),
.A2(n_704),
.B(n_737),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_798),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_827),
.A2(n_829),
.B1(n_781),
.B2(n_792),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_829),
.B(n_706),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_819),
.A2(n_698),
.B(n_509),
.C(n_331),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_772),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_762),
.B(n_706),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_844),
.A2(n_824),
.B(n_814),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_821),
.Y(n_952)
);

OAI21xp33_ASAP7_75t_L g953 ( 
.A1(n_870),
.A2(n_356),
.B(n_255),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_861),
.A2(n_722),
.B(n_604),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_800),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_854),
.B(n_738),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_863),
.A2(n_722),
.B(n_604),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_790),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_821),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_869),
.A2(n_722),
.B(n_604),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_842),
.A2(n_495),
.B(n_493),
.C(n_482),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_876),
.A2(n_722),
.B(n_604),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_879),
.A2(n_581),
.B(n_718),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_836),
.A2(n_324),
.B(n_328),
.C(n_329),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_757),
.A2(n_581),
.B(n_718),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_824),
.A2(n_823),
.B(n_809),
.Y(n_966)
);

BUFx12f_ASAP7_75t_L g967 ( 
.A(n_811),
.Y(n_967)
);

INVx6_ASAP7_75t_L g968 ( 
.A(n_807),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_780),
.A2(n_718),
.B(n_730),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_782),
.A2(n_718),
.B(n_495),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_860),
.B(n_738),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_836),
.A2(n_743),
.B1(n_738),
.B2(n_737),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_823),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_816),
.A2(n_859),
.B1(n_858),
.B2(n_847),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_804),
.Y(n_975)
);

O2A1O1Ixp5_ASAP7_75t_SL g976 ( 
.A1(n_856),
.A2(n_486),
.B(n_493),
.C(n_489),
.Y(n_976)
);

OAI21xp33_ASAP7_75t_L g977 ( 
.A1(n_870),
.A2(n_353),
.B(n_262),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_839),
.A2(n_330),
.B(n_334),
.C(n_335),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_825),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_839),
.A2(n_372),
.B(n_403),
.C(n_401),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_796),
.B(n_743),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_786),
.A2(n_487),
.B(n_484),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_847),
.A2(n_737),
.B1(n_704),
.B2(n_235),
.Y(n_983)
);

AOI21x1_ASAP7_75t_L g984 ( 
.A1(n_846),
.A2(n_487),
.B(n_484),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_834),
.B(n_235),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_824),
.A2(n_704),
.B(n_348),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_860),
.B(n_858),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_851),
.Y(n_988)
);

OAI21x1_ASAP7_75t_L g989 ( 
.A1(n_825),
.A2(n_704),
.B(n_87),
.Y(n_989)
);

NAND2x1_ASAP7_75t_L g990 ( 
.A(n_834),
.B(n_94),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_852),
.B(n_339),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_804),
.B(n_259),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_851),
.B(n_363),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_800),
.Y(n_994)
);

NOR2x1_ASAP7_75t_L g995 ( 
.A(n_822),
.B(n_296),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_807),
.B(n_363),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_834),
.A2(n_788),
.B(n_835),
.Y(n_997)
);

NOR2x1p5_ASAP7_75t_SL g998 ( 
.A(n_837),
.B(n_296),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_807),
.B(n_296),
.Y(n_999)
);

NOR2x1_ASAP7_75t_L g1000 ( 
.A(n_816),
.B(n_341),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_845),
.B(n_380),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_767),
.B(n_386),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_785),
.B(n_109),
.Y(n_1003)
);

OAI21x1_ASAP7_75t_L g1004 ( 
.A1(n_845),
.A2(n_156),
.B(n_111),
.Y(n_1004)
);

BUFx8_ASAP7_75t_L g1005 ( 
.A(n_848),
.Y(n_1005)
);

BUFx12f_ASAP7_75t_L g1006 ( 
.A(n_833),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_864),
.B(n_386),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_841),
.A2(n_389),
.B(n_403),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_758),
.A2(n_395),
.B(n_401),
.C(n_400),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_865),
.B(n_868),
.Y(n_1010)
);

AOI21x1_ASAP7_75t_L g1011 ( 
.A1(n_849),
.A2(n_409),
.B(n_341),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_816),
.A2(n_409),
.B1(n_341),
.B2(n_395),
.Y(n_1012)
);

AO21x1_ASAP7_75t_L g1013 ( 
.A1(n_855),
.A2(n_409),
.B(n_15),
.Y(n_1013)
);

BUFx12f_ASAP7_75t_L g1014 ( 
.A(n_800),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_857),
.A2(n_399),
.B(n_394),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_826),
.Y(n_1016)
);

NAND2xp33_ASAP7_75t_L g1017 ( 
.A(n_867),
.B(n_389),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_875),
.A2(n_399),
.B(n_394),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_880),
.A2(n_201),
.B1(n_173),
.B2(n_168),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_771),
.B(n_163),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_795),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_872),
.A2(n_14),
.B(n_16),
.C(n_18),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_871),
.B(n_19),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_868),
.B(n_21),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_877),
.B(n_21),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_877),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_878),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_866),
.B(n_810),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_902),
.B(n_935),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_973),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_987),
.B(n_778),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_919),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_966),
.A2(n_850),
.B(n_812),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_987),
.B(n_880),
.Y(n_1034)
);

OAI21x1_ASAP7_75t_L g1035 ( 
.A1(n_908),
.A2(n_850),
.B(n_815),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_895),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_902),
.B(n_871),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_950),
.B(n_843),
.Y(n_1038)
);

OAI22x1_ASAP7_75t_L g1039 ( 
.A1(n_1012),
.A2(n_853),
.B1(n_797),
.B2(n_25),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_907),
.B(n_797),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_904),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_934),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_993),
.B(n_22),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_909),
.Y(n_1044)
);

OR2x6_ASAP7_75t_SL g1045 ( 
.A(n_927),
.B(n_24),
.Y(n_1045)
);

NOR2xp67_ASAP7_75t_L g1046 ( 
.A(n_929),
.B(n_143),
.Y(n_1046)
);

AOI21xp33_ASAP7_75t_L g1047 ( 
.A1(n_974),
.A2(n_25),
.B(n_26),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_910),
.A2(n_867),
.B(n_159),
.Y(n_1048)
);

INVx5_ASAP7_75t_L g1049 ( 
.A(n_934),
.Y(n_1049)
);

AOI21x1_ASAP7_75t_L g1050 ( 
.A1(n_897),
.A2(n_157),
.B(n_147),
.Y(n_1050)
);

AO31x2_ASAP7_75t_L g1051 ( 
.A1(n_891),
.A2(n_26),
.A3(n_27),
.B(n_28),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_951),
.A2(n_145),
.B(n_142),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_901),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_1053)
);

AO31x2_ASAP7_75t_L g1054 ( 
.A1(n_887),
.A2(n_31),
.A3(n_33),
.B(n_34),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_886),
.A2(n_134),
.B(n_129),
.Y(n_1055)
);

NOR2x1_ASAP7_75t_R g1056 ( 
.A(n_1006),
.B(n_35),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_941),
.A2(n_122),
.B(n_117),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_947),
.A2(n_113),
.B1(n_110),
.B2(n_39),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_1004),
.A2(n_37),
.B(n_38),
.Y(n_1059)
);

NAND2x1p5_ASAP7_75t_L g1060 ( 
.A(n_883),
.B(n_37),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_975),
.B(n_42),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_893),
.A2(n_42),
.B(n_43),
.Y(n_1062)
);

AOI21xp33_ASAP7_75t_L g1063 ( 
.A1(n_991),
.A2(n_44),
.B(n_45),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_884),
.A2(n_44),
.B(n_46),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_896),
.A2(n_46),
.B(n_47),
.Y(n_1065)
);

AO21x1_ASAP7_75t_L g1066 ( 
.A1(n_1019),
.A2(n_48),
.B(n_49),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_939),
.B(n_48),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_971),
.A2(n_84),
.B1(n_52),
.B2(n_53),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_890),
.B(n_50),
.Y(n_1069)
);

OAI22x1_ASAP7_75t_L g1070 ( 
.A1(n_1023),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_975),
.B(n_66),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_914),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_981),
.B(n_69),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_920),
.A2(n_70),
.B(n_73),
.Y(n_1074)
);

OR2x6_ASAP7_75t_L g1075 ( 
.A(n_928),
.B(n_1014),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_923),
.A2(n_70),
.B(n_76),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_899),
.A2(n_78),
.B(n_79),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_911),
.B(n_971),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_958),
.B(n_882),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_882),
.B(n_901),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_934),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_1020),
.B(n_947),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_911),
.B(n_996),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1028),
.B(n_1020),
.Y(n_1084)
);

NOR2xp67_ASAP7_75t_L g1085 ( 
.A(n_956),
.B(n_1021),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_924),
.A2(n_997),
.B(n_989),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_933),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_887),
.A2(n_946),
.B(n_931),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_959),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_934),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1028),
.A2(n_991),
.B1(n_903),
.B2(n_916),
.Y(n_1091)
);

OAI21xp33_ASAP7_75t_L g1092 ( 
.A1(n_917),
.A2(n_1002),
.B(n_953),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_945),
.Y(n_1093)
);

OR2x6_ASAP7_75t_L g1094 ( 
.A(n_928),
.B(n_1021),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1001),
.B(n_888),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_888),
.B(n_894),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_968),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_926),
.A2(n_963),
.B(n_984),
.Y(n_1098)
);

AO31x2_ASAP7_75t_L g1099 ( 
.A1(n_1013),
.A2(n_1022),
.A3(n_905),
.B(n_980),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_1005),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_894),
.B(n_942),
.Y(n_1101)
);

AOI21x1_ASAP7_75t_SL g1102 ( 
.A1(n_1024),
.A2(n_1025),
.B(n_1003),
.Y(n_1102)
);

NAND2x1p5_ASAP7_75t_L g1103 ( 
.A(n_883),
.B(n_942),
.Y(n_1103)
);

OR2x6_ASAP7_75t_L g1104 ( 
.A(n_928),
.B(n_955),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_1010),
.A2(n_969),
.B(n_965),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_949),
.B(n_1002),
.Y(n_1106)
);

NAND2x1p5_ASAP7_75t_L g1107 ( 
.A(n_990),
.B(n_988),
.Y(n_1107)
);

AOI21x1_ASAP7_75t_L g1108 ( 
.A1(n_979),
.A2(n_1026),
.B(n_985),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_936),
.B(n_956),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_976),
.A2(n_944),
.B(n_913),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1007),
.B(n_925),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_970),
.A2(n_954),
.B(n_962),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_1005),
.Y(n_1113)
);

INVx2_ASAP7_75t_SL g1114 ( 
.A(n_915),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_957),
.A2(n_960),
.B(n_943),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_892),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1007),
.B(n_925),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_977),
.A2(n_930),
.B1(n_1003),
.B2(n_932),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_915),
.B(n_992),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1027),
.B(n_980),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_948),
.A2(n_964),
.B(n_978),
.C(n_938),
.Y(n_1121)
);

AOI21x1_ASAP7_75t_L g1122 ( 
.A1(n_999),
.A2(n_986),
.B(n_1011),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_921),
.A2(n_961),
.B(n_999),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_937),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_968),
.Y(n_1125)
);

INVx5_ASAP7_75t_L g1126 ( 
.A(n_968),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1009),
.A2(n_972),
.B(n_983),
.Y(n_1127)
);

INVxp67_ASAP7_75t_SL g1128 ( 
.A(n_994),
.Y(n_1128)
);

AOI21xp33_ASAP7_75t_L g1129 ( 
.A1(n_952),
.A2(n_1000),
.B(n_994),
.Y(n_1129)
);

INVxp67_ASAP7_75t_L g1130 ( 
.A(n_906),
.Y(n_1130)
);

AOI221xp5_ASAP7_75t_SL g1131 ( 
.A1(n_1018),
.A2(n_930),
.B1(n_1015),
.B2(n_1008),
.C(n_1017),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_906),
.B(n_903),
.Y(n_1132)
);

AO31x2_ASAP7_75t_L g1133 ( 
.A1(n_982),
.A2(n_940),
.A3(n_912),
.B(n_998),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_912),
.A2(n_995),
.B(n_1016),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_892),
.B(n_898),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_940),
.A2(n_889),
.B(n_967),
.C(n_987),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_940),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_940),
.A2(n_900),
.B(n_885),
.Y(n_1138)
);

NAND3xp33_ASAP7_75t_L g1139 ( 
.A(n_889),
.B(n_987),
.C(n_922),
.Y(n_1139)
);

INVxp67_ASAP7_75t_L g1140 ( 
.A(n_907),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_934),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_922),
.B(n_753),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_951),
.A2(n_1004),
.B(n_989),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_922),
.B(n_753),
.Y(n_1144)
);

BUFx4f_ASAP7_75t_L g1145 ( 
.A(n_892),
.Y(n_1145)
);

CKINVDCx11_ASAP7_75t_R g1146 ( 
.A(n_914),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_973),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_895),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_895),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_918),
.A2(n_922),
.B(n_801),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_907),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_934),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_922),
.A2(n_987),
.B1(n_753),
.B2(n_974),
.Y(n_1153)
);

AND2x2_ASAP7_75t_SL g1154 ( 
.A(n_987),
.B(n_922),
.Y(n_1154)
);

O2A1O1Ixp5_ASAP7_75t_L g1155 ( 
.A1(n_974),
.A2(n_891),
.B(n_987),
.C(n_887),
.Y(n_1155)
);

AO31x2_ASAP7_75t_L g1156 ( 
.A1(n_891),
.A2(n_887),
.A3(n_923),
.B(n_920),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_895),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_922),
.B(n_753),
.Y(n_1158)
);

AOI21xp33_ASAP7_75t_L g1159 ( 
.A1(n_922),
.A2(n_987),
.B(n_974),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_934),
.Y(n_1160)
);

BUFx8_ASAP7_75t_SL g1161 ( 
.A(n_914),
.Y(n_1161)
);

NOR2x1_ASAP7_75t_SL g1162 ( 
.A(n_934),
.B(n_834),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1109),
.B(n_1029),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1094),
.B(n_1130),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_1094),
.B(n_1130),
.Y(n_1165)
);

OAI21xp33_ASAP7_75t_L g1166 ( 
.A1(n_1092),
.A2(n_1031),
.B(n_1034),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_1094),
.B(n_1089),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1154),
.A2(n_1158),
.B1(n_1144),
.B2(n_1142),
.Y(n_1168)
);

INVx3_ASAP7_75t_SL g1169 ( 
.A(n_1032),
.Y(n_1169)
);

HB1xp67_ASAP7_75t_L g1170 ( 
.A(n_1044),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1031),
.B(n_1109),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1111),
.B(n_1117),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1036),
.Y(n_1173)
);

INVx3_ASAP7_75t_SL g1174 ( 
.A(n_1032),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_1089),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1041),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1030),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1081),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1154),
.B(n_1153),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_1126),
.Y(n_1180)
);

OA21x2_ASAP7_75t_L g1181 ( 
.A1(n_1138),
.A2(n_1110),
.B(n_1088),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_1081),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_1145),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_1084),
.B(n_1139),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_1081),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_1140),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1086),
.A2(n_1105),
.B(n_1143),
.Y(n_1187)
);

BUFx2_ASAP7_75t_SL g1188 ( 
.A(n_1126),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1119),
.B(n_1043),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1159),
.B(n_1150),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1037),
.A2(n_1091),
.B1(n_1082),
.B2(n_1118),
.Y(n_1191)
);

OR2x6_ASAP7_75t_SL g1192 ( 
.A(n_1072),
.B(n_1116),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1073),
.B(n_1106),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1073),
.B(n_1078),
.Y(n_1194)
);

BUFx10_ASAP7_75t_L g1195 ( 
.A(n_1072),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1038),
.B(n_1061),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_1114),
.Y(n_1197)
);

NAND2x1p5_ASAP7_75t_L g1198 ( 
.A(n_1049),
.B(n_1126),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1087),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1078),
.B(n_1083),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_1040),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1067),
.B(n_1069),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1118),
.A2(n_1136),
.B1(n_1055),
.B2(n_1065),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1140),
.B(n_1151),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1093),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1148),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_1126),
.Y(n_1207)
);

NOR2x1_ASAP7_75t_L g1208 ( 
.A(n_1085),
.B(n_1097),
.Y(n_1208)
);

NOR3xp33_ASAP7_75t_L g1209 ( 
.A(n_1063),
.B(n_1129),
.C(n_1047),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1081),
.Y(n_1210)
);

INVx3_ASAP7_75t_SL g1211 ( 
.A(n_1116),
.Y(n_1211)
);

O2A1O1Ixp5_ASAP7_75t_L g1212 ( 
.A1(n_1066),
.A2(n_1127),
.B(n_1155),
.C(n_1076),
.Y(n_1212)
);

OR2x6_ASAP7_75t_L g1213 ( 
.A(n_1104),
.B(n_1075),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1079),
.B(n_1095),
.Y(n_1214)
);

AND2x6_ASAP7_75t_L g1215 ( 
.A(n_1141),
.B(n_1152),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1121),
.A2(n_1155),
.B(n_1035),
.C(n_1033),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1141),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_1141),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1145),
.Y(n_1219)
);

BUFx2_ASAP7_75t_R g1220 ( 
.A(n_1161),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_SL g1221 ( 
.A1(n_1062),
.A2(n_1077),
.B(n_1074),
.C(n_1132),
.Y(n_1221)
);

INVxp67_ASAP7_75t_SL g1222 ( 
.A(n_1151),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_SL g1223 ( 
.A1(n_1132),
.A2(n_1058),
.B1(n_1135),
.B2(n_1128),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1149),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1124),
.B(n_1080),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1157),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1104),
.B(n_1075),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1071),
.B(n_1120),
.Y(n_1228)
);

INVx1_ASAP7_75t_SL g1229 ( 
.A(n_1125),
.Y(n_1229)
);

INVx1_ASAP7_75t_SL g1230 ( 
.A(n_1125),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1147),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1053),
.A2(n_1121),
.B(n_1136),
.C(n_1128),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_SL g1233 ( 
.A1(n_1134),
.A2(n_1064),
.B(n_1162),
.Y(n_1233)
);

INVx1_ASAP7_75t_SL g1234 ( 
.A(n_1125),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1103),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1039),
.A2(n_1046),
.B1(n_1131),
.B2(n_1068),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1104),
.A2(n_1070),
.B1(n_1075),
.B2(n_1107),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1045),
.B(n_1060),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1125),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1141),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1137),
.A2(n_1101),
.B1(n_1096),
.B2(n_1060),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1103),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1053),
.A2(n_1049),
.B1(n_1152),
.B2(n_1107),
.Y(n_1243)
);

OR2x6_ASAP7_75t_SL g1244 ( 
.A(n_1100),
.B(n_1161),
.Y(n_1244)
);

BUFx4_ASAP7_75t_SL g1245 ( 
.A(n_1113),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1097),
.B(n_1049),
.Y(n_1246)
);

NAND3xp33_ASAP7_75t_L g1247 ( 
.A(n_1152),
.B(n_1160),
.C(n_1090),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1123),
.A2(n_1146),
.B1(n_1042),
.B2(n_1090),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1100),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1042),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1143),
.A2(n_1123),
.B(n_1115),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1112),
.A2(n_1048),
.B(n_1057),
.Y(n_1252)
);

AND2x6_ASAP7_75t_L g1253 ( 
.A(n_1152),
.B(n_1160),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1099),
.B(n_1156),
.Y(n_1254)
);

BUFx12f_ASAP7_75t_L g1255 ( 
.A(n_1146),
.Y(n_1255)
);

OAI21xp33_ASAP7_75t_L g1256 ( 
.A1(n_1122),
.A2(n_1113),
.B(n_1108),
.Y(n_1256)
);

BUFx2_ASAP7_75t_SL g1257 ( 
.A(n_1056),
.Y(n_1257)
);

O2A1O1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1099),
.A2(n_1102),
.B(n_1156),
.C(n_1054),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1050),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1156),
.B(n_1133),
.Y(n_1260)
);

BUFx12f_ASAP7_75t_L g1261 ( 
.A(n_1054),
.Y(n_1261)
);

CKINVDCx16_ASAP7_75t_R g1262 ( 
.A(n_1102),
.Y(n_1262)
);

NAND3xp33_ASAP7_75t_L g1263 ( 
.A(n_1156),
.B(n_1054),
.C(n_1051),
.Y(n_1263)
);

NAND2x1p5_ASAP7_75t_L g1264 ( 
.A(n_1052),
.B(n_1059),
.Y(n_1264)
);

AOI221xp5_ASAP7_75t_L g1265 ( 
.A1(n_1051),
.A2(n_1052),
.B1(n_1133),
.B2(n_1059),
.C(n_1098),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1133),
.B(n_1051),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1098),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1142),
.B(n_1144),
.Y(n_1268)
);

OR2x6_ASAP7_75t_L g1269 ( 
.A(n_1104),
.B(n_1075),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1154),
.A2(n_922),
.B1(n_1034),
.B2(n_987),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1142),
.B(n_1144),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1126),
.Y(n_1272)
);

AOI222xp33_ASAP7_75t_L g1273 ( 
.A1(n_1154),
.A2(n_1023),
.B1(n_1034),
.B2(n_1153),
.C1(n_987),
.C2(n_953),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1142),
.B(n_1144),
.Y(n_1274)
);

INVxp33_ASAP7_75t_L g1275 ( 
.A(n_1044),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1089),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1031),
.A2(n_987),
.B1(n_922),
.B2(n_424),
.Y(n_1277)
);

O2A1O1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1159),
.A2(n_749),
.B(n_987),
.C(n_974),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1036),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1142),
.B(n_1144),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1142),
.B(n_1144),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_SL g1282 ( 
.A(n_1159),
.B(n_987),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1030),
.Y(n_1283)
);

NOR2xp67_ASAP7_75t_L g1284 ( 
.A(n_1140),
.B(n_1151),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1084),
.B(n_648),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1029),
.B(n_1111),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1142),
.B(n_1144),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1029),
.B(n_1031),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1044),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1031),
.B(n_749),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1154),
.A2(n_922),
.B1(n_1034),
.B2(n_987),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1161),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1044),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1159),
.A2(n_987),
.B(n_922),
.C(n_753),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1036),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1089),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1126),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_SL g1298 ( 
.A(n_1159),
.B(n_987),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1154),
.A2(n_922),
.B1(n_1034),
.B2(n_987),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1029),
.B(n_1031),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1029),
.B(n_1031),
.Y(n_1301)
);

NAND2x1_ASAP7_75t_L g1302 ( 
.A(n_1081),
.B(n_968),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1044),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1142),
.B(n_1144),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1094),
.B(n_1021),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1030),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1029),
.B(n_1111),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1126),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1036),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1044),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1159),
.A2(n_987),
.B1(n_1154),
.B2(n_1153),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1142),
.B(n_1144),
.Y(n_1312)
);

OR2x6_ASAP7_75t_L g1313 ( 
.A(n_1104),
.B(n_1075),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1142),
.B(n_1144),
.Y(n_1314)
);

CKINVDCx11_ASAP7_75t_R g1315 ( 
.A(n_1244),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1251),
.A2(n_1252),
.B(n_1187),
.Y(n_1316)
);

OAI21xp33_ASAP7_75t_L g1317 ( 
.A1(n_1290),
.A2(n_1171),
.B(n_1277),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1176),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1186),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1273),
.B(n_1268),
.Y(n_1320)
);

OAI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1282),
.A2(n_1298),
.B1(n_1194),
.B2(n_1237),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1245),
.Y(n_1322)
);

OA21x2_ASAP7_75t_L g1323 ( 
.A1(n_1212),
.A2(n_1265),
.B(n_1216),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1311),
.A2(n_1294),
.B1(n_1200),
.B2(n_1223),
.Y(n_1324)
);

AO21x1_ASAP7_75t_SL g1325 ( 
.A1(n_1236),
.A2(n_1202),
.B(n_1254),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1170),
.Y(n_1326)
);

AO21x1_ASAP7_75t_SL g1327 ( 
.A1(n_1266),
.A2(n_1254),
.B(n_1260),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1199),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1278),
.A2(n_1190),
.B(n_1282),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_SL g1330 ( 
.A1(n_1184),
.A2(n_1213),
.B1(n_1313),
.B2(n_1269),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1205),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1206),
.Y(n_1332)
);

INVxp67_ASAP7_75t_SL g1333 ( 
.A(n_1222),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1198),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1198),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1209),
.A2(n_1273),
.B1(n_1299),
.B2(n_1270),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1224),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_1293),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1226),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1279),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1175),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1295),
.Y(n_1342)
);

INVxp33_ASAP7_75t_L g1343 ( 
.A(n_1289),
.Y(n_1343)
);

INVxp67_ASAP7_75t_L g1344 ( 
.A(n_1303),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1309),
.Y(n_1345)
);

BUFx12f_ASAP7_75t_L g1346 ( 
.A(n_1255),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1231),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1298),
.A2(n_1238),
.B1(n_1203),
.B2(n_1299),
.Y(n_1348)
);

BUFx12f_ASAP7_75t_L g1349 ( 
.A(n_1292),
.Y(n_1349)
);

AO21x1_ASAP7_75t_L g1350 ( 
.A1(n_1203),
.A2(n_1191),
.B(n_1190),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1283),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1310),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1268),
.B(n_1271),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1271),
.B(n_1274),
.Y(n_1354)
);

BUFx8_ASAP7_75t_L g1355 ( 
.A(n_1249),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_SL g1356 ( 
.A1(n_1270),
.A2(n_1291),
.B1(n_1191),
.B2(n_1179),
.Y(n_1356)
);

CKINVDCx6p67_ASAP7_75t_R g1357 ( 
.A(n_1169),
.Y(n_1357)
);

BUFx8_ASAP7_75t_SL g1358 ( 
.A(n_1183),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1180),
.Y(n_1359)
);

BUFx8_ASAP7_75t_SL g1360 ( 
.A(n_1219),
.Y(n_1360)
);

BUFx12f_ASAP7_75t_L g1361 ( 
.A(n_1195),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1306),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_SL g1363 ( 
.A1(n_1291),
.A2(n_1179),
.B1(n_1168),
.B2(n_1301),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1274),
.A2(n_1314),
.B1(n_1312),
.B2(n_1304),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1250),
.Y(n_1365)
);

NAND2x1_ASAP7_75t_L g1366 ( 
.A(n_1233),
.B(n_1215),
.Y(n_1366)
);

CKINVDCx20_ASAP7_75t_R g1367 ( 
.A(n_1174),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1225),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_1180),
.Y(n_1369)
);

INVx5_ASAP7_75t_L g1370 ( 
.A(n_1215),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1280),
.B(n_1281),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_1180),
.Y(n_1372)
);

AO21x1_ASAP7_75t_L g1373 ( 
.A1(n_1232),
.A2(n_1258),
.B(n_1168),
.Y(n_1373)
);

NAND2x1p5_ASAP7_75t_L g1374 ( 
.A(n_1207),
.B(n_1272),
.Y(n_1374)
);

AO21x1_ASAP7_75t_SL g1375 ( 
.A1(n_1266),
.A2(n_1260),
.B(n_1312),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1166),
.A2(n_1163),
.B1(n_1314),
.B2(n_1287),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1280),
.B(n_1281),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1181),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1204),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_1207),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1286),
.Y(n_1381)
);

CKINVDCx11_ASAP7_75t_R g1382 ( 
.A(n_1192),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1287),
.A2(n_1304),
.B1(n_1300),
.B2(n_1288),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1307),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1214),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1193),
.A2(n_1196),
.B1(n_1285),
.B2(n_1189),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1172),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1228),
.B(n_1284),
.Y(n_1388)
);

INVx5_ASAP7_75t_L g1389 ( 
.A(n_1215),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1272),
.B(n_1297),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1197),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1178),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1201),
.A2(n_1241),
.B1(n_1248),
.B2(n_1275),
.Y(n_1393)
);

INVx6_ASAP7_75t_L g1394 ( 
.A(n_1272),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_SL g1395 ( 
.A1(n_1227),
.A2(n_1261),
.B1(n_1243),
.B2(n_1164),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1178),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1164),
.A2(n_1165),
.B1(n_1313),
.B2(n_1213),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1276),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1227),
.A2(n_1313),
.B1(n_1269),
.B2(n_1213),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1165),
.A2(n_1269),
.B1(n_1262),
.B2(n_1305),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1256),
.A2(n_1243),
.B1(n_1167),
.B2(n_1195),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1182),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_1211),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_1257),
.Y(n_1404)
);

INVx1_ASAP7_75t_SL g1405 ( 
.A(n_1296),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1235),
.B(n_1242),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1305),
.B(n_1167),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1221),
.A2(n_1263),
.B1(n_1208),
.B2(n_1239),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1267),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1182),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1185),
.B(n_1210),
.Y(n_1411)
);

INVx6_ASAP7_75t_L g1412 ( 
.A(n_1297),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1215),
.Y(n_1413)
);

AOI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1263),
.A2(n_1247),
.B(n_1302),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1220),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1210),
.Y(n_1416)
);

INVx6_ASAP7_75t_L g1417 ( 
.A(n_1297),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1188),
.A2(n_1247),
.B1(n_1308),
.B2(n_1229),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1264),
.B(n_1229),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_SL g1420 ( 
.A1(n_1230),
.A2(n_1234),
.B1(n_1308),
.B2(n_1239),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1217),
.A2(n_1218),
.B(n_1259),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1217),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1230),
.A2(n_1234),
.B1(n_1246),
.B2(n_1218),
.Y(n_1423)
);

AOI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1259),
.A2(n_1253),
.B(n_1240),
.Y(n_1424)
);

INVx6_ASAP7_75t_L g1425 ( 
.A(n_1240),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1253),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1253),
.Y(n_1427)
);

AO21x1_ASAP7_75t_L g1428 ( 
.A1(n_1253),
.A2(n_1203),
.B(n_1153),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1292),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1171),
.A2(n_987),
.B1(n_1154),
.B2(n_1159),
.Y(n_1430)
);

CKINVDCx8_ASAP7_75t_R g1431 ( 
.A(n_1188),
.Y(n_1431)
);

AO21x1_ASAP7_75t_L g1432 ( 
.A1(n_1203),
.A2(n_1153),
.B(n_1278),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1173),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_1292),
.Y(n_1434)
);

NAND3xp33_ASAP7_75t_SL g1435 ( 
.A(n_1290),
.B(n_749),
.C(n_753),
.Y(n_1435)
);

CKINVDCx6p67_ASAP7_75t_R g1436 ( 
.A(n_1255),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1173),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1173),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1277),
.A2(n_1290),
.B1(n_922),
.B2(n_1171),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1173),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1212),
.A2(n_1265),
.B(n_1138),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1173),
.Y(n_1442)
);

BUFx4f_ASAP7_75t_L g1443 ( 
.A(n_1180),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1251),
.A2(n_1252),
.B(n_1187),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1177),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1273),
.B(n_1154),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1171),
.A2(n_987),
.B1(n_1154),
.B2(n_1159),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1290),
.B(n_1171),
.Y(n_1448)
);

CKINVDCx11_ASAP7_75t_R g1449 ( 
.A(n_1244),
.Y(n_1449)
);

INVx4_ASAP7_75t_L g1450 ( 
.A(n_1180),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1273),
.B(n_1154),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1175),
.Y(n_1452)
);

INVx3_ASAP7_75t_L g1453 ( 
.A(n_1198),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1277),
.A2(n_1290),
.B1(n_922),
.B2(n_1171),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1173),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1173),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1171),
.A2(n_987),
.B1(n_1154),
.B2(n_1159),
.Y(n_1457)
);

NOR2x1_ASAP7_75t_R g1458 ( 
.A(n_1255),
.B(n_616),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1171),
.A2(n_987),
.B1(n_1290),
.B2(n_1154),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1273),
.B(n_1154),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1186),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1277),
.A2(n_1290),
.B1(n_922),
.B2(n_1171),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1198),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1173),
.Y(n_1464)
);

BUFx2_ASAP7_75t_R g1465 ( 
.A(n_1244),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1171),
.A2(n_987),
.B1(n_1154),
.B2(n_1159),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1170),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1179),
.B(n_1270),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1173),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1173),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1173),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1173),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1448),
.B(n_1383),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1352),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1366),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1371),
.B(n_1377),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1371),
.B(n_1377),
.Y(n_1477)
);

AO21x2_ASAP7_75t_L g1478 ( 
.A1(n_1329),
.A2(n_1444),
.B(n_1316),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_1352),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1317),
.B(n_1353),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1439),
.B(n_1454),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1378),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1354),
.B(n_1385),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1419),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1413),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1373),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1373),
.Y(n_1487)
);

INVx5_ASAP7_75t_L g1488 ( 
.A(n_1370),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1323),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1462),
.B(n_1368),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1467),
.Y(n_1491)
);

AO31x2_ASAP7_75t_L g1492 ( 
.A1(n_1432),
.A2(n_1350),
.A3(n_1428),
.B(n_1324),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_SL g1493 ( 
.A(n_1465),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1323),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1323),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1468),
.B(n_1336),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1319),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1364),
.B(n_1376),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1461),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1350),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1468),
.B(n_1356),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1326),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1421),
.A2(n_1414),
.B(n_1409),
.Y(n_1503)
);

INVxp67_ASAP7_75t_SL g1504 ( 
.A(n_1333),
.Y(n_1504)
);

AO21x2_ASAP7_75t_L g1505 ( 
.A1(n_1432),
.A2(n_1428),
.B(n_1321),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1388),
.B(n_1343),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1421),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1446),
.B(n_1451),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1347),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1413),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1441),
.B(n_1320),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1408),
.A2(n_1320),
.B(n_1446),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1441),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1451),
.B(n_1460),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1460),
.B(n_1363),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1441),
.B(n_1379),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1407),
.B(n_1399),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1338),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1318),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1375),
.B(n_1348),
.Y(n_1520)
);

OA21x2_ASAP7_75t_L g1521 ( 
.A1(n_1430),
.A2(n_1466),
.B(n_1447),
.Y(n_1521)
);

OR2x6_ASAP7_75t_L g1522 ( 
.A(n_1330),
.B(n_1400),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1328),
.Y(n_1523)
);

OAI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1435),
.A2(n_1393),
.B1(n_1343),
.B2(n_1357),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1331),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1459),
.B(n_1386),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1332),
.Y(n_1527)
);

BUFx12f_ASAP7_75t_L g1528 ( 
.A(n_1322),
.Y(n_1528)
);

AO21x2_ASAP7_75t_L g1529 ( 
.A1(n_1424),
.A2(n_1472),
.B(n_1471),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1337),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1339),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1370),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1375),
.B(n_1327),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1340),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1342),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1327),
.B(n_1325),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1345),
.Y(n_1537)
);

CKINVDCx20_ASAP7_75t_R g1538 ( 
.A(n_1429),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1387),
.B(n_1406),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1391),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1433),
.Y(n_1541)
);

AO21x2_ASAP7_75t_L g1542 ( 
.A1(n_1437),
.A2(n_1470),
.B(n_1469),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1370),
.Y(n_1543)
);

BUFx6f_ASAP7_75t_L g1544 ( 
.A(n_1370),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1438),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1440),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1344),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1442),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1455),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1370),
.Y(n_1550)
);

INVx3_ASAP7_75t_L g1551 ( 
.A(n_1389),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1456),
.Y(n_1552)
);

INVx2_ASAP7_75t_SL g1553 ( 
.A(n_1394),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1397),
.A2(n_1401),
.B(n_1445),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1464),
.Y(n_1555)
);

OA21x2_ASAP7_75t_L g1556 ( 
.A1(n_1457),
.A2(n_1351),
.B(n_1362),
.Y(n_1556)
);

BUFx10_ASAP7_75t_L g1557 ( 
.A(n_1394),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1406),
.B(n_1384),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1389),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1365),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1420),
.Y(n_1561)
);

INVx2_ASAP7_75t_SL g1562 ( 
.A(n_1394),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1392),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1418),
.A2(n_1427),
.B(n_1426),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1396),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1381),
.B(n_1411),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1402),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1410),
.Y(n_1568)
);

AO21x2_ASAP7_75t_L g1569 ( 
.A1(n_1423),
.A2(n_1416),
.B(n_1422),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1407),
.B(n_1389),
.Y(n_1570)
);

CKINVDCx8_ASAP7_75t_R g1571 ( 
.A(n_1322),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1429),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1395),
.B(n_1407),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1398),
.B(n_1405),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1389),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1369),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1389),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1341),
.B(n_1452),
.Y(n_1578)
);

INVx2_ASAP7_75t_SL g1579 ( 
.A(n_1412),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1334),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1334),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1335),
.B(n_1453),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1341),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1453),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1453),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1463),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1359),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1374),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1374),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1431),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1390),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1450),
.B(n_1372),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1450),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1481),
.A2(n_1458),
.B(n_1372),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1511),
.B(n_1452),
.Y(n_1595)
);

INVxp67_ASAP7_75t_L g1596 ( 
.A(n_1502),
.Y(n_1596)
);

NOR2x1_ASAP7_75t_L g1597 ( 
.A(n_1529),
.B(n_1403),
.Y(n_1597)
);

NOR2x1_ASAP7_75t_SL g1598 ( 
.A(n_1488),
.B(n_1361),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1507),
.B(n_1359),
.Y(n_1599)
);

INVx4_ASAP7_75t_L g1600 ( 
.A(n_1488),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1484),
.B(n_1380),
.Y(n_1601)
);

AOI21xp33_ASAP7_75t_L g1602 ( 
.A1(n_1524),
.A2(n_1380),
.B(n_1361),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1484),
.B(n_1382),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1476),
.B(n_1382),
.Y(n_1604)
);

INVxp67_ASAP7_75t_L g1605 ( 
.A(n_1497),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1474),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1511),
.B(n_1357),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1507),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1542),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1516),
.B(n_1436),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1516),
.B(n_1436),
.Y(n_1611)
);

AOI221xp5_ASAP7_75t_L g1612 ( 
.A1(n_1498),
.A2(n_1415),
.B1(n_1403),
.B2(n_1367),
.C(n_1404),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1479),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1485),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1490),
.A2(n_1443),
.B(n_1431),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1507),
.B(n_1367),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1508),
.B(n_1425),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1542),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1482),
.B(n_1355),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1507),
.B(n_1404),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1508),
.B(n_1425),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1533),
.B(n_1434),
.Y(n_1622)
);

NOR2x1_ASAP7_75t_L g1623 ( 
.A(n_1529),
.B(n_1434),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1489),
.B(n_1355),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1521),
.A2(n_1315),
.B1(n_1449),
.B2(n_1346),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1514),
.B(n_1425),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1542),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1479),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1514),
.B(n_1477),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1520),
.B(n_1417),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1489),
.B(n_1355),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1509),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1475),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1512),
.B(n_1412),
.Y(n_1634)
);

NOR3xp33_ASAP7_75t_L g1635 ( 
.A(n_1480),
.B(n_1315),
.C(n_1449),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1473),
.B(n_1483),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1512),
.B(n_1412),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1512),
.B(n_1443),
.Y(n_1638)
);

INVx2_ASAP7_75t_SL g1639 ( 
.A(n_1523),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1499),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1494),
.B(n_1358),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1513),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1494),
.B(n_1358),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1512),
.B(n_1443),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1566),
.B(n_1346),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1566),
.B(n_1349),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1495),
.B(n_1360),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1519),
.B(n_1349),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1491),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1525),
.B(n_1360),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1525),
.B(n_1527),
.Y(n_1651)
);

BUFx2_ASAP7_75t_L g1652 ( 
.A(n_1485),
.Y(n_1652)
);

INVxp67_ASAP7_75t_SL g1653 ( 
.A(n_1504),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1521),
.A2(n_1517),
.B1(n_1515),
.B2(n_1501),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1491),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1496),
.A2(n_1561),
.B1(n_1526),
.B2(n_1515),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1506),
.B(n_1501),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1495),
.B(n_1523),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1530),
.B(n_1531),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1496),
.B(n_1547),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1549),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1561),
.A2(n_1493),
.B1(n_1522),
.B2(n_1573),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1530),
.B(n_1531),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1536),
.B(n_1503),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1634),
.B(n_1637),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1629),
.B(n_1603),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1634),
.B(n_1536),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1660),
.B(n_1549),
.Y(n_1668)
);

AOI221x1_ASAP7_75t_L g1669 ( 
.A1(n_1635),
.A2(n_1486),
.B1(n_1487),
.B2(n_1574),
.C(n_1500),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1610),
.B(n_1587),
.Y(n_1670)
);

OAI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1625),
.A2(n_1561),
.B1(n_1522),
.B2(n_1573),
.Y(n_1671)
);

NAND4xp25_ASAP7_75t_L g1672 ( 
.A(n_1636),
.B(n_1540),
.C(n_1518),
.D(n_1500),
.Y(n_1672)
);

NOR3xp33_ASAP7_75t_L g1673 ( 
.A(n_1602),
.B(n_1590),
.C(n_1578),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1637),
.B(n_1486),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1640),
.B(n_1534),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1640),
.B(n_1657),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1596),
.B(n_1535),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_SL g1678 ( 
.A1(n_1656),
.A2(n_1521),
.B1(n_1505),
.B2(n_1522),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1605),
.B(n_1535),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1610),
.B(n_1590),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1632),
.Y(n_1681)
);

AOI211xp5_ASAP7_75t_L g1682 ( 
.A1(n_1656),
.A2(n_1487),
.B(n_1583),
.C(n_1539),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1629),
.B(n_1517),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1653),
.B(n_1537),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1603),
.B(n_1517),
.Y(n_1685)
);

AOI221xp5_ASAP7_75t_L g1686 ( 
.A1(n_1654),
.A2(n_1539),
.B1(n_1558),
.B2(n_1505),
.C(n_1546),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1638),
.B(n_1644),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1662),
.A2(n_1521),
.B1(n_1505),
.B2(n_1522),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1616),
.B(n_1517),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1606),
.B(n_1541),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1604),
.A2(n_1522),
.B1(n_1558),
.B2(n_1556),
.Y(n_1691)
);

OA211x2_ASAP7_75t_L g1692 ( 
.A1(n_1612),
.A2(n_1492),
.B(n_1488),
.C(n_1544),
.Y(n_1692)
);

OAI21xp5_ASAP7_75t_SL g1693 ( 
.A1(n_1615),
.A2(n_1590),
.B(n_1570),
.Y(n_1693)
);

OAI21xp33_ASAP7_75t_L g1694 ( 
.A1(n_1623),
.A2(n_1554),
.B(n_1552),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1594),
.A2(n_1590),
.B1(n_1488),
.B2(n_1571),
.Y(n_1695)
);

NOR3xp33_ASAP7_75t_L g1696 ( 
.A(n_1611),
.B(n_1564),
.C(n_1575),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1645),
.A2(n_1556),
.B1(n_1554),
.B2(n_1528),
.Y(n_1697)
);

NAND4xp25_ASAP7_75t_L g1698 ( 
.A(n_1594),
.B(n_1545),
.C(n_1548),
.D(n_1546),
.Y(n_1698)
);

AOI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1638),
.A2(n_1644),
.B1(n_1650),
.B2(n_1648),
.C(n_1621),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1619),
.A2(n_1488),
.B1(n_1571),
.B2(n_1544),
.Y(n_1700)
);

NAND3xp33_ASAP7_75t_SL g1701 ( 
.A(n_1611),
.B(n_1607),
.C(n_1538),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1651),
.B(n_1529),
.Y(n_1702)
);

OAI21xp5_ASAP7_75t_SL g1703 ( 
.A1(n_1623),
.A2(n_1570),
.B(n_1577),
.Y(n_1703)
);

OAI21xp33_ASAP7_75t_L g1704 ( 
.A1(n_1597),
.A2(n_1545),
.B(n_1541),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1664),
.B(n_1510),
.Y(n_1705)
);

OAI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1619),
.A2(n_1544),
.B1(n_1577),
.B2(n_1575),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1597),
.A2(n_1544),
.B(n_1570),
.Y(n_1707)
);

OAI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1641),
.A2(n_1544),
.B1(n_1510),
.B2(n_1551),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_SL g1709 ( 
.A1(n_1650),
.A2(n_1544),
.B1(n_1570),
.B2(n_1532),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1641),
.A2(n_1559),
.B1(n_1532),
.B2(n_1550),
.Y(n_1710)
);

NAND4xp25_ASAP7_75t_L g1711 ( 
.A(n_1607),
.B(n_1548),
.C(n_1552),
.D(n_1555),
.Y(n_1711)
);

OAI221xp5_ASAP7_75t_SL g1712 ( 
.A1(n_1595),
.A2(n_1492),
.B1(n_1555),
.B2(n_1560),
.C(n_1581),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1643),
.A2(n_1551),
.B1(n_1532),
.B2(n_1543),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1632),
.Y(n_1714)
);

NAND3xp33_ASAP7_75t_L g1715 ( 
.A(n_1643),
.B(n_1585),
.C(n_1581),
.Y(n_1715)
);

NAND3xp33_ASAP7_75t_L g1716 ( 
.A(n_1647),
.B(n_1585),
.C(n_1556),
.Y(n_1716)
);

OAI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1647),
.A2(n_1550),
.B1(n_1551),
.B2(n_1532),
.Y(n_1717)
);

AOI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1648),
.A2(n_1560),
.B1(n_1563),
.B2(n_1565),
.C(n_1567),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1651),
.B(n_1478),
.Y(n_1719)
);

OAI221xp5_ASAP7_75t_SL g1720 ( 
.A1(n_1645),
.A2(n_1631),
.B1(n_1624),
.B2(n_1646),
.C(n_1630),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_SL g1721 ( 
.A1(n_1616),
.A2(n_1598),
.B1(n_1646),
.B2(n_1622),
.Y(n_1721)
);

NAND3xp33_ASAP7_75t_L g1722 ( 
.A(n_1609),
.B(n_1556),
.C(n_1584),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1620),
.B(n_1582),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1613),
.B(n_1492),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_SL g1725 ( 
.A1(n_1622),
.A2(n_1551),
.B(n_1550),
.Y(n_1725)
);

NAND4xp25_ASAP7_75t_L g1726 ( 
.A(n_1624),
.B(n_1563),
.C(n_1565),
.D(n_1567),
.Y(n_1726)
);

NOR3xp33_ASAP7_75t_L g1727 ( 
.A(n_1631),
.B(n_1564),
.C(n_1588),
.Y(n_1727)
);

NAND3xp33_ASAP7_75t_L g1728 ( 
.A(n_1609),
.B(n_1584),
.C(n_1586),
.Y(n_1728)
);

NAND3xp33_ASAP7_75t_L g1729 ( 
.A(n_1618),
.B(n_1586),
.C(n_1576),
.Y(n_1729)
);

AND2x2_ASAP7_75t_SL g1730 ( 
.A(n_1614),
.B(n_1475),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1628),
.B(n_1649),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1620),
.B(n_1580),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1655),
.B(n_1492),
.Y(n_1733)
);

OAI21xp33_ASAP7_75t_L g1734 ( 
.A1(n_1618),
.A2(n_1627),
.B(n_1621),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1659),
.B(n_1478),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1622),
.A2(n_1528),
.B1(n_1569),
.B2(n_1568),
.Y(n_1736)
);

NOR3xp33_ASAP7_75t_L g1737 ( 
.A(n_1600),
.B(n_1588),
.C(n_1589),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1674),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1674),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1681),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1714),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1702),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1668),
.B(n_1661),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1702),
.Y(n_1744)
);

AND2x4_ASAP7_75t_SL g1745 ( 
.A(n_1705),
.B(n_1600),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1690),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1719),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1684),
.Y(n_1748)
);

AND2x4_ASAP7_75t_SL g1749 ( 
.A(n_1705),
.B(n_1600),
.Y(n_1749)
);

OR2x2_ASAP7_75t_L g1750 ( 
.A(n_1687),
.B(n_1724),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1677),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1731),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1733),
.B(n_1719),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1665),
.B(n_1687),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1730),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_SL g1756 ( 
.A(n_1695),
.B(n_1620),
.Y(n_1756)
);

INVx2_ASAP7_75t_SL g1757 ( 
.A(n_1705),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1735),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1665),
.B(n_1664),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1679),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1667),
.B(n_1664),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1675),
.Y(n_1762)
);

INVx4_ASAP7_75t_L g1763 ( 
.A(n_1730),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1728),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1667),
.B(n_1666),
.Y(n_1765)
);

INVx5_ASAP7_75t_L g1766 ( 
.A(n_1689),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1683),
.B(n_1664),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1732),
.B(n_1614),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1729),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1734),
.Y(n_1770)
);

INVxp67_ASAP7_75t_SL g1771 ( 
.A(n_1670),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1722),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1676),
.B(n_1639),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1715),
.Y(n_1774)
);

INVxp67_ASAP7_75t_SL g1775 ( 
.A(n_1716),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1704),
.B(n_1694),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1711),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1727),
.B(n_1608),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1712),
.B(n_1658),
.Y(n_1779)
);

NOR2xp67_ASAP7_75t_L g1780 ( 
.A(n_1698),
.B(n_1608),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1723),
.B(n_1652),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1685),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1670),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1699),
.B(n_1608),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1726),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1686),
.B(n_1663),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1680),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1723),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1703),
.B(n_1642),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1696),
.B(n_1663),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1736),
.B(n_1599),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1710),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1706),
.Y(n_1793)
);

OAI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1776),
.A2(n_1678),
.B(n_1669),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1740),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1777),
.B(n_1672),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1789),
.Y(n_1797)
);

NAND2x1_ASAP7_75t_L g1798 ( 
.A(n_1763),
.B(n_1778),
.Y(n_1798)
);

NOR2x1p5_ASAP7_75t_L g1799 ( 
.A(n_1763),
.B(n_1701),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1789),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1740),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1747),
.Y(n_1802)
);

INVxp67_ASAP7_75t_SL g1803 ( 
.A(n_1783),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1747),
.Y(n_1804)
);

AND2x4_ASAP7_75t_L g1805 ( 
.A(n_1766),
.B(n_1737),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1741),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1741),
.Y(n_1807)
);

AND2x4_ASAP7_75t_L g1808 ( 
.A(n_1766),
.B(n_1707),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1752),
.B(n_1751),
.Y(n_1809)
);

NAND5xp2_ASAP7_75t_L g1810 ( 
.A(n_1775),
.B(n_1688),
.C(n_1693),
.D(n_1682),
.E(n_1721),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1742),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1787),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1759),
.B(n_1725),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1750),
.B(n_1772),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1763),
.B(n_1673),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1759),
.B(n_1709),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1742),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1751),
.B(n_1718),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1759),
.B(n_1697),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1759),
.B(n_1697),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1747),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1758),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1766),
.B(n_1633),
.Y(n_1823)
);

NOR3xp33_ASAP7_75t_SL g1824 ( 
.A(n_1756),
.B(n_1572),
.C(n_1720),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1750),
.B(n_1691),
.Y(n_1825)
);

NOR2xp33_ASAP7_75t_L g1826 ( 
.A(n_1777),
.B(n_1622),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1744),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1744),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1754),
.B(n_1691),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1772),
.B(n_1736),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1758),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1754),
.B(n_1620),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1772),
.B(n_1713),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1738),
.Y(n_1834)
);

INVx2_ASAP7_75t_SL g1835 ( 
.A(n_1766),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1785),
.B(n_1617),
.Y(n_1836)
);

AOI32xp33_ASAP7_75t_L g1837 ( 
.A1(n_1776),
.A2(n_1671),
.A3(n_1688),
.B1(n_1626),
.B2(n_1617),
.Y(n_1837)
);

OAI21xp33_ASAP7_75t_L g1838 ( 
.A1(n_1775),
.A2(n_1785),
.B(n_1774),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1758),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1739),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1748),
.Y(n_1841)
);

BUFx2_ASAP7_75t_L g1842 ( 
.A(n_1763),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1760),
.B(n_1601),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1788),
.Y(n_1844)
);

AOI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1780),
.A2(n_1692),
.B1(n_1700),
.B2(n_1708),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1748),
.Y(n_1846)
);

OAI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1794),
.A2(n_1780),
.B1(n_1755),
.B2(n_1786),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1825),
.B(n_1786),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1813),
.B(n_1761),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1795),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1795),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1796),
.B(n_1770),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1801),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1801),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1838),
.B(n_1770),
.Y(n_1855)
);

NOR2x1_ASAP7_75t_L g1856 ( 
.A(n_1799),
.B(n_1769),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1806),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1812),
.B(n_1774),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1825),
.B(n_1779),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1806),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1807),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1830),
.B(n_1779),
.Y(n_1862)
);

NOR2x1_ASAP7_75t_L g1863 ( 
.A(n_1799),
.B(n_1769),
.Y(n_1863)
);

NOR2xp67_ASAP7_75t_L g1864 ( 
.A(n_1835),
.B(n_1766),
.Y(n_1864)
);

NAND4xp25_ASAP7_75t_SL g1865 ( 
.A(n_1837),
.B(n_1755),
.C(n_1784),
.D(n_1788),
.Y(n_1865)
);

AOI32xp33_ASAP7_75t_L g1866 ( 
.A1(n_1842),
.A2(n_1784),
.A3(n_1793),
.B1(n_1788),
.B2(n_1764),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1832),
.B(n_1767),
.Y(n_1867)
);

AND2x4_ASAP7_75t_L g1868 ( 
.A(n_1842),
.B(n_1778),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1813),
.B(n_1761),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1818),
.B(n_1771),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1830),
.B(n_1743),
.Y(n_1871)
);

AOI21xp33_ASAP7_75t_SL g1872 ( 
.A1(n_1815),
.A2(n_1764),
.B(n_1781),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1803),
.B(n_1790),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1836),
.B(n_1790),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1816),
.B(n_1757),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1807),
.Y(n_1876)
);

INVxp67_ASAP7_75t_L g1877 ( 
.A(n_1814),
.Y(n_1877)
);

NOR2xp33_ASAP7_75t_SL g1878 ( 
.A(n_1835),
.B(n_1600),
.Y(n_1878)
);

BUFx2_ASAP7_75t_L g1879 ( 
.A(n_1832),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1814),
.B(n_1743),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1805),
.B(n_1778),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1810),
.B(n_1760),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1797),
.B(n_1800),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1809),
.B(n_1829),
.Y(n_1884)
);

AND2x4_ASAP7_75t_SL g1885 ( 
.A(n_1824),
.B(n_1768),
.Y(n_1885)
);

INVx1_ASAP7_75t_SL g1886 ( 
.A(n_1833),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1841),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1829),
.B(n_1746),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1802),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1837),
.B(n_1766),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1841),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1846),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1816),
.B(n_1767),
.Y(n_1893)
);

INVx1_ASAP7_75t_SL g1894 ( 
.A(n_1833),
.Y(n_1894)
);

INVx2_ASAP7_75t_SL g1895 ( 
.A(n_1798),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1846),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1826),
.B(n_1746),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1802),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1819),
.B(n_1757),
.Y(n_1899)
);

INVxp67_ASAP7_75t_L g1900 ( 
.A(n_1797),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1850),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1889),
.Y(n_1902)
);

INVxp67_ASAP7_75t_SL g1903 ( 
.A(n_1856),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1871),
.B(n_1800),
.Y(n_1904)
);

INVx1_ASAP7_75t_SL g1905 ( 
.A(n_1886),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1882),
.B(n_1834),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1889),
.Y(n_1907)
);

NOR2x1_ASAP7_75t_L g1908 ( 
.A(n_1863),
.B(n_1798),
.Y(n_1908)
);

INVx1_ASAP7_75t_SL g1909 ( 
.A(n_1894),
.Y(n_1909)
);

CKINVDCx16_ASAP7_75t_R g1910 ( 
.A(n_1882),
.Y(n_1910)
);

INVx1_ASAP7_75t_SL g1911 ( 
.A(n_1895),
.Y(n_1911)
);

OR2x2_ASAP7_75t_L g1912 ( 
.A(n_1880),
.B(n_1844),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1870),
.B(n_1852),
.Y(n_1913)
);

HB1xp67_ASAP7_75t_L g1914 ( 
.A(n_1877),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1855),
.B(n_1819),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1866),
.B(n_1834),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1849),
.B(n_1820),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1851),
.Y(n_1918)
);

INVx1_ASAP7_75t_SL g1919 ( 
.A(n_1895),
.Y(n_1919)
);

AOI22xp33_ASAP7_75t_L g1920 ( 
.A1(n_1865),
.A2(n_1820),
.B1(n_1808),
.B2(n_1805),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1862),
.B(n_1859),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1858),
.B(n_1840),
.Y(n_1922)
);

AOI22x1_ASAP7_75t_L g1923 ( 
.A1(n_1848),
.A2(n_1805),
.B1(n_1808),
.B2(n_1823),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1888),
.B(n_1844),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1849),
.B(n_1869),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1898),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1869),
.B(n_1808),
.Y(n_1927)
);

INVx5_ASAP7_75t_L g1928 ( 
.A(n_1868),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1872),
.B(n_1840),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1853),
.Y(n_1930)
);

CKINVDCx16_ASAP7_75t_R g1931 ( 
.A(n_1847),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1877),
.B(n_1792),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1900),
.Y(n_1933)
);

BUFx3_ASAP7_75t_L g1934 ( 
.A(n_1868),
.Y(n_1934)
);

BUFx6f_ASAP7_75t_L g1935 ( 
.A(n_1868),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1884),
.B(n_1811),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1893),
.B(n_1808),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1874),
.B(n_1782),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1898),
.Y(n_1939)
);

AOI22x1_ASAP7_75t_L g1940 ( 
.A1(n_1875),
.A2(n_1879),
.B1(n_1900),
.B2(n_1890),
.Y(n_1940)
);

AOI221x1_ASAP7_75t_L g1941 ( 
.A1(n_1906),
.A2(n_1873),
.B1(n_1887),
.B2(n_1896),
.C(n_1892),
.Y(n_1941)
);

O2A1O1Ixp5_ASAP7_75t_L g1942 ( 
.A1(n_1903),
.A2(n_1890),
.B(n_1883),
.C(n_1881),
.Y(n_1942)
);

AOI221xp5_ASAP7_75t_L g1943 ( 
.A1(n_1931),
.A2(n_1881),
.B1(n_1885),
.B2(n_1891),
.C(n_1897),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1933),
.Y(n_1944)
);

AOI21xp33_ASAP7_75t_L g1945 ( 
.A1(n_1940),
.A2(n_1881),
.B(n_1878),
.Y(n_1945)
);

A2O1A1Ixp33_ASAP7_75t_L g1946 ( 
.A1(n_1908),
.A2(n_1885),
.B(n_1845),
.C(n_1864),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1914),
.Y(n_1947)
);

OAI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1931),
.A2(n_1875),
.B1(n_1766),
.B2(n_1899),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1910),
.B(n_1899),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1910),
.B(n_1867),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1901),
.Y(n_1951)
);

OAI222xp33_ASAP7_75t_L g1952 ( 
.A1(n_1940),
.A2(n_1781),
.B1(n_1792),
.B2(n_1791),
.C1(n_1782),
.C2(n_1854),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1925),
.B(n_1857),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1905),
.B(n_1860),
.Y(n_1954)
);

OAI31xp33_ASAP7_75t_L g1955 ( 
.A1(n_1916),
.A2(n_1823),
.A3(n_1861),
.B(n_1876),
.Y(n_1955)
);

NOR2xp33_ASAP7_75t_L g1956 ( 
.A(n_1913),
.B(n_1843),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1901),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1935),
.Y(n_1958)
);

AOI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1915),
.A2(n_1792),
.B1(n_1823),
.B2(n_1791),
.Y(n_1959)
);

OAI22xp5_ASAP7_75t_L g1960 ( 
.A1(n_1920),
.A2(n_1753),
.B1(n_1823),
.B2(n_1745),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1918),
.Y(n_1961)
);

OA21x2_ASAP7_75t_L g1962 ( 
.A1(n_1929),
.A2(n_1821),
.B(n_1804),
.Y(n_1962)
);

OR2x2_ASAP7_75t_L g1963 ( 
.A(n_1905),
.B(n_1811),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1935),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1909),
.B(n_1762),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1918),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1909),
.B(n_1762),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1925),
.B(n_1765),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1930),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1947),
.B(n_1917),
.Y(n_1970)
);

INVxp67_ASAP7_75t_L g1971 ( 
.A(n_1947),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1949),
.B(n_1917),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1943),
.A2(n_1908),
.B1(n_1921),
.B2(n_1923),
.Y(n_1973)
);

INVx1_ASAP7_75t_SL g1974 ( 
.A(n_1950),
.Y(n_1974)
);

NAND2x1p5_ASAP7_75t_L g1975 ( 
.A(n_1958),
.B(n_1928),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1969),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1944),
.B(n_1921),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1958),
.B(n_1934),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1969),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1963),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1946),
.B(n_1928),
.Y(n_1981)
);

INVxp67_ASAP7_75t_L g1982 ( 
.A(n_1964),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1964),
.B(n_1934),
.Y(n_1983)
);

NAND2x1_ASAP7_75t_L g1984 ( 
.A(n_1948),
.B(n_1935),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1963),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1954),
.B(n_1934),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1951),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1957),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1961),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1966),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1953),
.Y(n_1991)
);

AOI22xp33_ASAP7_75t_L g1992 ( 
.A1(n_1960),
.A2(n_1923),
.B1(n_1935),
.B2(n_1904),
.Y(n_1992)
);

OAI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1981),
.A2(n_1942),
.B(n_1941),
.Y(n_1993)
);

OAI21xp33_ASAP7_75t_L g1994 ( 
.A1(n_1973),
.A2(n_1977),
.B(n_1992),
.Y(n_1994)
);

O2A1O1Ixp33_ASAP7_75t_L g1995 ( 
.A1(n_1971),
.A2(n_1952),
.B(n_1946),
.C(n_1945),
.Y(n_1995)
);

OAI22xp33_ASAP7_75t_L g1996 ( 
.A1(n_1984),
.A2(n_1941),
.B1(n_1928),
.B2(n_1935),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1974),
.B(n_1953),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1978),
.B(n_1968),
.Y(n_1998)
);

NAND2xp33_ASAP7_75t_SL g1999 ( 
.A(n_1970),
.B(n_1935),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1978),
.B(n_1968),
.Y(n_2000)
);

OAI22xp5_ASAP7_75t_L g2001 ( 
.A1(n_1972),
.A2(n_1928),
.B1(n_1959),
.B2(n_1956),
.Y(n_2001)
);

NAND4xp25_ASAP7_75t_L g2002 ( 
.A(n_1986),
.B(n_1955),
.C(n_1911),
.D(n_1919),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_SL g2003 ( 
.A(n_1975),
.B(n_1928),
.Y(n_2003)
);

OAI211xp5_ASAP7_75t_SL g2004 ( 
.A1(n_1971),
.A2(n_1919),
.B(n_1911),
.C(n_1967),
.Y(n_2004)
);

OAI21xp5_ASAP7_75t_L g2005 ( 
.A1(n_1975),
.A2(n_1965),
.B(n_1928),
.Y(n_2005)
);

OAI211xp5_ASAP7_75t_SL g2006 ( 
.A1(n_1983),
.A2(n_1980),
.B(n_1985),
.C(n_1982),
.Y(n_2006)
);

OAI221xp5_ASAP7_75t_SL g2007 ( 
.A1(n_1991),
.A2(n_1982),
.B1(n_1989),
.B2(n_1988),
.C(n_1987),
.Y(n_2007)
);

NAND3xp33_ASAP7_75t_L g2008 ( 
.A(n_1990),
.B(n_1962),
.C(n_1904),
.Y(n_2008)
);

NAND3xp33_ASAP7_75t_L g2009 ( 
.A(n_1993),
.B(n_1979),
.C(n_1976),
.Y(n_2009)
);

AOI211xp5_ASAP7_75t_L g2010 ( 
.A1(n_1995),
.A2(n_1932),
.B(n_1922),
.C(n_1930),
.Y(n_2010)
);

NAND4xp75_ASAP7_75t_L g2011 ( 
.A(n_2003),
.B(n_1962),
.C(n_1927),
.D(n_1907),
.Y(n_2011)
);

AOI211x1_ASAP7_75t_L g2012 ( 
.A1(n_1994),
.A2(n_1996),
.B(n_2005),
.C(n_2002),
.Y(n_2012)
);

NOR3x1_ASAP7_75t_L g2013 ( 
.A(n_1997),
.B(n_2000),
.C(n_1998),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_SL g2014 ( 
.A(n_1999),
.B(n_1924),
.Y(n_2014)
);

NOR3xp33_ASAP7_75t_L g2015 ( 
.A(n_2006),
.B(n_1936),
.C(n_1907),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_2008),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_2001),
.B(n_1938),
.Y(n_2017)
);

NOR2xp67_ASAP7_75t_L g2018 ( 
.A(n_2004),
.B(n_1902),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_L g2019 ( 
.A(n_2007),
.B(n_1936),
.Y(n_2019)
);

OAI211xp5_ASAP7_75t_SL g2020 ( 
.A1(n_1994),
.A2(n_1939),
.B(n_1902),
.C(n_1907),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_2018),
.B(n_1924),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_SL g2022 ( 
.A(n_2016),
.B(n_1937),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_2012),
.B(n_1937),
.Y(n_2023)
);

OAI211xp5_ASAP7_75t_L g2024 ( 
.A1(n_2019),
.A2(n_1962),
.B(n_1926),
.C(n_1902),
.Y(n_2024)
);

OAI21xp5_ASAP7_75t_L g2025 ( 
.A1(n_2009),
.A2(n_1927),
.B(n_1926),
.Y(n_2025)
);

NOR4xp25_ASAP7_75t_L g2026 ( 
.A(n_2020),
.B(n_1939),
.C(n_1926),
.D(n_1912),
.Y(n_2026)
);

NAND3xp33_ASAP7_75t_L g2027 ( 
.A(n_2015),
.B(n_1939),
.C(n_1912),
.Y(n_2027)
);

NOR2xp33_ASAP7_75t_L g2028 ( 
.A(n_2017),
.B(n_1804),
.Y(n_2028)
);

NOR4xp25_ASAP7_75t_L g2029 ( 
.A(n_2014),
.B(n_1817),
.C(n_1827),
.D(n_1828),
.Y(n_2029)
);

AO22x2_ASAP7_75t_L g2030 ( 
.A1(n_2023),
.A2(n_2011),
.B1(n_2013),
.B2(n_2010),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_2022),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_2021),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_2027),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2028),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_2025),
.Y(n_2035)
);

NOR2x1_ASAP7_75t_L g2036 ( 
.A(n_2024),
.B(n_1817),
.Y(n_2036)
);

AOI22xp5_ASAP7_75t_L g2037 ( 
.A1(n_2026),
.A2(n_1778),
.B1(n_1745),
.B2(n_1749),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2029),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_2031),
.B(n_1827),
.Y(n_2039)
);

OAI21xp5_ASAP7_75t_L g2040 ( 
.A1(n_2033),
.A2(n_1773),
.B(n_1828),
.Y(n_2040)
);

NOR3xp33_ASAP7_75t_L g2041 ( 
.A(n_2035),
.B(n_1773),
.C(n_1717),
.Y(n_2041)
);

OR2x2_ASAP7_75t_L g2042 ( 
.A(n_2032),
.B(n_2034),
.Y(n_2042)
);

AOI22xp33_ASAP7_75t_SL g2043 ( 
.A1(n_2030),
.A2(n_1598),
.B1(n_1749),
.B2(n_1745),
.Y(n_2043)
);

NAND2x1_ASAP7_75t_L g2044 ( 
.A(n_2036),
.B(n_1821),
.Y(n_2044)
);

NAND2x1p5_ASAP7_75t_L g2045 ( 
.A(n_2042),
.B(n_2038),
.Y(n_2045)
);

XNOR2xp5_ASAP7_75t_L g2046 ( 
.A(n_2039),
.B(n_2030),
.Y(n_2046)
);

NOR2x1_ASAP7_75t_L g2047 ( 
.A(n_2044),
.B(n_2037),
.Y(n_2047)
);

AND3x2_ASAP7_75t_L g2048 ( 
.A(n_2041),
.B(n_1592),
.C(n_1831),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_2048),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_2045),
.Y(n_2050)
);

NAND4xp25_ASAP7_75t_SL g2051 ( 
.A(n_2050),
.B(n_2047),
.C(n_2043),
.D(n_2040),
.Y(n_2051)
);

OAI221xp5_ASAP7_75t_L g2052 ( 
.A1(n_2051),
.A2(n_2046),
.B1(n_2049),
.B2(n_1822),
.C(n_1831),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2051),
.Y(n_2053)
);

AOI21xp33_ASAP7_75t_L g2054 ( 
.A1(n_2053),
.A2(n_2049),
.B(n_1562),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_2052),
.B(n_1822),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_2055),
.B(n_1839),
.Y(n_2056)
);

AOI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_2056),
.A2(n_2054),
.B1(n_1839),
.B2(n_1753),
.Y(n_2057)
);

NAND5xp2_ASAP7_75t_L g2058 ( 
.A(n_2057),
.B(n_1593),
.C(n_1626),
.D(n_1589),
.E(n_1591),
.Y(n_2058)
);

OAI221xp5_ASAP7_75t_R g2059 ( 
.A1(n_2058),
.A2(n_1749),
.B1(n_1557),
.B2(n_1579),
.C(n_1562),
.Y(n_2059)
);

AOI211xp5_ASAP7_75t_L g2060 ( 
.A1(n_2059),
.A2(n_1579),
.B(n_1553),
.C(n_1717),
.Y(n_2060)
);


endmodule