module fake_jpeg_12323_n_236 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_9),
.B(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_3),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_39),
.B(n_62),
.Y(n_90)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_66),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_13),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_44),
.B(n_57),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_45),
.Y(n_83)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_27),
.Y(n_49)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_11),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_24),
.B(n_1),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_32),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_102),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_24),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_71),
.B(n_79),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_38),
.B1(n_30),
.B2(n_17),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g114 ( 
.A1(n_72),
.A2(n_77),
.B1(n_99),
.B2(n_5),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_20),
.B1(n_31),
.B2(n_25),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_75),
.A2(n_81),
.B1(n_94),
.B2(n_101),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_38),
.B1(n_30),
.B2(n_17),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_65),
.A2(n_41),
.B1(n_43),
.B2(n_31),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_SL g82 ( 
.A(n_49),
.Y(n_82)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_25),
.B1(n_20),
.B2(n_29),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_32),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_97),
.B(n_98),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_29),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_48),
.A2(n_37),
.B1(n_15),
.B2(n_26),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_56),
.A2(n_37),
.B1(n_26),
.B2(n_3),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_1),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_2),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_4),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_106),
.B(n_121),
.Y(n_146)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_107),
.Y(n_154)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_4),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_111),
.B(n_116),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_122),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_5),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_5),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_118),
.B(n_120),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_7),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_124),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_8),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_77),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_96),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_123),
.B(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_103),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_130),
.Y(n_151)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_128),
.A2(n_134),
.B1(n_137),
.B2(n_107),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_70),
.B(n_72),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_132),
.Y(n_156)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_85),
.A2(n_87),
.B(n_100),
.C(n_69),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_112),
.B(n_133),
.C(n_132),
.Y(n_163)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_92),
.C(n_100),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_143),
.C(n_144),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_69),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_91),
.B1(n_92),
.B2(n_105),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_144),
.A2(n_126),
.B1(n_136),
.B2(n_137),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_91),
.B1(n_87),
.B2(n_89),
.Y(n_147)
);

AO21x1_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_163),
.B(n_145),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_95),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_153),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_135),
.A2(n_95),
.B1(n_114),
.B2(n_106),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_149),
.A2(n_162),
.B1(n_133),
.B2(n_145),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_95),
.Y(n_153)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

A2O1A1O1Ixp25_ASAP7_75t_L g159 ( 
.A1(n_108),
.A2(n_129),
.B(n_109),
.C(n_115),
.D(n_117),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_159),
.B(n_153),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_129),
.A2(n_131),
.B1(n_124),
.B2(n_128),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_127),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_179),
.C(n_139),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_134),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_167),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_122),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_172),
.Y(n_189)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_171),
.B(n_173),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_138),
.B(n_150),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_162),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_175),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_156),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_160),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_177),
.Y(n_195)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_152),
.B(n_146),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_182),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_155),
.C(n_163),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_183),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_141),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_149),
.A2(n_148),
.B1(n_140),
.B2(n_141),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_196),
.C(n_182),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_191),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_161),
.B(n_154),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_199),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_157),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_168),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_193),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_161),
.C(n_154),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_177),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

OAI32xp33_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_171),
.A3(n_175),
.B1(n_166),
.B2(n_183),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_185),
.A2(n_181),
.B1(n_165),
.B2(n_179),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_202),
.A2(n_190),
.B1(n_187),
.B2(n_184),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_189),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_209),
.Y(n_212)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_206),
.C(n_208),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_196),
.C(n_194),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_170),
.C(n_165),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_200),
.Y(n_213)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_198),
.C(n_195),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_216),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_198),
.B(n_189),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_215),
.A2(n_208),
.B(n_207),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_195),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_218),
.A2(n_209),
.B1(n_201),
.B2(n_199),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_222),
.Y(n_227)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_221),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_214),
.A2(n_210),
.B(n_207),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_212),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_226),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_212),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_223),
.C(n_211),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_230),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_223),
.C(n_211),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_216),
.Y(n_233)
);

AOI21x1_ASAP7_75t_L g234 ( 
.A1(n_233),
.A2(n_215),
.B(n_228),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_232),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_167),
.Y(n_236)
);


endmodule