module fake_jpeg_1101_n_130 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_26),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_48),
.Y(n_58)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_54),
.Y(n_60)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_40),
.Y(n_68)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_59),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_53),
.A2(n_37),
.B1(n_35),
.B2(n_42),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_63),
.B(n_66),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_55),
.B1(n_35),
.B2(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_38),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_38),
.B(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_46),
.C(n_40),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_0),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_47),
.B1(n_44),
.B2(n_43),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_66),
.Y(n_80)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_45),
.Y(n_87)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_77),
.B(n_0),
.Y(n_86)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_79),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_81),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_65),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_79),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_93),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_1),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_87),
.B(n_4),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_76),
.A2(n_59),
.B(n_36),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_88),
.A2(n_89),
.B(n_73),
.Y(n_96)
);

AO21x1_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_59),
.B(n_16),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_73),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_18),
.Y(n_93)
);

NOR4xp25_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_22),
.C(n_33),
.D(n_32),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_101),
.C(n_107),
.Y(n_110)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_102),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_104),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_72),
.B(n_2),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_1),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_105),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_2),
.B(n_3),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_3),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_15),
.C(n_30),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_91),
.C(n_84),
.Y(n_111)
);

AOI21x1_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_31),
.B(n_29),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_108),
.B(n_7),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_112),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_SL g112 ( 
.A(n_100),
.B(n_28),
.C(n_27),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_25),
.B(n_24),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_115),
.Y(n_122)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_101),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_120),
.B1(n_114),
.B2(n_110),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_109),
.A2(n_107),
.B1(n_106),
.B2(n_9),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_113),
.C(n_116),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_123),
.B(n_124),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_122),
.C(n_120),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_112),
.A3(n_110),
.B1(n_118),
.B2(n_23),
.C1(n_12),
.C2(n_7),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

OAI321xp33_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_8),
.A3(n_9),
.B1(n_11),
.B2(n_13),
.C(n_14),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_8),
.Y(n_130)
);


endmodule