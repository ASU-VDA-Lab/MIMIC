module fake_jpeg_28987_n_447 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_447);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_447;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_10),
.Y(n_29)
);

INVxp33_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_23),
.B(n_9),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_48),
.B(n_51),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_9),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_54),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_23),
.B(n_7),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_85),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_25),
.B(n_7),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_25),
.B(n_10),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_59),
.Y(n_135)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_30),
.B(n_10),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_65),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_5),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_69),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_5),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_70),
.B(n_81),
.Y(n_136)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

BUFx4f_ASAP7_75t_SL g100 ( 
.A(n_77),
.Y(n_100)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_34),
.B(n_5),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_84),
.Y(n_121)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_33),
.B(n_11),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_89),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g112 ( 
.A(n_87),
.Y(n_112)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_88),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_91),
.Y(n_120)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_33),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_28),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_93),
.B(n_96),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_91),
.A2(n_39),
.B1(n_46),
.B2(n_43),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_95),
.A2(n_106),
.B1(n_108),
.B2(n_0),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_28),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_52),
.A2(n_68),
.B1(n_90),
.B2(n_55),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_103),
.A2(n_122),
.B1(n_142),
.B2(n_130),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_59),
.A2(n_39),
.B1(n_46),
.B2(n_43),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_32),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_107),
.B(n_130),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_84),
.A2(n_39),
.B1(n_46),
.B2(n_43),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_88),
.A2(n_22),
.B1(n_41),
.B2(n_37),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_143),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_62),
.B(n_34),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_128),
.B(n_133),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_57),
.B(n_22),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_63),
.A2(n_46),
.B1(n_41),
.B2(n_37),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_74),
.B(n_35),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_73),
.B(n_35),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_145),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_72),
.A2(n_32),
.B1(n_43),
.B2(n_45),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_SL g143 ( 
.A1(n_76),
.A2(n_44),
.B(n_45),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_79),
.B(n_33),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_92),
.A2(n_44),
.B(n_43),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_146),
.B(n_121),
.C(n_129),
.Y(n_198)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_147),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_144),
.A2(n_75),
.B1(n_77),
.B2(n_102),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_148),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_94),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_149),
.B(n_174),
.Y(n_216)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_150),
.Y(n_214)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_152),
.Y(n_217)
);

O2A1O1Ixp33_ASAP7_75t_SL g153 ( 
.A1(n_146),
.A2(n_87),
.B(n_83),
.C(n_80),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_153),
.A2(n_157),
.B1(n_159),
.B2(n_178),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_45),
.Y(n_154)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_154),
.B(n_158),
.CI(n_100),
.CON(n_224),
.SN(n_224)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_155),
.A2(n_168),
.B1(n_180),
.B2(n_188),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_107),
.A2(n_45),
.B1(n_47),
.B2(n_2),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_93),
.B(n_45),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_144),
.A2(n_47),
.B1(n_1),
.B2(n_2),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_161),
.Y(n_219)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_102),
.A2(n_11),
.B1(n_1),
.B2(n_3),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_164),
.Y(n_231)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

INVx8_ASAP7_75t_L g229 ( 
.A(n_165),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_110),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_167),
.B(n_172),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_98),
.A2(n_12),
.B1(n_3),
.B2(n_4),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_139),
.Y(n_169)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_116),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_94),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_98),
.A2(n_3),
.B1(n_4),
.B2(n_11),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_101),
.A2(n_3),
.B1(n_4),
.B2(n_13),
.Y(n_180)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

O2A1O1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_145),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_194),
.Y(n_200)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_105),
.Y(n_184)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_186),
.Y(n_225)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_126),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_187),
.A2(n_193),
.B1(n_196),
.B2(n_127),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_114),
.A2(n_13),
.B1(n_14),
.B2(n_0),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_189),
.Y(n_206)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_99),
.A2(n_0),
.B1(n_14),
.B2(n_122),
.Y(n_190)
);

AO22x2_ASAP7_75t_SL g230 ( 
.A1(n_190),
.A2(n_100),
.B1(n_105),
.B2(n_137),
.Y(n_230)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_140),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_191),
.Y(n_227)
);

AND2x4_ASAP7_75t_L g192 ( 
.A(n_96),
.B(n_0),
.Y(n_192)
);

AND2x2_ASAP7_75t_SL g241 ( 
.A(n_192),
.B(n_183),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_113),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_99),
.A2(n_0),
.B1(n_121),
.B2(n_101),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_L g195 ( 
.A1(n_114),
.A2(n_134),
.B1(n_111),
.B2(n_132),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_195),
.A2(n_134),
.B1(n_111),
.B2(n_135),
.Y(n_202)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_140),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_120),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_197),
.B(n_104),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_198),
.A2(n_109),
.B(n_97),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_136),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_199),
.B(n_203),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_202),
.A2(n_228),
.B1(n_240),
.B2(n_195),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_121),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_207),
.B(n_224),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_112),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_212),
.B(n_232),
.Y(n_257)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_151),
.B(n_100),
.C(n_112),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_158),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_179),
.A2(n_132),
.B1(n_135),
.B2(n_112),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_181),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_105),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_154),
.B(n_151),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_236),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_151),
.B(n_137),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_238),
.A2(n_156),
.B1(n_166),
.B2(n_193),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_170),
.A2(n_115),
.B(n_137),
.C(n_127),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_239),
.B(n_242),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_155),
.A2(n_104),
.B1(n_137),
.B2(n_194),
.Y(n_240)
);

XNOR2x1_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_232),
.Y(n_265)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_243),
.Y(n_285)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_201),
.Y(n_244)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_244),
.Y(n_288)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_247),
.Y(n_290)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_208),
.Y(n_248)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_248),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_225),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_249),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_230),
.A2(n_153),
.B1(n_190),
.B2(n_157),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_250),
.A2(n_254),
.B1(n_266),
.B2(n_267),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_163),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_251),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_210),
.B(n_189),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_252),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_233),
.A2(n_198),
.B1(n_159),
.B2(n_190),
.Y(n_254)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

INVx13_ASAP7_75t_L g316 ( 
.A(n_255),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_256),
.B(n_265),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_158),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_259),
.B(n_224),
.C(n_241),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_216),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_260),
.B(n_263),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_261),
.A2(n_269),
.B1(n_271),
.B2(n_233),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_262),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_207),
.B(n_152),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_200),
.B(n_190),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_264),
.Y(n_282)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_208),
.Y(n_268)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_268),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_230),
.A2(n_147),
.B1(n_150),
.B2(n_162),
.Y(n_269)
);

BUFx12_ASAP7_75t_L g270 ( 
.A(n_218),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_270),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_230),
.A2(n_177),
.B1(n_175),
.B2(n_191),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_212),
.A2(n_169),
.B(n_165),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_272),
.A2(n_217),
.B(n_221),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_199),
.B(n_182),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_L g306 ( 
.A1(n_273),
.A2(n_278),
.B(n_200),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_226),
.Y(n_274)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_274),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_213),
.A2(n_176),
.B(n_184),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_275),
.A2(n_271),
.B(n_269),
.Y(n_310)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_211),
.Y(n_276)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_211),
.Y(n_277)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_277),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_224),
.B(n_203),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_236),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_280),
.Y(n_293)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_220),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_205),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_227),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_283),
.A2(n_289),
.B1(n_310),
.B2(n_314),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_213),
.B1(n_231),
.B2(n_219),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_303),
.C(n_259),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_254),
.A2(n_267),
.B1(n_204),
.B2(n_246),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_294),
.A2(n_305),
.B1(n_215),
.B2(n_235),
.Y(n_338)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_296),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_245),
.B(n_241),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_299),
.B(n_309),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_253),
.B(n_239),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_279),
.A2(n_231),
.B1(n_219),
.B2(n_202),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_306),
.Y(n_319)
);

AND2x6_ASAP7_75t_L g307 ( 
.A(n_253),
.B(n_274),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_307),
.B(n_311),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_308),
.Y(n_327)
);

O2A1O1Ixp33_ASAP7_75t_L g309 ( 
.A1(n_275),
.A2(n_264),
.B(n_257),
.C(n_272),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_278),
.A2(n_258),
.B(n_257),
.Y(n_311)
);

O2A1O1Ixp33_ASAP7_75t_L g312 ( 
.A1(n_258),
.A2(n_206),
.B(n_221),
.C(n_227),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_312),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_261),
.A2(n_245),
.B1(n_265),
.B2(n_256),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_289),
.A2(n_249),
.B1(n_243),
.B2(n_247),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_317),
.A2(n_343),
.B1(n_345),
.B2(n_297),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_287),
.A2(n_260),
.B1(n_268),
.B2(n_248),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_318),
.A2(n_329),
.B1(n_330),
.B2(n_338),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_321),
.B(n_322),
.C(n_326),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_280),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_296),
.Y(n_323)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_323),
.Y(n_346)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_285),
.Y(n_324)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_324),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_295),
.B(n_277),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_295),
.B(n_292),
.C(n_303),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_328),
.B(n_333),
.C(n_334),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_287),
.A2(n_276),
.B1(n_244),
.B2(n_222),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_294),
.A2(n_255),
.B1(n_222),
.B2(n_262),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_285),
.Y(n_331)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_331),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_220),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_301),
.B(n_235),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_283),
.A2(n_206),
.B1(n_217),
.B2(n_229),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_335),
.A2(n_286),
.B(n_297),
.Y(n_362)
);

AO22x1_ASAP7_75t_L g336 ( 
.A1(n_309),
.A2(n_270),
.B1(n_281),
.B2(n_214),
.Y(n_336)
);

AO21x2_ASAP7_75t_L g351 ( 
.A1(n_336),
.A2(n_291),
.B(n_300),
.Y(n_351)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_290),
.Y(n_337)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_337),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_301),
.B(n_215),
.C(n_218),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_339),
.B(n_341),
.C(n_344),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_299),
.B(n_313),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_310),
.A2(n_282),
.B1(n_315),
.B2(n_312),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_293),
.B(n_270),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_282),
.A2(n_308),
.B1(n_305),
.B2(n_291),
.Y(n_345)
);

AO21x1_ASAP7_75t_L g349 ( 
.A1(n_340),
.A2(n_293),
.B(n_307),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_349),
.B(n_352),
.Y(n_379)
);

INVx11_ASAP7_75t_L g373 ( 
.A(n_351),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_336),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_300),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_353),
.B(n_368),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_341),
.B(n_284),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_354),
.B(n_356),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_336),
.Y(n_355)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_355),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_319),
.B(n_286),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_343),
.B(n_332),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_358),
.B(n_361),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_360),
.A2(n_338),
.B1(n_337),
.B2(n_331),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_345),
.B(n_270),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_362),
.A2(n_339),
.B1(n_344),
.B2(n_288),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_342),
.A2(n_290),
.B1(n_304),
.B2(n_302),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_363),
.A2(n_365),
.B1(n_329),
.B2(n_323),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_342),
.A2(n_304),
.B1(n_302),
.B2(n_298),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_L g366 ( 
.A(n_340),
.B(n_298),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_366),
.A2(n_325),
.B1(n_327),
.B2(n_320),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_326),
.B(n_237),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_322),
.B(n_237),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_334),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_353),
.B(n_333),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_371),
.B(n_372),
.C(n_385),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_321),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_374),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_346),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_375),
.B(n_367),
.Y(n_400)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_348),
.Y(n_376)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_376),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_377),
.A2(n_382),
.B1(n_362),
.B2(n_346),
.Y(n_404)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_348),
.Y(n_378)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_378),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_357),
.A2(n_335),
.B1(n_320),
.B2(n_324),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_381),
.A2(n_357),
.B1(n_355),
.B2(n_352),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_384),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_350),
.B(n_347),
.C(n_359),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_359),
.B(n_316),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_388),
.B(n_389),
.C(n_368),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_347),
.B(n_316),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_376),
.Y(n_390)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_390),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_393),
.B(n_397),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_394),
.B(n_396),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_379),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_370),
.B(n_369),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_400),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_370),
.B(n_349),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_401),
.B(n_402),
.C(n_403),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_365),
.C(n_363),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_371),
.B(n_349),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_404),
.B(n_405),
.Y(n_418)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_378),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_373),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_406),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_402),
.B(n_372),
.C(n_389),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_409),
.B(n_417),
.Y(n_421)
);

BUFx24_ASAP7_75t_SL g412 ( 
.A(n_399),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_412),
.B(n_415),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_396),
.A2(n_379),
.B(n_387),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_414),
.A2(n_390),
.B(n_373),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_391),
.B(n_380),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_388),
.C(n_384),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_410),
.B(n_386),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_420),
.Y(n_430)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_411),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_423),
.B(n_424),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_418),
.A2(n_416),
.B1(n_404),
.B2(n_406),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_407),
.A2(n_405),
.B(n_392),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_425),
.A2(n_427),
.B(n_428),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_407),
.B(n_395),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_426),
.B(n_409),
.C(n_417),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_413),
.A2(n_360),
.B1(n_401),
.B2(n_403),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_414),
.A2(n_395),
.B1(n_398),
.B2(n_392),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_429),
.Y(n_437)
);

AOI322xp5_ASAP7_75t_L g431 ( 
.A1(n_428),
.A2(n_398),
.A3(n_364),
.B1(n_367),
.B2(n_420),
.C1(n_424),
.C2(n_421),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_431),
.A2(n_434),
.B1(n_435),
.B2(n_205),
.Y(n_439)
);

NAND5xp2_ASAP7_75t_L g434 ( 
.A(n_422),
.B(n_377),
.C(n_351),
.D(n_408),
.E(n_393),
.Y(n_434)
);

AOI322xp5_ASAP7_75t_L g435 ( 
.A1(n_427),
.A2(n_351),
.A3(n_382),
.B1(n_364),
.B2(n_397),
.C1(n_383),
.C2(n_408),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_433),
.A2(n_426),
.B(n_351),
.Y(n_436)
);

A2O1A1O1Ixp25_ASAP7_75t_L g442 ( 
.A1(n_436),
.A2(n_432),
.B(n_435),
.C(n_201),
.D(n_223),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_430),
.A2(n_351),
.B1(n_288),
.B2(n_262),
.Y(n_438)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_438),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_439),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_442),
.B(n_440),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_441),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_443),
.B(n_444),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_445),
.A2(n_437),
.B(n_214),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_446),
.B(n_223),
.Y(n_447)
);


endmodule