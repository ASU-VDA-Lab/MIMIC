module real_aes_7214_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_417;
wire n_449;
wire n_363;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_552;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
OAI22xp5_ASAP7_75t_SL g182 ( .A1(n_0), .A2(n_183), .B1(n_184), .B2(n_185), .Y(n_182) );
INVx1_ASAP7_75t_L g185 ( .A(n_0), .Y(n_185) );
INVx1_ASAP7_75t_L g286 ( .A(n_1), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_2), .Y(n_157) );
INVx1_ASAP7_75t_L g168 ( .A(n_3), .Y(n_168) );
AOI22xp33_ASAP7_75t_L g126 ( .A1(n_4), .A2(n_31), .B1(n_127), .B2(n_131), .Y(n_126) );
AOI21xp33_ASAP7_75t_L g297 ( .A1(n_5), .A2(n_216), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g206 ( .A(n_6), .Y(n_206) );
AND2x6_ASAP7_75t_L g221 ( .A(n_6), .B(n_204), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_6), .B(n_544), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_7), .A2(n_266), .B(n_267), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_8), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g303 ( .A(n_9), .Y(n_303) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_10), .A2(n_29), .B1(n_91), .B2(n_96), .Y(n_99) );
INVx1_ASAP7_75t_L g241 ( .A(n_11), .Y(n_241) );
INVx1_ASAP7_75t_L g274 ( .A(n_12), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g84 ( .A1(n_13), .A2(n_50), .B1(n_85), .B2(n_102), .Y(n_84) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_14), .B(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g137 ( .A(n_15), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_16), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_17), .B(n_231), .Y(n_347) );
AO22x2_ASAP7_75t_L g101 ( .A1(n_18), .A2(n_30), .B1(n_91), .B2(n_92), .Y(n_101) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_19), .B(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_20), .B(n_296), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_21), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_22), .A2(n_271), .B(n_273), .C(n_275), .Y(n_270) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_23), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_24), .B(n_256), .Y(n_287) );
AOI22xp5_ASAP7_75t_SL g539 ( .A1(n_24), .A2(n_81), .B1(n_176), .B2(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_24), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_25), .A2(n_81), .B1(n_176), .B2(n_551), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_25), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g106 ( .A1(n_26), .A2(n_53), .B1(n_107), .B2(n_112), .Y(n_106) );
INVx1_ASAP7_75t_L g313 ( .A(n_27), .Y(n_313) );
INVx2_ASAP7_75t_L g219 ( .A(n_28), .Y(n_219) );
OAI221xp5_ASAP7_75t_L g197 ( .A1(n_30), .A2(n_42), .B1(n_52), .B2(n_198), .C(n_199), .Y(n_197) );
INVxp67_ASAP7_75t_L g200 ( .A(n_30), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_32), .A2(n_221), .B(n_223), .C(n_226), .Y(n_222) );
INVx1_ASAP7_75t_L g311 ( .A(n_33), .Y(n_311) );
OAI22xp5_ASAP7_75t_SL g188 ( .A1(n_34), .A2(n_189), .B1(n_190), .B2(n_191), .Y(n_188) );
INVx1_ASAP7_75t_L g190 ( .A(n_34), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_34), .B(n_256), .Y(n_346) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_35), .A2(n_180), .B1(n_181), .B2(n_182), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_35), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_36), .Y(n_150) );
CKINVDCx16_ASAP7_75t_R g314 ( .A(n_37), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_38), .B(n_216), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_39), .A2(n_223), .B1(n_289), .B2(n_310), .Y(n_309) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_40), .Y(n_243) );
CKINVDCx16_ASAP7_75t_R g282 ( .A(n_41), .Y(n_282) );
AO22x2_ASAP7_75t_L g90 ( .A1(n_42), .A2(n_61), .B1(n_91), .B2(n_92), .Y(n_90) );
INVxp67_ASAP7_75t_L g201 ( .A(n_42), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g300 ( .A1(n_43), .A2(n_301), .B(n_302), .C(n_304), .Y(n_300) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_44), .Y(n_350) );
INVx1_ASAP7_75t_L g299 ( .A(n_45), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g117 ( .A1(n_46), .A2(n_51), .B1(n_118), .B2(n_121), .Y(n_117) );
INVx1_ASAP7_75t_L g204 ( .A(n_47), .Y(n_204) );
INVx1_ASAP7_75t_L g240 ( .A(n_48), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_49), .Y(n_198) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_52), .A2(n_66), .B1(n_91), .B2(n_96), .Y(n_95) );
INVxp67_ASAP7_75t_L g189 ( .A(n_54), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_SL g321 ( .A1(n_55), .A2(n_231), .B(n_304), .C(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g184 ( .A(n_56), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g316 ( .A(n_57), .Y(n_316) );
INVx1_ASAP7_75t_L g343 ( .A(n_58), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_59), .A2(n_81), .B1(n_175), .B2(n_176), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_59), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g344 ( .A1(n_60), .A2(n_221), .B(n_223), .C(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_62), .B(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g238 ( .A(n_63), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_64), .B(n_231), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g284 ( .A1(n_65), .A2(n_221), .B(n_223), .C(n_285), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_67), .A2(n_187), .B1(n_188), .B2(n_192), .Y(n_186) );
INVx1_ASAP7_75t_L g192 ( .A(n_67), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_68), .B(n_249), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g292 ( .A(n_69), .Y(n_292) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_70), .A2(n_221), .B(n_223), .C(n_252), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_71), .Y(n_261) );
INVx1_ASAP7_75t_L g320 ( .A(n_72), .Y(n_320) );
CKINVDCx16_ASAP7_75t_R g268 ( .A(n_73), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_74), .B(n_228), .Y(n_253) );
INVx1_ASAP7_75t_L g91 ( .A(n_75), .Y(n_91) );
INVx1_ASAP7_75t_L g93 ( .A(n_75), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_76), .B(n_245), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_77), .A2(n_216), .B(n_319), .Y(n_318) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_194), .B1(n_207), .B2(n_530), .C(n_538), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_177), .Y(n_79) );
INVx1_ASAP7_75t_L g176 ( .A(n_81), .Y(n_176) );
AND2x2_ASAP7_75t_SL g81 ( .A(n_82), .B(n_135), .Y(n_81) );
NOR2xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_116), .Y(n_82) );
NAND2xp33_ASAP7_75t_SL g83 ( .A(n_84), .B(n_106), .Y(n_83) );
BUFx3_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_97), .Y(n_87) );
AND2x6_ASAP7_75t_L g109 ( .A(n_88), .B(n_110), .Y(n_109) );
AND2x4_ASAP7_75t_L g119 ( .A(n_88), .B(n_120), .Y(n_119) );
AND2x6_ASAP7_75t_L g148 ( .A(n_88), .B(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_94), .Y(n_88) );
AND2x2_ASAP7_75t_L g105 ( .A(n_89), .B(n_95), .Y(n_105) );
INVx2_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_90), .B(n_95), .Y(n_115) );
AND2x2_ASAP7_75t_L g124 ( .A(n_90), .B(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g156 ( .A(n_90), .B(n_99), .Y(n_156) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g96 ( .A(n_93), .Y(n_96) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g125 ( .A(n_95), .Y(n_125) );
INVx1_ASAP7_75t_L g155 ( .A(n_95), .Y(n_155) );
AND2x4_ASAP7_75t_L g104 ( .A(n_97), .B(n_105), .Y(n_104) );
AND2x4_ASAP7_75t_L g113 ( .A(n_97), .B(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g123 ( .A(n_97), .B(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g97 ( .A(n_98), .B(n_100), .Y(n_97) );
OR2x2_ASAP7_75t_L g111 ( .A(n_98), .B(n_101), .Y(n_111) );
AND2x2_ASAP7_75t_L g120 ( .A(n_98), .B(n_101), .Y(n_120) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x2_ASAP7_75t_L g149 ( .A(n_99), .B(n_101), .Y(n_149) );
AND2x2_ASAP7_75t_L g154 ( .A(n_100), .B(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g167 ( .A(n_100), .Y(n_167) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g134 ( .A(n_101), .Y(n_134) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g140 ( .A(n_105), .Y(n_140) );
NAND2x1p5_ASAP7_75t_L g143 ( .A(n_105), .B(n_120), .Y(n_143) );
INVx4_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx11_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g139 ( .A(n_111), .B(n_140), .Y(n_139) );
BUFx3_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OR2x6_ASAP7_75t_L g133 ( .A(n_115), .B(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_126), .Y(n_116) );
BUFx3_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g130 ( .A(n_120), .B(n_124), .Y(n_130) );
BUFx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g174 ( .A(n_125), .Y(n_174) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx5_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx8_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx4f_ASAP7_75t_SL g131 ( .A(n_132), .Y(n_131) );
INVx6_ASAP7_75t_SL g132 ( .A(n_133), .Y(n_132) );
NOR3xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_144), .C(n_163), .Y(n_135) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_138), .B1(n_141), .B2(n_142), .Y(n_136) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
OAI221xp5_ASAP7_75t_SL g144 ( .A1(n_145), .A2(n_150), .B1(n_151), .B2(n_157), .C(n_158), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx4_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g172 ( .A(n_149), .Y(n_172) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_154), .B(n_156), .Y(n_153) );
INVx1_ASAP7_75t_L g162 ( .A(n_155), .Y(n_162) );
AND2x4_ASAP7_75t_L g161 ( .A(n_156), .B(n_162), .Y(n_161) );
NAND2x1p5_ASAP7_75t_L g166 ( .A(n_156), .B(n_167), .Y(n_166) );
BUFx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OAI22xp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B1(n_168), .B2(n_169), .Y(n_163) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
CKINVDCx16_ASAP7_75t_R g170 ( .A(n_171), .Y(n_170) );
OR2x6_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
OAI22xp5_ASAP7_75t_SL g177 ( .A1(n_178), .A2(n_179), .B1(n_186), .B2(n_193), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_179), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_182), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_184), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_186), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g191 ( .A(n_189), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_189), .B(n_229), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_195), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_196), .Y(n_195) );
AND3x1_ASAP7_75t_SL g196 ( .A(n_197), .B(n_202), .C(n_205), .Y(n_196) );
INVxp67_ASAP7_75t_L g544 ( .A(n_197), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
INVx1_ASAP7_75t_SL g546 ( .A(n_202), .Y(n_546) );
OAI21xp5_ASAP7_75t_L g548 ( .A1(n_202), .A2(n_533), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g555 ( .A(n_202), .Y(n_555) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_203), .B(n_206), .Y(n_549) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
OR2x2_ASAP7_75t_SL g554 ( .A(n_205), .B(n_555), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_SL g208 ( .A(n_209), .B(n_499), .Y(n_208) );
NOR3xp33_ASAP7_75t_L g209 ( .A(n_210), .B(n_392), .C(n_465), .Y(n_209) );
OAI211xp5_ASAP7_75t_SL g210 ( .A1(n_211), .A2(n_278), .B(n_324), .C(n_376), .Y(n_210) );
INVxp67_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_246), .Y(n_212) );
AND2x2_ASAP7_75t_L g340 ( .A(n_213), .B(n_341), .Y(n_340) );
INVx3_ASAP7_75t_L g359 ( .A(n_213), .Y(n_359) );
INVx2_ASAP7_75t_L g374 ( .A(n_213), .Y(n_374) );
INVx1_ASAP7_75t_L g404 ( .A(n_213), .Y(n_404) );
AND2x2_ASAP7_75t_L g454 ( .A(n_213), .B(n_375), .Y(n_454) );
AOI32xp33_ASAP7_75t_L g481 ( .A1(n_213), .A2(n_409), .A3(n_482), .B1(n_484), .B2(n_485), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_213), .B(n_330), .Y(n_487) );
AND2x2_ASAP7_75t_L g514 ( .A(n_213), .B(n_357), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_213), .B(n_523), .Y(n_522) );
OR2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_242), .Y(n_213) );
AOI21xp5_ASAP7_75t_SL g214 ( .A1(n_215), .A2(n_222), .B(n_235), .Y(n_214) );
BUFx2_ASAP7_75t_L g266 ( .A(n_216), .Y(n_266) );
AND2x4_ASAP7_75t_L g216 ( .A(n_217), .B(n_221), .Y(n_216) );
NAND2x1p5_ASAP7_75t_L g283 ( .A(n_217), .B(n_221), .Y(n_283) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_220), .Y(n_217) );
INVx1_ASAP7_75t_L g535 ( .A(n_218), .Y(n_535) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g224 ( .A(n_219), .Y(n_224) );
INVx1_ASAP7_75t_L g290 ( .A(n_219), .Y(n_290) );
INVx1_ASAP7_75t_L g225 ( .A(n_220), .Y(n_225) );
INVx3_ASAP7_75t_L g229 ( .A(n_220), .Y(n_229) );
INVx1_ASAP7_75t_L g231 ( .A(n_220), .Y(n_231) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_220), .Y(n_256) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_220), .Y(n_272) );
INVx4_ASAP7_75t_SL g276 ( .A(n_221), .Y(n_276) );
BUFx3_ASAP7_75t_L g532 ( .A(n_221), .Y(n_532) );
INVx5_ASAP7_75t_L g269 ( .A(n_223), .Y(n_269) );
AND2x6_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
BUFx3_ASAP7_75t_L g234 ( .A(n_224), .Y(n_234) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_224), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_230), .B(n_232), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g285 ( .A1(n_228), .A2(n_286), .B(n_287), .C(n_288), .Y(n_285) );
INVx5_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_229), .B(n_303), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_232), .A2(n_346), .B(n_347), .Y(n_345) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g275 ( .A(n_234), .Y(n_275) );
INVx1_ASAP7_75t_L g348 ( .A(n_235), .Y(n_348) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_236), .A2(n_281), .B(n_291), .Y(n_280) );
AO21x2_ASAP7_75t_L g307 ( .A1(n_236), .A2(n_308), .B(n_315), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_236), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_237), .Y(n_245) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
AND2x2_ASAP7_75t_SL g249 ( .A(n_238), .B(n_239), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
NOR2xp33_ASAP7_75t_SL g242 ( .A(n_243), .B(n_244), .Y(n_242) );
INVx3_ASAP7_75t_L g296 ( .A(n_244), .Y(n_296) );
INVx4_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
OA21x2_ASAP7_75t_L g317 ( .A1(n_245), .A2(n_318), .B(n_323), .Y(n_317) );
AND2x2_ASAP7_75t_L g403 ( .A(n_246), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g425 ( .A(n_246), .Y(n_425) );
AND2x2_ASAP7_75t_L g510 ( .A(n_246), .B(n_340), .Y(n_510) );
AND2x2_ASAP7_75t_L g513 ( .A(n_246), .B(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_263), .Y(n_246) );
INVx2_ASAP7_75t_L g332 ( .A(n_247), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_247), .B(n_357), .Y(n_363) );
AND2x2_ASAP7_75t_L g373 ( .A(n_247), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g409 ( .A(n_247), .Y(n_409) );
AO21x2_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_250), .B(n_260), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g262 ( .A(n_249), .Y(n_262) );
OA21x2_ASAP7_75t_L g264 ( .A1(n_249), .A2(n_265), .B(n_277), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_259), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B(n_257), .Y(n_252) );
INVx4_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g301 ( .A(n_256), .Y(n_301) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx3_ASAP7_75t_L g304 ( .A(n_258), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_262), .B(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_262), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g351 ( .A(n_263), .B(n_332), .Y(n_351) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g333 ( .A(n_264), .Y(n_333) );
AND2x2_ASAP7_75t_L g375 ( .A(n_264), .B(n_357), .Y(n_375) );
AND2x2_ASAP7_75t_L g444 ( .A(n_264), .B(n_341), .Y(n_444) );
O2A1O1Ixp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_269), .B(n_270), .C(n_276), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g298 ( .A1(n_269), .A2(n_276), .B(n_299), .C(n_300), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_L g319 ( .A1(n_269), .A2(n_276), .B(n_320), .C(n_321), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_271), .B(n_274), .Y(n_273) );
INVx4_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OAI22xp5_ASAP7_75t_SL g310 ( .A1(n_272), .A2(n_311), .B1(n_312), .B2(n_313), .Y(n_310) );
INVx2_ASAP7_75t_L g312 ( .A(n_272), .Y(n_312) );
OAI22xp33_ASAP7_75t_L g308 ( .A1(n_276), .A2(n_283), .B1(n_309), .B2(n_314), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_293), .Y(n_278) );
OR2x2_ASAP7_75t_L g338 ( .A(n_279), .B(n_307), .Y(n_338) );
INVx1_ASAP7_75t_L g417 ( .A(n_279), .Y(n_417) );
AND2x2_ASAP7_75t_L g431 ( .A(n_279), .B(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_279), .B(n_306), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_279), .B(n_429), .Y(n_483) );
AND2x2_ASAP7_75t_L g491 ( .A(n_279), .B(n_492), .Y(n_491) );
INVx3_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx3_ASAP7_75t_L g328 ( .A(n_280), .Y(n_328) );
AND2x2_ASAP7_75t_L g398 ( .A(n_280), .B(n_307), .Y(n_398) );
OAI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B(n_284), .Y(n_281) );
OAI21xp5_ASAP7_75t_L g342 ( .A1(n_283), .A2(n_343), .B(n_344), .Y(n_342) );
OAI322xp33_ASAP7_75t_L g538 ( .A1(n_286), .A2(n_539), .A3(n_541), .B1(n_545), .B2(n_547), .C1(n_550), .C2(n_552), .Y(n_538) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx3_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_293), .B(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g525 ( .A(n_293), .Y(n_525) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_306), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_294), .B(n_369), .Y(n_391) );
OR2x2_ASAP7_75t_L g420 ( .A(n_294), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g452 ( .A(n_294), .B(n_432), .Y(n_452) );
INVx1_ASAP7_75t_SL g472 ( .A(n_294), .Y(n_472) );
AND2x2_ASAP7_75t_L g476 ( .A(n_294), .B(n_337), .Y(n_476) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_SL g329 ( .A(n_295), .B(n_306), .Y(n_329) );
AND2x2_ASAP7_75t_L g336 ( .A(n_295), .B(n_317), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_295), .B(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g379 ( .A(n_295), .B(n_361), .Y(n_379) );
INVx1_ASAP7_75t_SL g386 ( .A(n_295), .Y(n_386) );
BUFx2_ASAP7_75t_L g397 ( .A(n_295), .Y(n_397) );
AND2x2_ASAP7_75t_L g413 ( .A(n_295), .B(n_328), .Y(n_413) );
AND2x2_ASAP7_75t_L g428 ( .A(n_295), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g492 ( .A(n_295), .B(n_307), .Y(n_492) );
OA21x2_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_297), .B(n_305), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_306), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g416 ( .A(n_306), .B(n_417), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g433 ( .A1(n_306), .A2(n_434), .B1(n_437), .B2(n_440), .C(n_445), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_306), .B(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_317), .Y(n_306) );
INVx3_ASAP7_75t_L g361 ( .A(n_307), .Y(n_361) );
INVx2_ASAP7_75t_L g537 ( .A(n_312), .Y(n_537) );
BUFx2_ASAP7_75t_L g371 ( .A(n_317), .Y(n_371) );
AND2x2_ASAP7_75t_L g385 ( .A(n_317), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g402 ( .A(n_317), .Y(n_402) );
OR2x2_ASAP7_75t_L g421 ( .A(n_317), .B(n_361), .Y(n_421) );
INVx3_ASAP7_75t_L g429 ( .A(n_317), .Y(n_429) );
AND2x2_ASAP7_75t_L g432 ( .A(n_317), .B(n_361), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_330), .B1(n_334), .B2(n_339), .C(n_352), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_327), .B(n_401), .Y(n_526) );
OR2x2_ASAP7_75t_L g529 ( .A(n_327), .B(n_360), .Y(n_529) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
OAI221xp5_ASAP7_75t_SL g352 ( .A1(n_328), .A2(n_353), .B1(n_360), .B2(n_362), .C(n_365), .Y(n_352) );
AND2x2_ASAP7_75t_L g369 ( .A(n_328), .B(n_361), .Y(n_369) );
AND2x2_ASAP7_75t_L g377 ( .A(n_328), .B(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_328), .B(n_385), .Y(n_384) );
NAND2x1_ASAP7_75t_L g427 ( .A(n_328), .B(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g479 ( .A(n_328), .B(n_421), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_330), .A2(n_439), .B1(n_468), .B2(n_470), .Y(n_467) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AOI322xp5_ASAP7_75t_L g376 ( .A1(n_331), .A2(n_340), .A3(n_377), .B1(n_380), .B2(n_383), .C1(n_387), .C2(n_390), .Y(n_376) );
OR2x2_ASAP7_75t_L g388 ( .A(n_331), .B(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_332), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g367 ( .A(n_332), .B(n_341), .Y(n_367) );
INVx1_ASAP7_75t_L g382 ( .A(n_332), .Y(n_382) );
AND2x2_ASAP7_75t_L g448 ( .A(n_332), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g358 ( .A(n_333), .B(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g449 ( .A(n_333), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_333), .B(n_357), .Y(n_523) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_337), .B(n_472), .Y(n_471) );
INVx3_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g423 ( .A(n_338), .B(n_370), .Y(n_423) );
OR2x2_ASAP7_75t_L g520 ( .A(n_338), .B(n_371), .Y(n_520) );
INVx1_ASAP7_75t_L g501 ( .A(n_339), .Y(n_501) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_351), .Y(n_339) );
INVx4_ASAP7_75t_L g389 ( .A(n_340), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_340), .B(n_408), .Y(n_414) );
INVx2_ASAP7_75t_L g357 ( .A(n_341), .Y(n_357) );
AO21x2_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_348), .B(n_349), .Y(n_341) );
INVx1_ASAP7_75t_L g439 ( .A(n_351), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_351), .B(n_411), .Y(n_480) );
AOI21xp33_ASAP7_75t_L g426 ( .A1(n_353), .A2(n_427), .B(n_430), .Y(n_426) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_358), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g411 ( .A(n_357), .Y(n_411) );
INVx1_ASAP7_75t_L g438 ( .A(n_357), .Y(n_438) );
INVx1_ASAP7_75t_L g364 ( .A(n_358), .Y(n_364) );
AND2x2_ASAP7_75t_L g366 ( .A(n_358), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g462 ( .A(n_359), .B(n_448), .Y(n_462) );
AND2x2_ASAP7_75t_L g484 ( .A(n_359), .B(n_444), .Y(n_484) );
BUFx2_ASAP7_75t_L g436 ( .A(n_361), .Y(n_436) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
AOI32xp33_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_368), .A3(n_369), .B1(n_370), .B2(n_372), .Y(n_365) );
INVx1_ASAP7_75t_L g446 ( .A(n_366), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_366), .A2(n_494), .B1(n_495), .B2(n_497), .Y(n_493) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_369), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_369), .B(n_428), .Y(n_469) );
AND2x2_ASAP7_75t_L g516 ( .A(n_369), .B(n_401), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_370), .B(n_417), .Y(n_464) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g517 ( .A(n_372), .Y(n_517) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
INVx1_ASAP7_75t_L g442 ( .A(n_373), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_375), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g489 ( .A(n_375), .B(n_409), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_375), .B(n_404), .Y(n_496) );
INVx1_ASAP7_75t_SL g478 ( .A(n_377), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_378), .B(n_429), .Y(n_456) );
NOR4xp25_ASAP7_75t_L g502 ( .A(n_378), .B(n_401), .C(n_503), .D(n_506), .Y(n_502) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_379), .B(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVxp67_ASAP7_75t_L g459 ( .A(n_382), .Y(n_459) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OAI21xp33_ASAP7_75t_L g509 ( .A1(n_385), .A2(n_476), .B(n_510), .Y(n_509) );
AND2x4_ASAP7_75t_L g401 ( .A(n_386), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g450 ( .A(n_389), .Y(n_450) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND4xp25_ASAP7_75t_SL g392 ( .A(n_393), .B(n_418), .C(n_433), .D(n_453), .Y(n_392) );
O2A1O1Ixp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_399), .B(n_403), .C(n_405), .Y(n_393) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_398), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g485 ( .A(n_398), .B(n_428), .Y(n_485) );
AND2x2_ASAP7_75t_L g494 ( .A(n_398), .B(n_472), .Y(n_494) );
INVx3_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_401), .B(n_436), .Y(n_498) );
AND2x2_ASAP7_75t_L g410 ( .A(n_404), .B(n_411), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_412), .B1(n_414), .B2(n_415), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_410), .Y(n_407) );
AND2x2_ASAP7_75t_L g508 ( .A(n_408), .B(n_454), .Y(n_508) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_410), .B(n_459), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_411), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
O2A1O1Ixp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_422), .B(n_424), .C(n_426), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g453 ( .A1(n_419), .A2(n_454), .B1(n_455), .B2(n_457), .C(n_460), .Y(n_453) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OAI221xp5_ASAP7_75t_L g511 ( .A1(n_427), .A2(n_512), .B1(n_515), .B2(n_517), .C(n_518), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_428), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_436), .B(n_505), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g466 ( .A(n_438), .Y(n_466) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_441), .A2(n_461), .B1(n_463), .B2(n_464), .Y(n_460) );
OR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AOI21xp33_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B(n_451), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_450), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_450), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OAI221xp5_ASAP7_75t_L g524 ( .A1(n_461), .A2(n_487), .B1(n_525), .B2(n_526), .C(n_527), .Y(n_524) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g506 ( .A(n_463), .Y(n_506) );
OAI211xp5_ASAP7_75t_SL g465 ( .A1(n_466), .A2(n_467), .B(n_473), .C(n_493), .Y(n_465) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AOI211xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_476), .B(n_477), .C(n_486), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B(n_480), .C(n_481), .Y(n_477) );
INVx1_ASAP7_75t_L g505 ( .A(n_483), .Y(n_505) );
OAI21xp5_ASAP7_75t_SL g527 ( .A1(n_484), .A2(n_510), .B(n_528), .Y(n_527) );
AOI21xp33_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_488), .B(n_490), .Y(n_486) );
INVx1_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
INVxp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OAI21xp5_ASAP7_75t_SL g519 ( .A1(n_496), .A2(n_520), .B(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NOR3xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_511), .C(n_524), .Y(n_499) );
OAI211xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B(n_507), .C(n_509), .Y(n_500) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
CKINVDCx14_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
CKINVDCx16_ASAP7_75t_R g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
CKINVDCx14_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_543), .Y(n_542) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
CKINVDCx16_ASAP7_75t_R g547 ( .A(n_548), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_553), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_554), .Y(n_553) );
endmodule