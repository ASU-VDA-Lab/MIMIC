module real_jpeg_29072_n_16 (n_333, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_333;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_0),
.A2(n_36),
.B1(n_63),
.B2(n_66),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_0),
.A2(n_36),
.B1(n_46),
.B2(n_47),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_1),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_126),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_1),
.A2(n_63),
.B1(n_66),
.B2(n_126),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_126),
.Y(n_264)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_2),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_2),
.A2(n_146),
.B(n_159),
.Y(n_158)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_2),
.Y(n_224)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_4),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_131),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_131),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_4),
.A2(n_63),
.B1(n_66),
.B2(n_131),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_6),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_6),
.A2(n_51),
.B1(n_63),
.B2(n_66),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_51),
.Y(n_284)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_8),
.A2(n_11),
.B(n_63),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_9),
.A2(n_34),
.B1(n_46),
.B2(n_47),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_9),
.A2(n_34),
.B1(n_63),
.B2(n_66),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_54),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_54),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_10),
.A2(n_54),
.B1(n_63),
.B2(n_66),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_11),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_11),
.B(n_32),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_L g176 ( 
.A1(n_11),
.A2(n_32),
.B(n_172),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_129),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_11),
.B(n_89),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_11),
.A2(n_110),
.B1(n_111),
.B2(n_223),
.Y(n_226)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_45),
.Y(n_56)
);

INVx11_ASAP7_75t_SL g65 ( 
.A(n_14),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_15),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_124),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_15),
.A2(n_46),
.B1(n_47),
.B2(n_124),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_15),
.A2(n_63),
.B1(n_66),
.B2(n_124),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_96),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_94),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_81),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_81),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_71),
.C(n_75),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_20),
.A2(n_21),
.B1(n_71),
.B2(n_319),
.Y(n_323)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_38),
.B1(n_39),
.B2(n_70),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_22),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_23),
.A2(n_37),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_23),
.A2(n_37),
.B1(n_137),
.B2(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_23),
.A2(n_264),
.B(n_283),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_24),
.B(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_24),
.A2(n_85),
.B(n_86),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_24),
.A2(n_30),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_24),
.A2(n_86),
.B(n_284),
.Y(n_308)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_25),
.B(n_32),
.Y(n_143)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

HAxp5_ASAP7_75t_SL g128 ( 
.A(n_27),
.B(n_129),
.CON(n_128),
.SN(n_128)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_29),
.A2(n_31),
.B1(n_128),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_30),
.B(n_284),
.Y(n_283)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

AOI32xp33_ASAP7_75t_L g170 ( 
.A1(n_31),
.A2(n_46),
.A3(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_33),
.A2(n_37),
.B(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_35),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_37),
.B(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_37),
.B(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_57),
.B2(n_69),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_41),
.B(n_57),
.C(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_52),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_42),
.A2(n_77),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_50),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_43),
.A2(n_55),
.B1(n_123),
.B2(n_125),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_43),
.A2(n_55),
.B1(n_123),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_43),
.A2(n_55),
.B1(n_155),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_43),
.A2(n_55),
.B1(n_79),
.B2(n_302),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_43)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_44),
.Y(n_171)
);

NAND2xp33_ASAP7_75t_SL g173 ( 
.A(n_44),
.B(n_47),
.Y(n_173)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_47),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_47),
.A2(n_61),
.B(n_129),
.C(n_200),
.Y(n_199)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_50),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_52),
.A2(n_89),
.B(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_57),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_57),
.A2(n_69),
.B1(n_76),
.B2(n_317),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_62),
.B(n_67),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_58),
.A2(n_67),
.B(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_58),
.A2(n_62),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_58),
.A2(n_180),
.B(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_58),
.A2(n_62),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_58),
.A2(n_62),
.B1(n_179),
.B2(n_198),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_58),
.A2(n_62),
.B1(n_105),
.B2(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_58),
.A2(n_119),
.B(n_257),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_66),
.Y(n_62)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_62),
.B(n_129),
.Y(n_221)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_111),
.Y(n_110)
);

BUFx4f_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_66),
.B(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_68),
.B(n_120),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_71),
.C(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_71),
.A2(n_316),
.B1(n_318),
.B2(n_319),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_71),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_75),
.B(n_323),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_76),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B(n_80),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_77),
.A2(n_80),
.B(n_90),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_87),
.B2(n_88),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI321xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_312),
.A3(n_324),
.B1(n_330),
.B2(n_331),
.C(n_333),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_294),
.B(n_311),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_270),
.B(n_293),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_160),
.B(n_247),
.C(n_269),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_147),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_101),
.B(n_147),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_132),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_116),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_103),
.B(n_116),
.C(n_132),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_109),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_104),
.B(n_109),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_106),
.B(n_190),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_108),
.B(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_112),
.B(n_113),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_115),
.Y(n_159)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_110),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_110),
.A2(n_208),
.B(n_209),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_110),
.A2(n_215),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_110),
.A2(n_224),
.B(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_115),
.Y(n_114)
);

INVx11_ASAP7_75t_L g210 ( 
.A(n_111),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_111),
.B(n_129),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_114),
.A2(n_168),
.B(n_169),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_127),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_127),
.B(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_130),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_141),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_134),
.B(n_139),
.C(n_141),
.Y(n_267)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_144),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.C(n_153),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_148),
.A2(n_149),
.B1(n_242),
.B2(n_244),
.Y(n_241)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_153),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.C(n_157),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_154),
.B(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_185),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_156),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_159),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_246),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_239),
.B(n_245),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_191),
.B(n_238),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_181),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_164),
.B(n_181),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_174),
.C(n_177),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_165),
.A2(n_166),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_170),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_168),
.B(n_210),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_168),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_169),
.A2(n_210),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_182),
.B(n_188),
.C(n_189),
.Y(n_240)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_232),
.B(n_237),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_211),
.B(n_231),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_201),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_194),
.B(n_201),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_199),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_195),
.A2(n_196),
.B1(n_199),
.B2(n_218),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_199),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_207),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_206),
.C(n_207),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_208),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_209),
.B(n_255),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_219),
.B(n_230),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_213),
.B(n_217),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_225),
.B(n_229),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_221),
.B(n_222),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_233),
.B(n_234),
.Y(n_237)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_240),
.B(n_241),
.Y(n_245)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_242),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_248),
.B(n_249),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_267),
.B2(n_268),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_258),
.B2(n_259),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_259),
.C(n_268),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_256),
.Y(n_276)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_262),
.C(n_266),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_266),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_267),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_271),
.B(n_272),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_292),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_285),
.B2(n_286),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_286),
.C(n_292),
.Y(n_295)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_276),
.B(n_279),
.C(n_281),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_280),
.Y(n_302)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_287),
.A2(n_288),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_290),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_288),
.A2(n_305),
.B(n_308),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_290),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_295),
.B(n_296),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_309),
.B2(n_310),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_304),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_299),
.B(n_304),
.C(n_310),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B(n_303),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_301),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_314),
.C(n_320),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_303),
.A2(n_314),
.B1(n_315),
.B2(n_329),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_303),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_309),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_322),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_313),
.B(n_322),
.Y(n_331)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_316),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_320),
.A2(n_321),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);


endmodule