module fake_jpeg_6922_n_76 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_76);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_67;
wire n_75;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_8),
.B(n_6),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_10),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_0),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_23),
.A2(n_19),
.B(n_20),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_11),
.B(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_25),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVxp33_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_31),
.B(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_27),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_25),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_13),
.B1(n_16),
.B2(n_24),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_41),
.B(n_46),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_35),
.A2(n_14),
.B1(n_20),
.B2(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_42),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_28),
.C(n_32),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_28),
.A2(n_14),
.B1(n_18),
.B2(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_32),
.B(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_13),
.Y(n_52)
);

NOR2x1_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_36),
.Y(n_49)
);

AO22x1_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_37),
.B1(n_40),
.B2(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_13),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_52),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_41),
.C(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_55),
.B(n_39),
.Y(n_60)
);

AOI322xp5_ASAP7_75t_SL g66 ( 
.A1(n_60),
.A2(n_53),
.A3(n_12),
.B1(n_8),
.B2(n_7),
.C1(n_5),
.C2(n_54),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_49),
.B2(n_50),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_66),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_65),
.B(n_56),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_64),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_62),
.C(n_53),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_61),
.C(n_32),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_68),
.B(n_63),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_71),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_40),
.B(n_69),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_74),
.A2(n_47),
.B1(n_29),
.B2(n_7),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_75),
.B(n_73),
.Y(n_76)
);


endmodule