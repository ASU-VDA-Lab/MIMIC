module real_aes_207_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_789;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g520 ( .A(n_0), .B(n_217), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_1), .B(n_109), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_2), .Y(n_124) );
INVx1_ASAP7_75t_L g151 ( .A(n_3), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_4), .B(n_523), .Y(n_542) );
NAND2xp33_ASAP7_75t_SL g513 ( .A(n_5), .B(n_172), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_6), .B(n_185), .Y(n_208) );
INVx1_ASAP7_75t_L g505 ( .A(n_7), .Y(n_505) );
INVx1_ASAP7_75t_L g242 ( .A(n_8), .Y(n_242) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_9), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_10), .Y(n_259) );
AND2x2_ASAP7_75t_L g540 ( .A(n_11), .B(n_141), .Y(n_540) );
INVx2_ASAP7_75t_L g142 ( .A(n_12), .Y(n_142) );
AND3x1_ASAP7_75t_L g106 ( .A(n_13), .B(n_34), .C(n_107), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_13), .Y(n_119) );
INVx1_ASAP7_75t_L g218 ( .A(n_14), .Y(n_218) );
AOI221x1_ASAP7_75t_L g508 ( .A1(n_15), .A2(n_174), .B1(n_509), .B2(n_511), .C(n_512), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_16), .B(n_523), .Y(n_576) );
INVx1_ASAP7_75t_L g105 ( .A(n_17), .Y(n_105) );
INVx1_ASAP7_75t_L g215 ( .A(n_18), .Y(n_215) );
INVx1_ASAP7_75t_SL g163 ( .A(n_19), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_20), .B(n_166), .Y(n_188) );
AOI33xp33_ASAP7_75t_L g233 ( .A1(n_21), .A2(n_49), .A3(n_148), .B1(n_159), .B2(n_234), .B3(n_235), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_22), .A2(n_511), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_23), .B(n_217), .Y(n_545) );
AOI221xp5_ASAP7_75t_SL g585 ( .A1(n_24), .A2(n_39), .B1(n_511), .B2(n_523), .C(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g252 ( .A(n_25), .Y(n_252) );
OR2x2_ASAP7_75t_L g143 ( .A(n_26), .B(n_88), .Y(n_143) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_26), .A2(n_88), .B(n_142), .Y(n_176) );
INVxp67_ASAP7_75t_L g507 ( .A(n_27), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_28), .B(n_220), .Y(n_580) );
AND2x2_ASAP7_75t_L g534 ( .A(n_29), .B(n_140), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_30), .B(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_31), .A2(n_511), .B(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_32), .B(n_220), .Y(n_587) );
AND2x2_ASAP7_75t_L g153 ( .A(n_33), .B(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g158 ( .A(n_33), .Y(n_158) );
AND2x2_ASAP7_75t_L g172 ( .A(n_33), .B(n_151), .Y(n_172) );
OR2x6_ASAP7_75t_L g121 ( .A(n_34), .B(n_122), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_35), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_36), .B(n_146), .Y(n_279) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_37), .A2(n_175), .B1(n_181), .B2(n_185), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_38), .B(n_190), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_40), .A2(n_80), .B1(n_156), .B2(n_511), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_41), .B(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_42), .B(n_217), .Y(n_532) );
AOI22xp33_ASAP7_75t_SL g788 ( .A1(n_43), .A2(n_787), .B1(n_789), .B2(n_791), .Y(n_788) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_44), .B(n_192), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_45), .B(n_166), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_46), .Y(n_184) );
AND2x2_ASAP7_75t_L g524 ( .A(n_47), .B(n_140), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_48), .B(n_140), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_50), .B(n_166), .Y(n_283) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_51), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_51), .A2(n_61), .B1(n_431), .B2(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g149 ( .A(n_52), .Y(n_149) );
INVx1_ASAP7_75t_L g168 ( .A(n_52), .Y(n_168) );
AND2x2_ASAP7_75t_L g284 ( .A(n_53), .B(n_140), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g240 ( .A1(n_54), .A2(n_72), .B1(n_146), .B2(n_156), .C(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_55), .B(n_146), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_56), .B(n_523), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_57), .B(n_175), .Y(n_261) );
AOI21xp5_ASAP7_75t_SL g197 ( .A1(n_58), .A2(n_156), .B(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g561 ( .A(n_59), .B(n_140), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_60), .B(n_220), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_61), .Y(n_806) );
INVx1_ASAP7_75t_L g211 ( .A(n_62), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_63), .B(n_217), .Y(n_559) );
AND2x2_ASAP7_75t_SL g581 ( .A(n_64), .B(n_141), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_65), .A2(n_511), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g282 ( .A(n_66), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_67), .B(n_220), .Y(n_546) );
AND2x2_ASAP7_75t_SL g553 ( .A(n_68), .B(n_192), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_69), .A2(n_156), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g154 ( .A(n_70), .Y(n_154) );
INVx1_ASAP7_75t_L g170 ( .A(n_70), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_71), .B(n_146), .Y(n_236) );
AND2x2_ASAP7_75t_L g173 ( .A(n_73), .B(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g212 ( .A(n_74), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_75), .A2(n_156), .B(n_162), .Y(n_155) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_76), .A2(n_101), .B1(n_110), .B2(n_808), .Y(n_100) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_77), .A2(n_156), .B(n_187), .C(n_191), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_78), .A2(n_83), .B1(n_146), .B2(n_523), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_79), .B(n_523), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_81), .B(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g123 ( .A(n_81), .Y(n_123) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_82), .B(n_174), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_84), .A2(n_156), .B1(n_231), .B2(n_232), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_85), .B(n_217), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_86), .B(n_217), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_87), .A2(n_511), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g199 ( .A(n_89), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_90), .B(n_220), .Y(n_558) );
AND2x2_ASAP7_75t_L g237 ( .A(n_91), .B(n_174), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_92), .A2(n_250), .B(n_251), .C(n_253), .Y(n_249) );
INVxp67_ASAP7_75t_L g510 ( .A(n_93), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_94), .B(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_95), .B(n_220), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_96), .A2(n_511), .B(n_578), .Y(n_577) );
BUFx2_ASAP7_75t_L g114 ( .A(n_97), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_98), .B(n_166), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_99), .Y(n_787) );
INVx1_ASAP7_75t_SL g808 ( .A(n_101), .Y(n_808) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_SL g103 ( .A(n_104), .B(n_106), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_105), .B(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OA21x2_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_125), .B(n_795), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_115), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_113), .B(n_796), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
INVxp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g796 ( .A1(n_116), .A2(n_797), .B(n_807), .Y(n_796) );
NOR2xp33_ASAP7_75t_SL g116 ( .A(n_117), .B(n_124), .Y(n_116) );
BUFx2_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g807 ( .A(n_118), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
AND2x6_ASAP7_75t_SL g495 ( .A(n_119), .B(n_121), .Y(n_495) );
OR2x6_ASAP7_75t_SL g786 ( .A(n_119), .B(n_120), .Y(n_786) );
OR2x2_ASAP7_75t_L g794 ( .A(n_119), .B(n_121), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_787), .B(n_788), .Y(n_125) );
INVxp67_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22x1_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_494), .B1(n_496), .B2(n_784), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_129), .A2(n_494), .B1(n_497), .B2(n_790), .Y(n_789) );
AND3x1_ASAP7_75t_L g129 ( .A(n_130), .B(n_488), .C(n_491), .Y(n_129) );
NAND5xp2_ASAP7_75t_L g130 ( .A(n_131), .B(n_388), .C(n_418), .D(n_432), .E(n_458), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OAI21xp33_ASAP7_75t_L g488 ( .A1(n_132), .A2(n_431), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g802 ( .A(n_132), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_337), .Y(n_132) );
NOR3xp33_ASAP7_75t_SL g133 ( .A(n_134), .B(n_285), .C(n_319), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_202), .B(n_224), .C(n_263), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_177), .Y(n_135) );
BUFx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_137), .B(n_275), .Y(n_340) );
AND2x2_ASAP7_75t_L g427 ( .A(n_137), .B(n_205), .Y(n_427) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OR2x2_ASAP7_75t_L g223 ( .A(n_138), .B(n_194), .Y(n_223) );
INVx1_ASAP7_75t_L g265 ( .A(n_138), .Y(n_265) );
INVx2_ASAP7_75t_L g270 ( .A(n_138), .Y(n_270) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_138), .Y(n_298) );
INVx1_ASAP7_75t_L g312 ( .A(n_138), .Y(n_312) );
AND2x2_ASAP7_75t_L g316 ( .A(n_138), .B(n_207), .Y(n_316) );
AND2x2_ASAP7_75t_L g397 ( .A(n_138), .B(n_206), .Y(n_397) );
AO21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_144), .B(n_173), .Y(n_138) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_139), .A2(n_528), .B(n_534), .Y(n_527) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_139), .A2(n_555), .B(n_561), .Y(n_554) );
AO21x2_ASAP7_75t_L g592 ( .A1(n_139), .A2(n_528), .B(n_534), .Y(n_592) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_140), .Y(n_139) );
OA21x2_ASAP7_75t_L g584 ( .A1(n_140), .A2(n_585), .B(n_589), .Y(n_584) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_SL g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x4_ASAP7_75t_L g185 ( .A(n_142), .B(n_143), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_155), .Y(n_144) );
INVx1_ASAP7_75t_L g262 ( .A(n_146), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_146), .A2(n_156), .B1(n_504), .B2(n_506), .Y(n_503) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_152), .Y(n_146) );
INVx1_ASAP7_75t_L g182 ( .A(n_147), .Y(n_182) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
OR2x6_ASAP7_75t_L g164 ( .A(n_148), .B(n_160), .Y(n_164) );
INVxp33_ASAP7_75t_L g234 ( .A(n_148), .Y(n_234) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g161 ( .A(n_149), .B(n_151), .Y(n_161) );
AND2x4_ASAP7_75t_L g220 ( .A(n_149), .B(n_169), .Y(n_220) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g183 ( .A(n_152), .Y(n_183) );
BUFx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x6_ASAP7_75t_L g511 ( .A(n_153), .B(n_161), .Y(n_511) );
INVx2_ASAP7_75t_L g160 ( .A(n_154), .Y(n_160) );
AND2x6_ASAP7_75t_L g217 ( .A(n_154), .B(n_167), .Y(n_217) );
INVxp67_ASAP7_75t_L g260 ( .A(n_156), .Y(n_260) );
AND2x4_ASAP7_75t_L g156 ( .A(n_157), .B(n_161), .Y(n_156) );
NOR2x1p5_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
INVx1_ASAP7_75t_L g235 ( .A(n_159), .Y(n_235) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
O2A1O1Ixp33_ASAP7_75t_SL g162 ( .A1(n_163), .A2(n_164), .B(n_165), .C(n_171), .Y(n_162) );
INVx2_ASAP7_75t_L g190 ( .A(n_164), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g198 ( .A1(n_164), .A2(n_171), .B(n_199), .C(n_200), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_164), .A2(n_211), .B1(n_212), .B2(n_213), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_SL g241 ( .A1(n_164), .A2(n_171), .B(n_242), .C(n_243), .Y(n_241) );
INVxp67_ASAP7_75t_L g250 ( .A(n_164), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g281 ( .A1(n_164), .A2(n_171), .B(n_282), .C(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g213 ( .A(n_166), .Y(n_213) );
AND2x4_ASAP7_75t_L g523 ( .A(n_166), .B(n_172), .Y(n_523) );
AND2x4_ASAP7_75t_L g166 ( .A(n_167), .B(n_169), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_171), .A2(n_188), .B(n_189), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_171), .B(n_185), .Y(n_221) );
INVx1_ASAP7_75t_L g231 ( .A(n_171), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_171), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_171), .A2(n_531), .B(n_532), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_171), .A2(n_545), .B(n_546), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_171), .A2(n_558), .B(n_559), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_171), .A2(n_579), .B(n_580), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_171), .A2(n_587), .B(n_588), .Y(n_586) );
INVx5_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_172), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_174), .A2(n_249), .B1(n_254), .B2(n_255), .Y(n_248) );
INVx3_ASAP7_75t_L g255 ( .A(n_174), .Y(n_255) );
INVx4_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_175), .B(n_258), .Y(n_257) );
AOI21x1_ASAP7_75t_L g516 ( .A1(n_175), .A2(n_517), .B(n_524), .Y(n_516) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
BUFx4f_ASAP7_75t_L g192 ( .A(n_176), .Y(n_192) );
AND2x4_ASAP7_75t_SL g177 ( .A(n_178), .B(n_193), .Y(n_177) );
HB1xp67_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g222 ( .A(n_179), .Y(n_222) );
AND2x2_ASAP7_75t_L g266 ( .A(n_179), .B(n_207), .Y(n_266) );
AND2x2_ASAP7_75t_L g287 ( .A(n_179), .B(n_194), .Y(n_287) );
INVx1_ASAP7_75t_L g310 ( .A(n_179), .Y(n_310) );
AND2x4_ASAP7_75t_L g377 ( .A(n_179), .B(n_206), .Y(n_377) );
AND2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_186), .Y(n_179) );
NOR3xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .C(n_184), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_185), .A2(n_197), .B(n_201), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_185), .B(n_505), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_185), .B(n_507), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_185), .B(n_510), .Y(n_509) );
NOR3xp33_ASAP7_75t_L g512 ( .A(n_185), .B(n_213), .C(n_513), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_185), .A2(n_542), .B(n_543), .Y(n_541) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_191), .A2(n_229), .B(n_237), .Y(n_228) );
AO21x2_ASAP7_75t_L g292 ( .A1(n_191), .A2(n_229), .B(n_237), .Y(n_292) );
AOI21x1_ASAP7_75t_L g549 ( .A1(n_191), .A2(n_550), .B(n_553), .Y(n_549) );
INVx2_ASAP7_75t_SL g191 ( .A(n_192), .Y(n_191) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_192), .A2(n_240), .B(n_244), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_192), .A2(n_576), .B(n_577), .Y(n_575) );
AND2x4_ASAP7_75t_L g393 ( .A(n_193), .B(n_310), .Y(n_393) );
OR2x2_ASAP7_75t_L g434 ( .A(n_193), .B(n_435), .Y(n_434) );
NOR2xp67_ASAP7_75t_SL g453 ( .A(n_193), .B(n_326), .Y(n_453) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_193), .B(n_385), .Y(n_471) );
INVx4_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2x1_ASAP7_75t_SL g271 ( .A(n_194), .B(n_207), .Y(n_271) );
AND2x4_ASAP7_75t_L g309 ( .A(n_194), .B(n_310), .Y(n_309) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_194), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_194), .B(n_269), .Y(n_347) );
INVx2_ASAP7_75t_L g361 ( .A(n_194), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g383 ( .A(n_194), .B(n_313), .Y(n_383) );
AND2x2_ASAP7_75t_L g475 ( .A(n_194), .B(n_333), .Y(n_475) );
OR2x6_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2x1_ASAP7_75t_L g203 ( .A(n_204), .B(n_223), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_205), .B(n_312), .Y(n_326) );
AND2x2_ASAP7_75t_SL g335 ( .A(n_205), .B(n_315), .Y(n_335) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_222), .Y(n_205) );
INVx1_ASAP7_75t_L g313 ( .A(n_206), .Y(n_313) );
INVx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g333 ( .A(n_207), .Y(n_333) );
AND2x4_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_214), .B(n_221), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_213), .B(n_252), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B1(n_218), .B2(n_219), .Y(n_214) );
INVxp67_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVxp67_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g366 ( .A(n_222), .Y(n_366) );
INVx2_ASAP7_75t_SL g411 ( .A(n_223), .Y(n_411) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_245), .Y(n_225) );
NAND2x1p5_ASAP7_75t_L g320 ( .A(n_226), .B(n_321), .Y(n_320) );
BUFx2_ASAP7_75t_L g357 ( .A(n_226), .Y(n_357) );
AND2x2_ASAP7_75t_L g481 ( .A(n_226), .B(n_306), .Y(n_481) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_238), .Y(n_226) );
AND2x4_ASAP7_75t_L g294 ( .A(n_227), .B(n_276), .Y(n_294) );
INVx1_ASAP7_75t_L g305 ( .A(n_227), .Y(n_305) );
AND2x2_ASAP7_75t_L g336 ( .A(n_227), .B(n_291), .Y(n_336) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_228), .B(n_239), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_228), .B(n_277), .Y(n_368) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_230), .B(n_236), .Y(n_229) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVxp67_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g274 ( .A(n_239), .Y(n_274) );
AND2x4_ASAP7_75t_L g342 ( .A(n_239), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g354 ( .A(n_239), .Y(n_354) );
INVx1_ASAP7_75t_L g396 ( .A(n_239), .Y(n_396) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_239), .Y(n_408) );
AND2x2_ASAP7_75t_L g424 ( .A(n_239), .B(n_247), .Y(n_424) );
BUFx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g371 ( .A(n_246), .B(n_329), .Y(n_371) );
INVx1_ASAP7_75t_SL g373 ( .A(n_246), .Y(n_373) );
AND2x2_ASAP7_75t_L g394 ( .A(n_246), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x4_ASAP7_75t_L g273 ( .A(n_247), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g301 ( .A(n_247), .Y(n_301) );
INVx2_ASAP7_75t_L g307 ( .A(n_247), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_247), .B(n_277), .Y(n_322) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_256), .Y(n_247) );
AO21x2_ASAP7_75t_L g277 ( .A1(n_255), .A2(n_278), .B(n_284), .Y(n_277) );
AO21x2_ASAP7_75t_L g291 ( .A1(n_255), .A2(n_278), .B(n_284), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_260), .B1(n_261), .B2(n_262), .Y(n_256) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_267), .B(n_272), .Y(n_263) );
INVx1_ASAP7_75t_L g403 ( .A(n_264), .Y(n_403) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g323 ( .A(n_266), .Y(n_323) );
AND2x2_ASAP7_75t_L g379 ( .A(n_266), .B(n_315), .Y(n_379) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_271), .Y(n_267) );
INVx1_ASAP7_75t_L g293 ( .A(n_268), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_268), .B(n_309), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_268), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g400 ( .A(n_268), .B(n_393), .Y(n_400) );
AND2x2_ASAP7_75t_L g474 ( .A(n_268), .B(n_475), .Y(n_474) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_269), .Y(n_462) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_270), .Y(n_382) );
AND2x2_ASAP7_75t_L g295 ( .A(n_271), .B(n_296), .Y(n_295) );
OAI21xp33_ASAP7_75t_L g483 ( .A1(n_271), .A2(n_484), .B(n_486), .Y(n_483) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
INVx3_ASAP7_75t_L g369 ( .A(n_273), .Y(n_369) );
NAND2x1_ASAP7_75t_SL g413 ( .A(n_273), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g416 ( .A(n_273), .B(n_294), .Y(n_416) );
AND2x2_ASAP7_75t_L g328 ( .A(n_275), .B(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g465 ( .A(n_275), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g476 ( .A(n_275), .B(n_424), .Y(n_476) );
INVx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2x1p5_ASAP7_75t_L g352 ( .A(n_276), .B(n_353), .Y(n_352) );
INVx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g407 ( .A(n_277), .B(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
OAI21xp5_ASAP7_75t_SL g285 ( .A1(n_286), .A2(n_299), .B(n_302), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_288), .B1(n_294), .B2(n_295), .Y(n_286) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_287), .Y(n_344) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_293), .Y(n_288) );
AND2x2_ASAP7_75t_L g317 ( .A(n_289), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g423 ( .A(n_289), .B(n_424), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_289), .A2(n_442), .B1(n_443), .B2(n_444), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_289), .B(n_450), .Y(n_449) );
AND2x4_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g306 ( .A(n_291), .B(n_307), .Y(n_306) );
NOR2xp67_ASAP7_75t_L g387 ( .A(n_291), .B(n_307), .Y(n_387) );
NOR2x1_ASAP7_75t_L g395 ( .A(n_291), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g343 ( .A(n_292), .Y(n_343) );
AND2x2_ASAP7_75t_L g351 ( .A(n_292), .B(n_307), .Y(n_351) );
INVx1_ASAP7_75t_L g414 ( .A(n_292), .Y(n_414) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2x1_ASAP7_75t_L g332 ( .A(n_297), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g444 ( .A(n_300), .B(n_329), .Y(n_444) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g318 ( .A(n_301), .Y(n_318) );
AND2x2_ASAP7_75t_L g341 ( .A(n_301), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g429 ( .A(n_301), .B(n_336), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_308), .B1(n_314), .B2(n_317), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g437 ( .A(n_304), .B(n_438), .Y(n_437) );
NAND2x1p5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
AND2x2_ASAP7_75t_L g467 ( .A(n_307), .B(n_354), .Y(n_467) );
AND2x2_ASAP7_75t_SL g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx2_ASAP7_75t_L g334 ( .A(n_309), .Y(n_334) );
OAI21xp33_ASAP7_75t_SL g480 ( .A1(n_309), .A2(n_481), .B(n_482), .Y(n_480) );
AND2x4_ASAP7_75t_SL g311 ( .A(n_312), .B(n_313), .Y(n_311) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_312), .Y(n_470) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
O2A1O1Ixp33_ASAP7_75t_SL g412 ( .A1(n_315), .A2(n_413), .B(n_415), .C(n_417), .Y(n_412) );
AND2x2_ASAP7_75t_SL g364 ( .A(n_316), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g417 ( .A(n_316), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_316), .B(n_393), .Y(n_457) );
INVx1_ASAP7_75t_SL g324 ( .A(n_317), .Y(n_324) );
AND2x2_ASAP7_75t_L g405 ( .A(n_318), .B(n_342), .Y(n_405) );
INVx1_ASAP7_75t_L g450 ( .A(n_318), .Y(n_450) );
OAI221xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_323), .B1(n_324), .B2(n_325), .C(n_327), .Y(n_319) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_320), .Y(n_439) );
INVx2_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g487 ( .A(n_322), .B(n_330), .Y(n_487) );
OR2x2_ASAP7_75t_L g346 ( .A(n_323), .B(n_347), .Y(n_346) );
NOR2x1_ASAP7_75t_L g359 ( .A(n_323), .B(n_360), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_323), .B(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g485 ( .A(n_323), .B(n_382), .Y(n_485) );
BUFx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI32xp33_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_331), .A3(n_334), .B1(n_335), .B2(n_336), .Y(n_327) );
INVx1_ASAP7_75t_L g348 ( .A(n_329), .Y(n_348) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_331), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g443 ( .A(n_332), .Y(n_443) );
OAI22xp33_ASAP7_75t_SL g425 ( .A1(n_334), .A2(n_426), .B1(n_428), .B2(n_430), .Y(n_425) );
INVx1_ASAP7_75t_L g456 ( .A(n_335), .Y(n_456) );
AOI211x1_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_344), .B(n_345), .C(n_362), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_339), .B(n_424), .Y(n_430) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g386 ( .A(n_342), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g452 ( .A(n_342), .Y(n_452) );
OAI222xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_348), .B1(n_349), .B2(n_355), .C1(n_356), .C2(n_358), .Y(n_345) );
INVxp67_ASAP7_75t_L g442 ( .A(n_346), .Y(n_442) );
OR2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_350), .B(n_435), .Y(n_482) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g398 ( .A(n_351), .B(n_395), .Y(n_398) );
INVx3_ASAP7_75t_L g438 ( .A(n_353), .Y(n_438) );
BUFx3_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g376 ( .A(n_361), .B(n_377), .Y(n_376) );
OAI221xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_367), .B1(n_370), .B2(n_375), .C(n_378), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
OAI21xp5_ASAP7_75t_L g420 ( .A1(n_364), .A2(n_421), .B(n_423), .Y(n_420) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g374 ( .A(n_368), .Y(n_374) );
OR2x2_ASAP7_75t_L g478 ( .A(n_369), .B(n_414), .Y(n_478) );
NOR2xp67_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_372), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
OAI21xp5_ASAP7_75t_L g472 ( .A1(n_375), .A2(n_404), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_376), .A2(n_448), .B(n_455), .Y(n_454) );
INVx4_ASAP7_75t_L g385 ( .A(n_377), .Y(n_385) );
OAI31xp33_ASAP7_75t_SL g378 ( .A1(n_379), .A2(n_380), .A3(n_384), .B(n_386), .Y(n_378) );
INVx1_ASAP7_75t_L g436 ( .A(n_380), .Y(n_436) );
NOR2x1_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g410 ( .A(n_385), .Y(n_410) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_401), .Y(n_388) );
NAND4xp25_ASAP7_75t_L g489 ( .A(n_389), .B(n_401), .C(n_420), .D(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_399), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_394), .B1(n_397), .B2(n_398), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g461 ( .A(n_393), .B(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_394), .B(n_414), .Y(n_422) );
INVx1_ASAP7_75t_SL g435 ( .A(n_397), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_402), .B(n_412), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B1(n_406), .B2(n_409), .Y(n_402) );
INVx3_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVxp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2x1_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_411), .A2(n_474), .B1(n_476), .B2(n_477), .Y(n_473) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NOR3xp33_ASAP7_75t_L g418 ( .A(n_419), .B(n_425), .C(n_431), .Y(n_418) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g490 ( .A(n_425), .Y(n_490) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI21xp33_ASAP7_75t_L g491 ( .A1(n_431), .A2(n_492), .B(n_493), .Y(n_491) );
INVxp33_ASAP7_75t_L g492 ( .A(n_432), .Y(n_492) );
AND2x2_ASAP7_75t_L g801 ( .A(n_432), .B(n_458), .Y(n_801) );
NOR2xp67_ASAP7_75t_L g432 ( .A(n_433), .B(n_440), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_436), .B1(n_437), .B2(n_439), .Y(n_433) );
OAI21xp5_ASAP7_75t_L g459 ( .A1(n_437), .A2(n_460), .B(n_463), .Y(n_459) );
INVx2_ASAP7_75t_L g447 ( .A(n_438), .Y(n_447) );
NAND3xp33_ASAP7_75t_SL g440 ( .A(n_441), .B(n_445), .C(n_454), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_448), .B1(n_451), .B2(n_453), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
INVxp33_ASAP7_75t_SL g493 ( .A(n_458), .Y(n_493) );
NOR3x1_ASAP7_75t_L g458 ( .A(n_459), .B(n_472), .C(n_479), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_468), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_480), .B(n_483), .Y(n_479) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g803 ( .A(n_489), .Y(n_803) );
CKINVDCx11_ASAP7_75t_R g494 ( .A(n_495), .Y(n_494) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_498), .B(n_661), .Y(n_497) );
NOR4xp25_ASAP7_75t_L g498 ( .A(n_499), .B(n_604), .C(n_643), .D(n_650), .Y(n_498) );
OAI221xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_525), .B1(n_562), .B2(n_571), .C(n_590), .Y(n_499) );
OR2x2_ASAP7_75t_L g734 ( .A(n_500), .B(n_596), .Y(n_734) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g649 ( .A(n_501), .B(n_574), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_501), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_SL g714 ( .A(n_501), .B(n_715), .Y(n_714) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_514), .Y(n_501) );
AND2x4_ASAP7_75t_SL g573 ( .A(n_502), .B(n_574), .Y(n_573) );
INVx3_ASAP7_75t_L g595 ( .A(n_502), .Y(n_595) );
AND2x2_ASAP7_75t_L g630 ( .A(n_502), .B(n_603), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_502), .B(n_515), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_502), .B(n_597), .Y(n_682) );
OR2x2_ASAP7_75t_L g760 ( .A(n_502), .B(n_574), .Y(n_760) );
AND2x4_ASAP7_75t_L g502 ( .A(n_503), .B(n_508), .Y(n_502) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g582 ( .A(n_515), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_515), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g608 ( .A(n_515), .Y(n_608) );
OR2x2_ASAP7_75t_L g613 ( .A(n_515), .B(n_597), .Y(n_613) );
AND2x2_ASAP7_75t_L g626 ( .A(n_515), .B(n_584), .Y(n_626) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_515), .Y(n_629) );
INVx1_ASAP7_75t_L g641 ( .A(n_515), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_515), .B(n_595), .Y(n_706) );
INVx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_522), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_526), .B(n_535), .Y(n_525) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g570 ( .A(n_527), .B(n_554), .Y(n_570) );
AND2x4_ASAP7_75t_L g600 ( .A(n_527), .B(n_539), .Y(n_600) );
INVx2_ASAP7_75t_L g634 ( .A(n_527), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_527), .B(n_554), .Y(n_692) );
AND2x2_ASAP7_75t_L g739 ( .A(n_527), .B(n_568), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_533), .Y(n_528) );
AOI222xp33_ASAP7_75t_L g727 ( .A1(n_535), .A2(n_599), .B1(n_642), .B2(n_702), .C1(n_728), .C2(n_730), .Y(n_727) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_547), .Y(n_536) );
AND2x2_ASAP7_75t_L g646 ( .A(n_537), .B(n_566), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_537), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g775 ( .A(n_537), .B(n_615), .Y(n_775) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_538), .A2(n_606), .B(n_610), .Y(n_605) );
AND2x2_ASAP7_75t_L g686 ( .A(n_538), .B(n_569), .Y(n_686) );
OR2x2_ASAP7_75t_L g711 ( .A(n_538), .B(n_570), .Y(n_711) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx5_ASAP7_75t_L g565 ( .A(n_539), .Y(n_565) );
AND2x2_ASAP7_75t_L g652 ( .A(n_539), .B(n_634), .Y(n_652) );
AND2x2_ASAP7_75t_L g678 ( .A(n_539), .B(n_554), .Y(n_678) );
OR2x2_ASAP7_75t_L g681 ( .A(n_539), .B(n_568), .Y(n_681) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_539), .Y(n_699) );
AND2x4_ASAP7_75t_SL g756 ( .A(n_539), .B(n_633), .Y(n_756) );
OR2x2_ASAP7_75t_L g765 ( .A(n_539), .B(n_592), .Y(n_765) );
OR2x6_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
INVx1_ASAP7_75t_L g598 ( .A(n_547), .Y(n_598) );
AOI221xp5_ASAP7_75t_SL g716 ( .A1(n_547), .A2(n_600), .B1(n_717), .B2(n_719), .C(n_720), .Y(n_716) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_554), .Y(n_547) );
OR2x2_ASAP7_75t_L g655 ( .A(n_548), .B(n_625), .Y(n_655) );
OR2x2_ASAP7_75t_L g665 ( .A(n_548), .B(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g691 ( .A(n_548), .B(n_692), .Y(n_691) );
AND2x4_ASAP7_75t_L g697 ( .A(n_548), .B(n_616), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_548), .B(n_680), .Y(n_709) );
INVx2_ASAP7_75t_L g722 ( .A(n_548), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g743 ( .A(n_548), .B(n_600), .Y(n_743) );
AND2x2_ASAP7_75t_L g747 ( .A(n_548), .B(n_569), .Y(n_747) );
AND2x2_ASAP7_75t_L g755 ( .A(n_548), .B(n_756), .Y(n_755) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g568 ( .A(n_549), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_554), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g599 ( .A(n_554), .B(n_568), .Y(n_599) );
INVx2_ASAP7_75t_L g616 ( .A(n_554), .Y(n_616) );
AND2x4_ASAP7_75t_L g633 ( .A(n_554), .B(n_634), .Y(n_633) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_554), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_560), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_563), .B(n_566), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g745 ( .A(n_564), .B(n_567), .Y(n_745) );
AND2x4_ASAP7_75t_L g591 ( .A(n_565), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g632 ( .A(n_565), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g659 ( .A(n_565), .B(n_599), .Y(n_659) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
AND2x2_ASAP7_75t_L g763 ( .A(n_567), .B(n_764), .Y(n_763) );
BUFx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g615 ( .A(n_568), .B(n_616), .Y(n_615) );
OAI21xp5_ASAP7_75t_SL g635 ( .A1(n_569), .A2(n_636), .B(n_642), .Y(n_635) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_582), .Y(n_572) );
INVx1_ASAP7_75t_SL g689 ( .A(n_573), .Y(n_689) );
AND2x2_ASAP7_75t_L g719 ( .A(n_573), .B(n_629), .Y(n_719) );
AND2x4_ASAP7_75t_L g730 ( .A(n_573), .B(n_731), .Y(n_730) );
OR2x2_ASAP7_75t_L g596 ( .A(n_574), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g603 ( .A(n_574), .Y(n_603) );
AND2x4_ASAP7_75t_L g609 ( .A(n_574), .B(n_595), .Y(n_609) );
INVx2_ASAP7_75t_L g620 ( .A(n_574), .Y(n_620) );
INVx1_ASAP7_75t_L g669 ( .A(n_574), .Y(n_669) );
OR2x2_ASAP7_75t_L g690 ( .A(n_574), .B(n_674), .Y(n_690) );
OR2x2_ASAP7_75t_L g704 ( .A(n_574), .B(n_584), .Y(n_704) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_574), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_574), .B(n_626), .Y(n_776) );
OR2x6_ASAP7_75t_L g574 ( .A(n_575), .B(n_581), .Y(n_574) );
INVx1_ASAP7_75t_L g621 ( .A(n_582), .Y(n_621) );
AND2x2_ASAP7_75t_L g754 ( .A(n_582), .B(n_620), .Y(n_754) );
AND2x2_ASAP7_75t_L g779 ( .A(n_582), .B(n_609), .Y(n_779) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g597 ( .A(n_584), .Y(n_597) );
BUFx3_ASAP7_75t_L g639 ( .A(n_584), .Y(n_639) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_584), .Y(n_666) );
INVx1_ASAP7_75t_L g675 ( .A(n_584), .Y(n_675) );
AOI33xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_593), .A3(n_598), .B1(n_599), .B2(n_600), .B3(n_601), .Y(n_590) );
AOI21x1_ASAP7_75t_SL g693 ( .A1(n_591), .A2(n_615), .B(n_677), .Y(n_693) );
INVx2_ASAP7_75t_L g723 ( .A(n_591), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_591), .B(n_722), .Y(n_729) );
AND2x2_ASAP7_75t_L g677 ( .A(n_592), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
AND2x2_ASAP7_75t_L g640 ( .A(n_595), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g741 ( .A(n_596), .Y(n_741) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_597), .Y(n_731) );
OAI32xp33_ASAP7_75t_L g780 ( .A1(n_598), .A2(n_600), .A3(n_776), .B1(n_781), .B2(n_783), .Y(n_780) );
AND2x2_ASAP7_75t_L g698 ( .A(n_599), .B(n_699), .Y(n_698) );
INVx2_ASAP7_75t_SL g688 ( .A(n_600), .Y(n_688) );
AND2x2_ASAP7_75t_L g753 ( .A(n_600), .B(n_697), .Y(n_753) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI221xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_614), .B1(n_617), .B2(n_631), .C(n_635), .Y(n_604) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_608), .B(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_609), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_609), .B(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_609), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g658 ( .A(n_613), .Y(n_658) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NOR3xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_622), .C(n_627), .Y(n_617) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g720 ( .A1(n_619), .A2(n_681), .B1(n_721), .B2(n_724), .Y(n_720) );
OR2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx1_ASAP7_75t_L g624 ( .A(n_620), .Y(n_624) );
NOR2x1p5_ASAP7_75t_L g638 ( .A(n_620), .B(n_639), .Y(n_638) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_620), .Y(n_660) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI322xp33_ASAP7_75t_L g687 ( .A1(n_623), .A2(n_665), .A3(n_688), .B1(n_689), .B2(n_690), .C1(n_691), .C2(n_693), .Y(n_687) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
A2O1A1Ixp33_ASAP7_75t_L g643 ( .A1(n_625), .A2(n_644), .B(n_645), .C(n_647), .Y(n_643) );
OR2x2_ASAP7_75t_L g735 ( .A(n_625), .B(n_689), .Y(n_735) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g642 ( .A(n_626), .B(n_630), .Y(n_642) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g648 ( .A(n_632), .B(n_649), .Y(n_648) );
INVx3_ASAP7_75t_SL g680 ( .A(n_633), .Y(n_680) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_637), .B(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_SL g684 ( .A(n_640), .Y(n_684) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_641), .Y(n_726) );
OR2x6_ASAP7_75t_SL g781 ( .A(n_644), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVxp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AOI211xp5_ASAP7_75t_L g771 ( .A1(n_649), .A2(n_772), .B(n_773), .C(n_780), .Y(n_771) );
O2A1O1Ixp33_ASAP7_75t_SL g650 ( .A1(n_651), .A2(n_653), .B(n_656), .C(n_660), .Y(n_650) );
OAI211xp5_ASAP7_75t_SL g662 ( .A1(n_651), .A2(n_663), .B(n_670), .C(n_694), .Y(n_662) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx3_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
NOR3xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_707), .C(n_751), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_667), .Y(n_663) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_666), .Y(n_758) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g713 ( .A(n_669), .Y(n_713) );
NOR3xp33_ASAP7_75t_SL g670 ( .A(n_671), .B(n_683), .C(n_687), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_676), .B1(n_679), .B2(n_682), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g715 ( .A(n_675), .Y(n_715) );
INVxp67_ASAP7_75t_SL g782 ( .A(n_675), .Y(n_782) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
INVx1_ASAP7_75t_SL g768 ( .A(n_681), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
OR2x2_ASAP7_75t_L g718 ( .A(n_684), .B(n_704), .Y(n_718) );
OR2x2_ASAP7_75t_L g769 ( .A(n_684), .B(n_770), .Y(n_769) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g767 ( .A(n_692), .Y(n_767) );
OR2x2_ASAP7_75t_L g783 ( .A(n_692), .B(n_722), .Y(n_783) );
OAI21xp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_698), .B(n_700), .Y(n_694) );
OAI31xp33_ASAP7_75t_L g708 ( .A1(n_695), .A2(n_709), .A3(n_710), .B(n_712), .Y(n_708) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_705), .Y(n_702) );
INVx1_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
AND2x4_ASAP7_75t_L g740 ( .A(n_705), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND4xp25_ASAP7_75t_SL g707 ( .A(n_708), .B(n_716), .C(n_727), .D(n_732), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_715), .Y(n_750) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
OR2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVxp67_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AOI221xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_736), .B1(n_740), .B2(n_742), .C(n_744), .Y(n_732) );
NAND2xp33_ASAP7_75t_SL g733 ( .A(n_734), .B(n_735), .Y(n_733) );
INVx1_ASAP7_75t_L g777 ( .A(n_736), .Y(n_777) );
AND2x2_ASAP7_75t_SL g736 ( .A(n_737), .B(n_739), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AOI21xp33_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B(n_748), .Y(n_744) );
INVx1_ASAP7_75t_L g772 ( .A(n_746), .Y(n_772) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g751 ( .A(n_752), .B(n_771), .Y(n_751) );
AOI221xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B1(n_755), .B2(n_757), .C(n_761), .Y(n_752) );
AND2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
INVx1_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
AOI21xp33_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_766), .B(n_769), .Y(n_761) );
INVxp33_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_776), .B1(n_777), .B2(n_778), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
CKINVDCx5p33_ASAP7_75t_R g784 ( .A(n_785), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_785), .Y(n_790) );
CKINVDCx11_ASAP7_75t_R g785 ( .A(n_786), .Y(n_785) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_792), .Y(n_791) );
CKINVDCx5p33_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
INVx3_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
OAI22xp33_ASAP7_75t_SL g797 ( .A1(n_798), .A2(n_799), .B1(n_804), .B2(n_805), .Y(n_797) );
INVxp67_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NAND3x1_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .C(n_803), .Y(n_800) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
endmodule