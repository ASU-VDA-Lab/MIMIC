module fake_jpeg_21334_n_280 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_182;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_0),
.C(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_38),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_0),
.C(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_44),
.Y(n_49)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_18),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_61),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_18),
.B1(n_31),
.B2(n_24),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_56),
.B1(n_64),
.B2(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_18),
.B1(n_31),
.B2(n_24),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_59),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_60),
.B(n_34),
.Y(n_67)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_31),
.B1(n_41),
.B2(n_26),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_66),
.A2(n_73),
.B1(n_78),
.B2(n_94),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_42),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_70),
.A2(n_79),
.B(n_82),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_40),
.B1(n_41),
.B2(n_26),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_72),
.A2(n_91),
.B1(n_101),
.B2(n_92),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_40),
.B1(n_17),
.B2(n_19),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_74),
.B(n_86),
.Y(n_121)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_42),
.B1(n_37),
.B2(n_38),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_39),
.B1(n_27),
.B2(n_34),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_39),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_84),
.B(n_93),
.Y(n_119)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_92),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_19),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_87),
.Y(n_105)
);

NAND3xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_30),
.C(n_21),
.Y(n_88)
);

OR2x2_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_97),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_26),
.B1(n_39),
.B2(n_30),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_100),
.B1(n_34),
.B2(n_27),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_58),
.A2(n_17),
.B1(n_25),
.B2(n_35),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_25),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_35),
.B1(n_32),
.B2(n_21),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_36),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_95),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_63),
.B(n_36),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_27),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_103),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_52),
.A2(n_39),
.B1(n_32),
.B2(n_28),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_47),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_52),
.B(n_34),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_78),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_50),
.B(n_34),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_108),
.B1(n_110),
.B2(n_124),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_76),
.A2(n_34),
.B1(n_28),
.B2(n_23),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_69),
.A2(n_28),
.B1(n_23),
.B2(n_33),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_122),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_70),
.A2(n_28),
.B1(n_2),
.B2(n_3),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_116),
.A2(n_128),
.B1(n_84),
.B2(n_81),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_103),
.C(n_69),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_100),
.A2(n_33),
.B1(n_29),
.B2(n_20),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_126),
.A2(n_131),
.B1(n_87),
.B2(n_82),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_70),
.A2(n_10),
.B1(n_2),
.B2(n_4),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_29),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_79),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_76),
.A2(n_29),
.B1(n_20),
.B2(n_4),
.Y(n_131)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_136),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_102),
.B(n_120),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_134),
.A2(n_143),
.B(n_151),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_89),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_135),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_127),
.Y(n_136)
);

INVx2_ASAP7_75t_R g137 ( 
.A(n_109),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_149),
.Y(n_162)
);

OR2x4_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_99),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_104),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_SL g170 ( 
.A1(n_141),
.A2(n_112),
.B(n_83),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_1),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_107),
.A2(n_82),
.B(n_79),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_99),
.B1(n_80),
.B2(n_68),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_144),
.A2(n_150),
.B1(n_157),
.B2(n_9),
.Y(n_183)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_148),
.Y(n_173)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_96),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_147),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_75),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_75),
.B(n_80),
.C(n_79),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_20),
.B(n_1),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_116),
.B(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_106),
.A2(n_110),
.B1(n_124),
.B2(n_132),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_10),
.B1(n_6),
.B2(n_7),
.Y(n_176)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_122),
.A2(n_77),
.B1(n_85),
.B2(n_90),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_119),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_159),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_105),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_175),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_169),
.B(n_170),
.Y(n_189)
);

AND2x6_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_105),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_163),
.B(n_164),
.Y(n_192)
);

CKINVDCx12_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_123),
.C(n_114),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_158),
.C(n_141),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_112),
.Y(n_169)
);

AND2x4_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_114),
.Y(n_174)
);

XOR2x2_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_139),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_10),
.B(n_2),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_176),
.A2(n_150),
.B1(n_144),
.B2(n_157),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_151),
.A2(n_11),
.B1(n_7),
.B2(n_8),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_180),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_8),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_185),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_183),
.A2(n_152),
.B1(n_138),
.B2(n_146),
.Y(n_199)
);

AO21x1_ASAP7_75t_L g185 ( 
.A1(n_134),
.A2(n_9),
.B(n_11),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_188),
.A2(n_204),
.B1(n_177),
.B2(n_166),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_186),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_200),
.Y(n_215)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_165),
.C(n_174),
.Y(n_223)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_196),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_197),
.A2(n_171),
.B(n_161),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_202),
.B1(n_203),
.B2(n_161),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_168),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_138),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_179),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_169),
.A2(n_136),
.B1(n_156),
.B2(n_153),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_183),
.A2(n_145),
.B1(n_159),
.B2(n_133),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_140),
.B1(n_12),
.B2(n_13),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_206),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_140),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_172),
.Y(n_225)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_208),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_204),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_209),
.B(n_224),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_212),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_194),
.B(n_162),
.Y(n_212)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_171),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_220),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_216),
.A2(n_190),
.B(n_185),
.Y(n_240)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_218),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_162),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_203),
.A2(n_174),
.B1(n_163),
.B2(n_181),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_197),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_174),
.C(n_189),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_228),
.C(n_230),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_192),
.C(n_187),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_206),
.C(n_189),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_234),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_215),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_193),
.C(n_198),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_220),
.C(n_198),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_238),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_240),
.A2(n_221),
.B(n_235),
.Y(n_248)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_241),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_217),
.B(n_190),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_242),
.B(n_238),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_211),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_247),
.Y(n_256)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_239),
.Y(n_246)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_248),
.A2(n_231),
.B1(n_237),
.B2(n_224),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_249),
.A2(n_229),
.B(n_233),
.Y(n_254)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_240),
.Y(n_250)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_236),
.C(n_233),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_255),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_248),
.A2(n_231),
.B1(n_213),
.B2(n_188),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_261),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_251),
.C(n_244),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_253),
.A2(n_210),
.B1(n_216),
.B2(n_228),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_265),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_256),
.A2(n_249),
.B(n_243),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_263),
.A2(n_260),
.B(n_258),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_251),
.C(n_252),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_229),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_258),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_268),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

AOI31xp67_ASAP7_75t_L g273 ( 
.A1(n_269),
.A2(n_271),
.A3(n_267),
.B(n_264),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_273),
.A2(n_208),
.B1(n_182),
.B2(n_257),
.Y(n_276)
);

NAND3xp33_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_219),
.C(n_245),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_241),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_276),
.C(n_218),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_277),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_272),
.C(n_180),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_279),
.B(n_11),
.Y(n_280)
);


endmodule