module fake_jpeg_22345_n_171 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_171);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_2),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_39),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_20),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_50),
.Y(n_60)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_31),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_5),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_52),
.B(n_21),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_28),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_56),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_22),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_61),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_22),
.B1(n_50),
.B2(n_16),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_69),
.B1(n_75),
.B2(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_44),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_63),
.B(n_67),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_40),
.B(n_32),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_27),
.B1(n_30),
.B2(n_29),
.Y(n_85)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

AND2x6_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_3),
.Y(n_68)
);

OAI32xp33_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_72),
.A3(n_74),
.B1(n_29),
.B2(n_24),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_37),
.B1(n_32),
.B2(n_36),
.Y(n_69)
);

AND2x6_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_4),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_5),
.B(n_6),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_73),
.A2(n_27),
.B1(n_7),
.B2(n_29),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_36),
.B1(n_38),
.B2(n_26),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_25),
.B1(n_16),
.B2(n_18),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_48),
.A2(n_25),
.B1(n_19),
.B2(n_18),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_82),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_79),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_21),
.B1(n_26),
.B2(n_19),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_23),
.B1(n_30),
.B2(n_29),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_49),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_55),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_30),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_85),
.A2(n_89),
.B1(n_92),
.B2(n_96),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_91),
.Y(n_111)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_102),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_38),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_62),
.Y(n_116)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_97),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

XNOR2x1_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_78),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_118),
.C(n_119),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_66),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_110),
.B(n_84),
.Y(n_127)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_114),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_78),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_91),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_87),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_65),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_72),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_90),
.B(n_102),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_123),
.B(n_127),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_133),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_112),
.C(n_119),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_68),
.C(n_92),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_130),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_109),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_132),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_93),
.B1(n_124),
.B2(n_107),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_137),
.B1(n_144),
.B2(n_96),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_142),
.C(n_81),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_132),
.A2(n_117),
.B1(n_105),
.B2(n_106),
.Y(n_137)
);

NAND2x1_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_113),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_141),
.A2(n_126),
.B1(n_95),
.B2(n_62),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_125),
.B1(n_120),
.B2(n_130),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_135),
.A2(n_123),
.B(n_121),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_147),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_146),
.A2(n_144),
.B1(n_100),
.B2(n_17),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_148),
.B(n_149),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_70),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_143),
.B(n_83),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_151),
.B(n_139),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_139),
.B(n_70),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_141),
.C(n_142),
.Y(n_157)
);

OAI21x1_ASAP7_75t_L g159 ( 
.A1(n_155),
.A2(n_145),
.B(n_9),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_137),
.B1(n_134),
.B2(n_136),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_158),
.B1(n_30),
.B2(n_24),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_17),
.Y(n_160)
);

AOI221xp5_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_160),
.B1(n_158),
.B2(n_11),
.C(n_12),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_153),
.A2(n_13),
.B(n_9),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_154),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_14),
.B(n_10),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_165),
.A2(n_166),
.B(n_167),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_157),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_159),
.A2(n_12),
.A3(n_14),
.B1(n_24),
.B2(n_23),
.C1(n_77),
.C2(n_7),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_166),
.C(n_77),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_168),
.Y(n_171)
);


endmodule