module fake_jpeg_14171_n_131 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_4),
.B(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_35),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_50),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_44),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_22),
.C(n_18),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_29),
.A2(n_24),
.B1(n_20),
.B2(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_29),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_24),
.B1(n_19),
.B2(n_18),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_22),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_29),
.A2(n_19),
.B1(n_21),
.B2(n_18),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_46),
.Y(n_61)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_52),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_63),
.Y(n_80)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_61),
.B1(n_67),
.B2(n_31),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_68),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_64),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_47),
.B(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_65),
.B(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_44),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_36),
.B1(n_18),
.B2(n_21),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_16),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_41),
.C(n_39),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_74),
.C(n_79),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_41),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_81),
.B1(n_69),
.B2(n_61),
.Y(n_86)
);

AND2x6_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_10),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_82),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_45),
.C(n_42),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_49),
.B1(n_53),
.B2(n_26),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_26),
.B(n_14),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_63),
.C(n_60),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_67),
.C(n_57),
.Y(n_92)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_93),
.B1(n_94),
.B2(n_42),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_65),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_83),
.B(n_68),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_92),
.C(n_70),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_28),
.Y(n_102)
);

AO22x1_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_67),
.B1(n_59),
.B2(n_62),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_95),
.B(n_23),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_61),
.B1(n_67),
.B2(n_64),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_73),
.A2(n_67),
.B1(n_36),
.B2(n_54),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_54),
.B1(n_53),
.B2(n_14),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_105),
.Y(n_108)
);

AOI31xp33_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_72),
.A3(n_76),
.B(n_81),
.Y(n_97)
);

OAI321xp33_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_89),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C(n_0),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_92),
.A2(n_71),
.B1(n_18),
.B2(n_53),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_104),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_91),
.A2(n_42),
.B1(n_28),
.B2(n_27),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_102),
.A2(n_2),
.B(n_3),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_27),
.B1(n_23),
.B2(n_16),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_103),
.B(n_84),
.Y(n_106)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

AOI221xp5_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_89),
.B1(n_95),
.B2(n_85),
.C(n_4),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

OA21x2_ASAP7_75t_SL g114 ( 
.A1(n_110),
.A2(n_102),
.B(n_100),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_0),
.C(n_2),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_113),
.C(n_104),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_101),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_6),
.C(n_7),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_114),
.A2(n_115),
.B1(n_118),
.B2(n_107),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_99),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_117),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_108),
.C(n_98),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_121),
.C(n_115),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_108),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_119),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

AOI322xp5_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_126),
.A3(n_120),
.B1(n_122),
.B2(n_98),
.C1(n_9),
.C2(n_8),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_116),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_6),
.C(n_9),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_127),
.A2(n_124),
.B(n_7),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_130),
.Y(n_131)
);


endmodule