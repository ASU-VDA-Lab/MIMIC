module fake_netlist_6_4777_n_1764 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1764);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1764;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_811;
wire n_683;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g155 ( 
.A(n_14),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_77),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_129),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_43),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_4),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_128),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_133),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_36),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_154),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_48),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_82),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_34),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_0),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_37),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_74),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_47),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_69),
.Y(n_176)
);

BUFx10_ASAP7_75t_L g177 ( 
.A(n_54),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_53),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_35),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_70),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_44),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_59),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_37),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_71),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_136),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_127),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_48),
.Y(n_188)
);

BUFx2_ASAP7_75t_SL g189 ( 
.A(n_86),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_101),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_97),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_135),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_56),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_150),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_62),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_44),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_16),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_120),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_75),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_64),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_38),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_104),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_65),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_68),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_106),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_63),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_66),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_25),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_134),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_124),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_4),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_102),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_72),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_79),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_16),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_51),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_153),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_131),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_98),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_84),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_28),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_96),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_50),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_46),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_23),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_100),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_61),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_14),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_26),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_9),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_90),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_24),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_105),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_88),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_114),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_94),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_35),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_51),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_47),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_118),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g242 ( 
.A(n_18),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_109),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_146),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_139),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_45),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_116),
.Y(n_247)
);

BUFx5_ASAP7_75t_L g248 ( 
.A(n_113),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_0),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_30),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_89),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_34),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_42),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_49),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_27),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_52),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_143),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_25),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_49),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_60),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_107),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_19),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_41),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_67),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_5),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_57),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_22),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_22),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_149),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_92),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_121),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_12),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_32),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_78),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_111),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_108),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_39),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_91),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_3),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_17),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_43),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_103),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_12),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_31),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_142),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_19),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_125),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_7),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_151),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_83),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_122),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_15),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_15),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_31),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_28),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_45),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_21),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_138),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_29),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_10),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_152),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_46),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_85),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_5),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_13),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_76),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_50),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_80),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_197),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_225),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_157),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_225),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_157),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_242),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_208),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_208),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_225),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_289),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_225),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_168),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_290),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_225),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_162),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_225),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_242),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_225),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g327 ( 
.A(n_155),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_176),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_242),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_160),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_161),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_209),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_209),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_209),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_209),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_212),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_212),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_160),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_212),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_212),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_304),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_304),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_262),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_199),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_161),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_262),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_292),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_292),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_164),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_165),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_175),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_239),
.Y(n_352)
);

INVxp33_ASAP7_75t_L g353 ( 
.A(n_184),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_239),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_199),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_216),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_217),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_176),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_176),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_222),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_224),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_181),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_183),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_226),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_185),
.Y(n_365)
);

INVxp33_ASAP7_75t_SL g366 ( 
.A(n_300),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_233),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_238),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_249),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_210),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_168),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_156),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_252),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_253),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_259),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_176),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_186),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_166),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_332),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_R g380 ( 
.A(n_318),
.B(n_187),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_320),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_340),
.B(n_205),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_310),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_320),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_310),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_332),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_333),
.Y(n_387)
);

AND2x2_ASAP7_75t_SL g388 ( 
.A(n_321),
.B(n_192),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_311),
.A2(n_163),
.B1(n_240),
.B2(n_182),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_312),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_320),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_320),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_328),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_333),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_312),
.Y(n_395)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_329),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_372),
.B(n_205),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_320),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_317),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_371),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_328),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_378),
.B(n_232),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_371),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_315),
.B(n_232),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_348),
.B(n_192),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_315),
.B(n_298),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_334),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_315),
.B(n_298),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_323),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_315),
.B(n_308),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_349),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_358),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_317),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_316),
.B(n_221),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_334),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_319),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_358),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_319),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_335),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_315),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_371),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_322),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_371),
.B(n_221),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_362),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_322),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_335),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_371),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_343),
.B(n_301),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_359),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_359),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_336),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_336),
.Y(n_432)
);

NOR2x1_ASAP7_75t_L g433 ( 
.A(n_331),
.B(n_189),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_313),
.A2(n_240),
.B1(n_284),
.B2(n_258),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_324),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_363),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_324),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_338),
.A2(n_182),
.B1(n_284),
.B2(n_258),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_326),
.B(n_301),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_337),
.B(n_308),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_376),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_376),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_337),
.B(n_191),
.Y(n_443)
);

BUFx10_ASAP7_75t_L g444 ( 
.A(n_409),
.Y(n_444)
);

AOI21x1_ASAP7_75t_L g445 ( 
.A1(n_439),
.A2(n_326),
.B(n_339),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_388),
.B(n_345),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_383),
.Y(n_447)
);

BUFx10_ASAP7_75t_L g448 ( 
.A(n_409),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_430),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_430),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_388),
.B(n_365),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_414),
.B(n_377),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_L g453 ( 
.A(n_397),
.B(n_195),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_423),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_388),
.B(n_345),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_423),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_398),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_388),
.B(n_366),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_430),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_393),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_414),
.B(n_321),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_404),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_430),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_423),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_383),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_383),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_423),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g468 ( 
.A1(n_414),
.A2(n_281),
.B1(n_352),
.B2(n_354),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_423),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_430),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_404),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_423),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_437),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_406),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_393),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_L g476 ( 
.A(n_397),
.B(n_204),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_393),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_389),
.Y(n_478)
);

INVx8_ASAP7_75t_L g479 ( 
.A(n_439),
.Y(n_479)
);

INVxp33_ASAP7_75t_L g480 ( 
.A(n_389),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_411),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_383),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_405),
.B(n_343),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_430),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_385),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_434),
.B(n_344),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_430),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_411),
.B(n_309),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_424),
.B(n_314),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_437),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_420),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_437),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_385),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_385),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_385),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_398),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_436),
.B(n_325),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_398),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_390),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_436),
.B(n_433),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_430),
.Y(n_501)
);

NAND3xp33_ASAP7_75t_L g502 ( 
.A(n_402),
.B(n_354),
.C(n_352),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_390),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_380),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g505 ( 
.A(n_434),
.Y(n_505)
);

NOR2xp67_ASAP7_75t_L g506 ( 
.A(n_393),
.B(n_339),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_390),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_393),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_396),
.Y(n_509)
);

NOR2x1p5_ASAP7_75t_L g510 ( 
.A(n_402),
.B(n_331),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_401),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_401),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_401),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_396),
.A2(n_303),
.B1(n_215),
.B2(n_241),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_433),
.B(n_330),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_390),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_398),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_401),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_401),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_380),
.B(n_355),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_420),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_405),
.B(n_428),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_412),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_395),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_406),
.B(n_206),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_441),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_439),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_398),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_395),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_441),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_395),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_396),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_395),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_408),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_441),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_408),
.B(n_214),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_399),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_399),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_412),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_399),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_399),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_413),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_413),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_420),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_413),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_441),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_410),
.A2(n_158),
.B1(n_261),
.B2(n_303),
.Y(n_547)
);

INVx5_ASAP7_75t_L g548 ( 
.A(n_441),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_443),
.B(n_327),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_412),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_410),
.B(n_219),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_405),
.B(n_215),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_413),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_439),
.A2(n_281),
.B1(n_288),
.B2(n_293),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_416),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_441),
.Y(n_556)
);

BUFx4f_ASAP7_75t_L g557 ( 
.A(n_441),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_443),
.B(n_241),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_416),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_382),
.B(n_220),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_416),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_416),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_382),
.B(n_243),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_428),
.B(n_346),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_418),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_418),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_418),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_418),
.Y(n_568)
);

AND3x2_ASAP7_75t_L g569 ( 
.A(n_428),
.B(n_306),
.C(n_172),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_420),
.B(n_427),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_412),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_439),
.B(n_306),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_427),
.B(n_223),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_441),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_440),
.B(n_353),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_422),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_442),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_422),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_L g579 ( 
.A(n_440),
.B(n_227),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_422),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_427),
.B(n_228),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_438),
.Y(n_582)
);

INVx5_ASAP7_75t_L g583 ( 
.A(n_442),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_427),
.B(n_235),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_439),
.B(n_243),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_381),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_379),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_412),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_442),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_379),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_462),
.B(n_422),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_462),
.A2(n_471),
.B1(n_474),
.B2(n_534),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_460),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_471),
.B(n_425),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_474),
.B(n_425),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_454),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_491),
.Y(n_597)
);

INVx8_ASAP7_75t_L g598 ( 
.A(n_479),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_460),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_458),
.B(n_425),
.Y(n_600)
);

AND2x6_ASAP7_75t_L g601 ( 
.A(n_522),
.B(n_171),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_534),
.B(n_425),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_549),
.B(n_435),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_L g604 ( 
.A(n_525),
.B(n_536),
.Y(n_604)
);

INVxp33_ASAP7_75t_L g605 ( 
.A(n_575),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_522),
.B(n_435),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_454),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_475),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_509),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_452),
.B(n_461),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_456),
.Y(n_611)
);

AO22x2_ASAP7_75t_L g612 ( 
.A1(n_547),
.A2(n_250),
.B1(n_299),
.B2(n_263),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_587),
.B(n_435),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_451),
.B(n_435),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_464),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_464),
.B(n_442),
.Y(n_616)
);

OA21x2_ASAP7_75t_L g617 ( 
.A1(n_473),
.A2(n_384),
.B(n_381),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_509),
.B(n_346),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_479),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_587),
.B(n_381),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_590),
.B(n_384),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_467),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_510),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_481),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_475),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_570),
.A2(n_391),
.B(n_384),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_467),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_520),
.B(n_488),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_446),
.A2(n_247),
.B1(n_261),
.B2(n_370),
.Y(n_629)
);

NAND3xp33_ASAP7_75t_L g630 ( 
.A(n_502),
.B(n_167),
.C(n_159),
.Y(n_630)
);

INVxp33_ASAP7_75t_L g631 ( 
.A(n_486),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_551),
.A2(n_392),
.B(n_391),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_455),
.B(n_247),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_475),
.Y(n_634)
);

AO22x2_ASAP7_75t_L g635 ( 
.A1(n_552),
.A2(n_265),
.B1(n_267),
.B2(n_280),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_477),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_590),
.B(n_391),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_504),
.B(n_236),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_560),
.B(n_245),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_532),
.B(n_347),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_469),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_477),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_469),
.B(n_392),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_477),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_472),
.B(n_392),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_472),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_473),
.B(n_400),
.Y(n_647)
);

A2O1A1Ixp33_ASAP7_75t_L g648 ( 
.A1(n_490),
.A2(n_234),
.B(n_271),
.C(n_270),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_563),
.B(n_169),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_558),
.B(n_170),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_490),
.B(n_400),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_492),
.B(n_400),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_492),
.B(n_403),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_508),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_483),
.B(n_251),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_508),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_510),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_585),
.B(n_180),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_564),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_564),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_508),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_527),
.B(n_442),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_586),
.Y(n_663)
);

BUFx4_ASAP7_75t_L g664 ( 
.A(n_486),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_483),
.B(n_403),
.Y(n_665)
);

BUFx5_ASAP7_75t_L g666 ( 
.A(n_527),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_586),
.B(n_403),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_586),
.B(n_442),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_527),
.B(n_442),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_527),
.B(n_442),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_500),
.B(n_188),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_515),
.B(n_532),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_572),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_572),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_453),
.B(n_198),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_572),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_511),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_491),
.B(n_417),
.Y(n_678)
);

O2A1O1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_476),
.A2(n_307),
.B(n_302),
.C(n_347),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_521),
.B(n_417),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_450),
.B(n_176),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_468),
.B(n_202),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_450),
.B(n_176),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_521),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_L g685 ( 
.A1(n_479),
.A2(n_285),
.B1(n_278),
.B2(n_173),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_521),
.B(n_417),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_544),
.B(n_417),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_450),
.B(n_176),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_511),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_579),
.B(n_229),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_489),
.B(n_230),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_544),
.B(n_417),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_450),
.B(n_248),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_512),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_544),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_444),
.B(n_256),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_497),
.B(n_231),
.Y(n_697)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_514),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_573),
.B(n_581),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_569),
.B(n_350),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_444),
.Y(n_701)
);

AND2x6_ASAP7_75t_SL g702 ( 
.A(n_478),
.B(n_350),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_444),
.B(n_264),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_444),
.B(n_266),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_448),
.B(n_274),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_514),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_554),
.A2(n_163),
.B1(n_211),
.B2(n_203),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_512),
.Y(n_708)
);

AND2x6_ASAP7_75t_SL g709 ( 
.A(n_478),
.B(n_351),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_448),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_512),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_513),
.Y(n_712)
);

AO22x2_ASAP7_75t_L g713 ( 
.A1(n_480),
.A2(n_213),
.B1(n_269),
.B2(n_260),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_459),
.B(n_429),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_459),
.B(n_248),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_459),
.B(n_248),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_448),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_445),
.B(n_351),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_479),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_459),
.B(n_429),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_513),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_448),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_582),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_584),
.B(n_246),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_505),
.A2(n_201),
.B1(n_174),
.B2(n_178),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_513),
.Y(n_726)
);

OAI221xp5_ASAP7_75t_L g727 ( 
.A1(n_493),
.A2(n_207),
.B1(n_200),
.B2(n_196),
.C(n_194),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_518),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_557),
.A2(n_398),
.B(n_421),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_463),
.B(n_429),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_518),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_479),
.B(n_275),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_493),
.B(n_254),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_518),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_519),
.Y(n_735)
);

OAI22xp33_ASAP7_75t_L g736 ( 
.A1(n_494),
.A2(n_300),
.B1(n_305),
.B2(n_268),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_463),
.B(n_470),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_494),
.B(n_255),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_470),
.B(n_386),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_457),
.B(n_276),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_519),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_519),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_499),
.B(n_272),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_470),
.B(n_386),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_445),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_523),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_470),
.B(n_387),
.Y(n_747)
);

AND2x6_ASAP7_75t_L g748 ( 
.A(n_487),
.B(n_179),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_487),
.B(n_501),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_523),
.Y(n_750)
);

OAI22xp33_ASAP7_75t_L g751 ( 
.A1(n_499),
.A2(n_305),
.B1(n_297),
.B2(n_296),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_487),
.B(n_248),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_523),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_487),
.B(n_248),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_506),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_659),
.B(n_356),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_605),
.B(n_438),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_610),
.B(n_557),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_596),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_618),
.B(n_356),
.Y(n_760)
);

NAND3xp33_ASAP7_75t_L g761 ( 
.A(n_650),
.B(n_277),
.C(n_273),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_610),
.B(n_507),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_598),
.Y(n_763)
);

INVx4_ASAP7_75t_L g764 ( 
.A(n_598),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_592),
.B(n_557),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_640),
.B(n_357),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_607),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_600),
.A2(n_557),
.B(n_484),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_598),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_R g770 ( 
.A(n_701),
.B(n_282),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_611),
.Y(n_771)
);

BUFx12f_ASAP7_75t_L g772 ( 
.A(n_702),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_603),
.B(n_507),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_615),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_622),
.Y(n_775)
);

OAI22xp33_ASAP7_75t_L g776 ( 
.A1(n_629),
.A2(n_660),
.B1(n_628),
.B2(n_698),
.Y(n_776)
);

INVx5_ASAP7_75t_L g777 ( 
.A(n_619),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_600),
.A2(n_484),
.B(n_449),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_722),
.Y(n_779)
);

BUFx4f_ASAP7_75t_L g780 ( 
.A(n_628),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_672),
.B(n_287),
.Y(n_781)
);

AND2x4_ASAP7_75t_SL g782 ( 
.A(n_710),
.B(n_161),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_609),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_606),
.B(n_516),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_623),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_602),
.B(n_516),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_591),
.B(n_524),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_627),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_672),
.B(n_357),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_594),
.B(n_524),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_641),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_646),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_663),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_597),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_593),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_673),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_657),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_724),
.B(n_619),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_723),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_674),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_700),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_724),
.A2(n_526),
.B1(n_501),
.B2(n_535),
.Y(n_802)
);

AND2x6_ASAP7_75t_L g803 ( 
.A(n_699),
.B(n_501),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_595),
.B(n_529),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_676),
.Y(n_805)
);

NOR2x1p5_ASAP7_75t_L g806 ( 
.A(n_624),
.B(n_630),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_599),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_658),
.A2(n_526),
.B1(n_501),
.B2(n_535),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_699),
.B(n_529),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_665),
.B(n_538),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_700),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_619),
.B(n_291),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_682),
.B(n_360),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_649),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_649),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_628),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_608),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_633),
.B(n_706),
.Y(n_818)
);

BUFx2_ASAP7_75t_L g819 ( 
.A(n_709),
.Y(n_819)
);

AOI22x1_ASAP7_75t_L g820 ( 
.A1(n_745),
.A2(n_526),
.B1(n_535),
.B2(n_546),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_745),
.B(n_538),
.Y(n_821)
);

CKINVDCx11_ASAP7_75t_R g822 ( 
.A(n_664),
.Y(n_822)
);

OR2x2_ASAP7_75t_L g823 ( 
.A(n_682),
.B(n_360),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_658),
.A2(n_526),
.B1(n_535),
.B2(n_546),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_619),
.B(n_457),
.Y(n_825)
);

OR2x6_ASAP7_75t_L g826 ( 
.A(n_717),
.B(n_361),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_614),
.B(n_540),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_614),
.B(n_540),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_719),
.B(n_457),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_643),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_597),
.B(n_684),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_635),
.Y(n_832)
);

BUFx4f_ASAP7_75t_L g833 ( 
.A(n_601),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_645),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_650),
.B(n_449),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_635),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_691),
.B(n_449),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_718),
.B(n_543),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_635),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_638),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_718),
.B(n_543),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_625),
.Y(n_842)
);

AND2x6_ASAP7_75t_L g843 ( 
.A(n_719),
.B(n_546),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_691),
.B(n_484),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_655),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_604),
.B(n_553),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_697),
.B(n_530),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_719),
.B(n_457),
.Y(n_848)
);

OR2x2_ASAP7_75t_L g849 ( 
.A(n_631),
.B(n_361),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_R g850 ( 
.A(n_695),
.B(n_671),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_721),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_719),
.B(n_457),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_726),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_613),
.B(n_553),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_734),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_748),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_725),
.B(n_555),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_666),
.B(n_457),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_725),
.B(n_555),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_731),
.B(n_559),
.Y(n_860)
);

NAND3xp33_ASAP7_75t_SL g861 ( 
.A(n_707),
.B(n_286),
.C(n_283),
.Y(n_861)
);

OR2x6_ASAP7_75t_L g862 ( 
.A(n_713),
.B(n_364),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_697),
.Y(n_863)
);

INVx5_ASAP7_75t_L g864 ( 
.A(n_601),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_735),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_620),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_601),
.A2(n_546),
.B1(n_556),
.B2(n_574),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_634),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_696),
.B(n_364),
.Y(n_869)
);

INVx1_ASAP7_75t_SL g870 ( 
.A(n_713),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_713),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_666),
.B(n_496),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_742),
.B(n_559),
.Y(n_873)
);

AO22x1_ASAP7_75t_L g874 ( 
.A1(n_671),
.A2(n_279),
.B1(n_295),
.B2(n_294),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_621),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_750),
.B(n_753),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_612),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_636),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_707),
.A2(n_257),
.B1(n_190),
.B2(n_244),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_612),
.B(n_367),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_642),
.Y(n_881)
);

AND2x6_ASAP7_75t_SL g882 ( 
.A(n_690),
.B(n_367),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_703),
.B(n_530),
.Y(n_883)
);

NOR2x1p5_ASAP7_75t_L g884 ( 
.A(n_637),
.B(n_368),
.Y(n_884)
);

NAND2x1p5_ASAP7_75t_L g885 ( 
.A(n_662),
.B(n_556),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_662),
.A2(n_589),
.B(n_530),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_612),
.B(n_368),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_667),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_739),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_704),
.B(n_530),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_705),
.B(n_369),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_601),
.A2(n_562),
.B1(n_566),
.B2(n_565),
.Y(n_892)
);

AO22x1_ASAP7_75t_L g893 ( 
.A1(n_690),
.A2(n_193),
.B1(n_218),
.B2(n_237),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_644),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_666),
.B(n_617),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_675),
.A2(n_574),
.B1(n_556),
.B2(n_577),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_733),
.B(n_369),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_744),
.Y(n_898)
);

AND2x2_ASAP7_75t_SL g899 ( 
.A(n_675),
.B(n_373),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_748),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_639),
.B(n_577),
.Y(n_901)
);

OR2x2_ASAP7_75t_SL g902 ( 
.A(n_736),
.B(n_373),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_748),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_666),
.B(n_562),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_666),
.B(n_565),
.Y(n_905)
);

OR2x2_ASAP7_75t_SL g906 ( 
.A(n_736),
.B(n_374),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_666),
.B(n_566),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_747),
.Y(n_908)
);

CKINVDCx6p67_ASAP7_75t_R g909 ( 
.A(n_748),
.Y(n_909)
);

AND2x6_ASAP7_75t_SL g910 ( 
.A(n_733),
.B(n_374),
.Y(n_910)
);

AND3x1_ASAP7_75t_L g911 ( 
.A(n_679),
.B(n_375),
.C(n_341),
.Y(n_911)
);

BUFx4f_ASAP7_75t_L g912 ( 
.A(n_748),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_617),
.B(n_567),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_647),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_651),
.Y(n_915)
);

INVx5_ASAP7_75t_L g916 ( 
.A(n_654),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_617),
.Y(n_917)
);

INVx5_ASAP7_75t_L g918 ( 
.A(n_656),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_652),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_616),
.B(n_375),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_653),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_738),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_661),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_738),
.B(n_496),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_751),
.B(n_577),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_616),
.B(n_574),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_743),
.Y(n_927)
);

INVxp67_ASAP7_75t_SL g928 ( 
.A(n_669),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_677),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_743),
.B(n_751),
.Y(n_930)
);

OR2x6_ASAP7_75t_L g931 ( 
.A(n_681),
.B(n_341),
.Y(n_931)
);

NAND2x1p5_ASAP7_75t_L g932 ( 
.A(n_669),
.B(n_577),
.Y(n_932)
);

INVx4_ASAP7_75t_L g933 ( 
.A(n_689),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_694),
.Y(n_934)
);

BUFx4f_ASAP7_75t_L g935 ( 
.A(n_708),
.Y(n_935)
);

AND2x2_ASAP7_75t_SL g936 ( 
.A(n_678),
.B(n_342),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_711),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_712),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_904),
.A2(n_670),
.B(n_668),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_811),
.B(n_816),
.Y(n_940)
);

BUFx10_ASAP7_75t_L g941 ( 
.A(n_882),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_775),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_814),
.B(n_755),
.Y(n_943)
);

A2O1A1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_930),
.A2(n_626),
.B(n_632),
.C(n_680),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_760),
.B(n_342),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_759),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_783),
.Y(n_947)
);

OAI21xp33_ASAP7_75t_L g948 ( 
.A1(n_813),
.A2(n_727),
.B(n_648),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_788),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_830),
.B(n_728),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_815),
.B(n_749),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_794),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_794),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_922),
.B(n_741),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_899),
.A2(n_670),
.B1(n_686),
.B2(n_687),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_904),
.A2(n_737),
.B(n_732),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_R g957 ( 
.A(n_779),
.B(n_692),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_905),
.A2(n_749),
.B(n_589),
.Y(n_958)
);

O2A1O1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_879),
.A2(n_685),
.B(n_752),
.C(n_715),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_905),
.A2(n_589),
.B(n_729),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_897),
.B(n_746),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_923),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_794),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_834),
.B(n_714),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_766),
.B(n_681),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_822),
.Y(n_966)
);

BUFx12f_ASAP7_75t_L g967 ( 
.A(n_772),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_907),
.A2(n_740),
.B(n_720),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_798),
.A2(n_730),
.B(n_528),
.Y(n_969)
);

OR2x6_ASAP7_75t_L g970 ( 
.A(n_799),
.B(n_763),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_801),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_849),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_923),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_758),
.A2(n_809),
.B(n_784),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_795),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_767),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_927),
.B(n_683),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_807),
.Y(n_978)
);

NOR3xp33_ASAP7_75t_SL g979 ( 
.A(n_757),
.B(n_754),
.C(n_752),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_777),
.Y(n_980)
);

OR2x6_ASAP7_75t_L g981 ( 
.A(n_763),
.B(n_683),
.Y(n_981)
);

INVx6_ASAP7_75t_L g982 ( 
.A(n_806),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_789),
.B(n_567),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_809),
.A2(n_528),
.B(n_517),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_771),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_863),
.B(n_688),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_914),
.B(n_578),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_850),
.B(n_818),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_762),
.A2(n_870),
.B1(n_823),
.B2(n_859),
.Y(n_989)
);

AO32x2_ASAP7_75t_L g990 ( 
.A1(n_877),
.A2(n_754),
.A3(n_716),
.B1(n_715),
.B2(n_693),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_776),
.B(n_177),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_817),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_870),
.B(n_688),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_839),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_762),
.A2(n_716),
.B1(n_693),
.B2(n_578),
.Y(n_995)
);

AOI21x1_ASAP7_75t_L g996 ( 
.A1(n_924),
.A2(n_503),
.B(n_447),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_842),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_857),
.A2(n_503),
.B1(n_447),
.B2(n_580),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_784),
.A2(n_496),
.B(n_498),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_777),
.A2(n_496),
.B(n_498),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_831),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_857),
.A2(n_537),
.B1(n_465),
.B2(n_580),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_774),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_915),
.B(n_465),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_777),
.A2(n_496),
.B(n_498),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_777),
.A2(n_496),
.B(n_498),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_840),
.B(n_498),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_837),
.A2(n_517),
.B(n_498),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_764),
.B(n_539),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_844),
.A2(n_517),
.B(n_528),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_919),
.B(n_466),
.Y(n_1011)
);

INVx4_ASAP7_75t_L g1012 ( 
.A(n_764),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_791),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_859),
.A2(n_541),
.B1(n_485),
.B2(n_576),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_891),
.B(n_177),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_770),
.Y(n_1016)
);

BUFx12f_ASAP7_75t_L g1017 ( 
.A(n_819),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_831),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_SL g1019 ( 
.A1(n_835),
.A2(n_537),
.B(n_466),
.C(n_576),
.Y(n_1019)
);

OR2x6_ASAP7_75t_L g1020 ( 
.A(n_769),
.B(n_517),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_847),
.A2(n_517),
.B(n_528),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_921),
.B(n_866),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_868),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_878),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_881),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_792),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_875),
.B(n_482),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_826),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_902),
.A2(n_906),
.B1(n_871),
.B2(n_832),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_894),
.Y(n_1030)
);

OA21x2_ASAP7_75t_L g1031 ( 
.A1(n_895),
.A2(n_545),
.B(n_482),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_861),
.A2(n_588),
.B1(n_539),
.B2(n_571),
.Y(n_1032)
);

NAND3xp33_ASAP7_75t_L g1033 ( 
.A(n_761),
.B(n_432),
.C(n_387),
.Y(n_1033)
);

INVx5_ASAP7_75t_L g1034 ( 
.A(n_843),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_910),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_845),
.B(n_517),
.Y(n_1036)
);

AOI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_862),
.A2(n_248),
.B1(n_177),
.B2(n_571),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_858),
.A2(n_528),
.B(n_583),
.Y(n_1038)
);

AOI21xp33_ASAP7_75t_L g1039 ( 
.A1(n_925),
.A2(n_531),
.B(n_485),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_780),
.B(n_528),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_851),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_888),
.B(n_495),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_872),
.A2(n_548),
.B(n_583),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_889),
.B(n_495),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_898),
.B(n_531),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_773),
.A2(n_583),
.B(n_548),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_836),
.A2(n_533),
.B1(n_541),
.B2(n_542),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_862),
.A2(n_533),
.B1(n_542),
.B2(n_545),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_879),
.A2(n_432),
.B(n_407),
.C(n_415),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_869),
.A2(n_588),
.B1(n_571),
.B2(n_550),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_797),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_773),
.A2(n_548),
.B(n_583),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_780),
.A2(n_588),
.B(n_550),
.C(n_539),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_935),
.Y(n_1054)
);

INVx4_ASAP7_75t_L g1055 ( 
.A(n_769),
.Y(n_1055)
);

AO32x2_ASAP7_75t_L g1056 ( 
.A1(n_933),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_1056)
);

NOR2xp67_ASAP7_75t_L g1057 ( 
.A(n_785),
.B(n_73),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_826),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_862),
.A2(n_892),
.B1(n_821),
.B2(n_810),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_826),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_908),
.B(n_561),
.Y(n_1061)
);

INVx3_ASAP7_75t_SL g1062 ( 
.A(n_869),
.Y(n_1062)
);

CKINVDCx16_ASAP7_75t_R g1063 ( 
.A(n_880),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_920),
.B(n_561),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_934),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_796),
.A2(n_800),
.B(n_805),
.C(n_890),
.Y(n_1066)
);

AOI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_781),
.A2(n_550),
.B1(n_568),
.B2(n_506),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_853),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_810),
.A2(n_548),
.B(n_583),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_782),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_768),
.A2(n_548),
.B(n_398),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_874),
.B(n_568),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_920),
.B(n_431),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_821),
.A2(n_431),
.B1(n_426),
.B2(n_394),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_928),
.B(n_1),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_855),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_SL g1077 ( 
.A1(n_765),
.A2(n_426),
.B(n_419),
.C(n_415),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_935),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_883),
.A2(n_419),
.B(n_407),
.C(n_394),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_901),
.A2(n_421),
.B(n_398),
.C(n_248),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_856),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_1071),
.A2(n_820),
.B(n_768),
.Y(n_1082)
);

OR2x6_ASAP7_75t_L g1083 ( 
.A(n_970),
.B(n_856),
.Y(n_1083)
);

OR2x2_ASAP7_75t_L g1084 ( 
.A(n_972),
.B(n_756),
.Y(n_1084)
);

AND3x4_ASAP7_75t_L g1085 ( 
.A(n_940),
.B(n_756),
.C(n_793),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_SL g1086 ( 
.A(n_1034),
.B(n_864),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1068),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_974),
.A2(n_864),
.B(n_833),
.Y(n_1088)
);

INVx6_ASAP7_75t_L g1089 ( 
.A(n_1054),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_1063),
.B(n_936),
.Y(n_1090)
);

AO21x2_ASAP7_75t_L g1091 ( 
.A1(n_1019),
.A2(n_895),
.B(n_778),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_946),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_996),
.A2(n_960),
.B(n_969),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_989),
.B(n_786),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_989),
.B(n_787),
.Y(n_1095)
);

OR2x6_ASAP7_75t_L g1096 ( 
.A(n_970),
.B(n_856),
.Y(n_1096)
);

AO31x2_ASAP7_75t_L g1097 ( 
.A1(n_1080),
.A2(n_778),
.A3(n_846),
.B(n_913),
.Y(n_1097)
);

AOI21xp33_ASAP7_75t_L g1098 ( 
.A1(n_991),
.A2(n_846),
.B(n_887),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_965),
.B(n_787),
.Y(n_1099)
);

AO31x2_ASAP7_75t_L g1100 ( 
.A1(n_944),
.A2(n_913),
.A3(n_827),
.B(n_828),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1015),
.B(n_884),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_1029),
.A2(n_812),
.B(n_876),
.C(n_865),
.Y(n_1102)
);

AO31x2_ASAP7_75t_L g1103 ( 
.A1(n_955),
.A2(n_827),
.A3(n_828),
.B(n_886),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_945),
.B(n_876),
.Y(n_1104)
);

O2A1O1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_1029),
.A2(n_790),
.B(n_804),
.C(n_825),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_976),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_948),
.A2(n_959),
.B(n_986),
.C(n_977),
.Y(n_1107)
);

OA21x2_ASAP7_75t_L g1108 ( 
.A1(n_1039),
.A2(n_790),
.B(n_804),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_1054),
.B(n_864),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_1016),
.Y(n_1110)
);

NOR2x1_ASAP7_75t_SL g1111 ( 
.A(n_1034),
.B(n_1020),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_982),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_1054),
.B(n_833),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_947),
.Y(n_1114)
);

AO31x2_ASAP7_75t_L g1115 ( 
.A1(n_955),
.A2(n_886),
.A3(n_854),
.B(n_860),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1059),
.A2(n_912),
.B1(n_860),
.B2(n_873),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1008),
.A2(n_912),
.B(n_854),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_951),
.B(n_803),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_985),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_943),
.B(n_933),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1010),
.A2(n_848),
.B(n_852),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_1062),
.B(n_929),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_982),
.Y(n_1123)
);

AOI221x1_ASAP7_75t_L g1124 ( 
.A1(n_1059),
.A2(n_917),
.B1(n_893),
.B2(n_873),
.C(n_938),
.Y(n_1124)
);

NAND3xp33_ASAP7_75t_L g1125 ( 
.A(n_979),
.B(n_911),
.C(n_808),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_1075),
.A2(n_900),
.B(n_903),
.C(n_824),
.Y(n_1126)
);

INVx4_ASAP7_75t_L g1127 ( 
.A(n_980),
.Y(n_1127)
);

AO21x2_ASAP7_75t_L g1128 ( 
.A1(n_1039),
.A2(n_829),
.B(n_896),
.Y(n_1128)
);

NAND2x1p5_ASAP7_75t_L g1129 ( 
.A(n_1034),
.B(n_916),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1021),
.A2(n_932),
.B(n_841),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1003),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_961),
.B(n_803),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1066),
.A2(n_802),
.B(n_867),
.C(n_937),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_983),
.A2(n_838),
.B1(n_841),
.B2(n_909),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1013),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_956),
.A2(n_932),
.B(n_838),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_1051),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_964),
.B(n_1007),
.Y(n_1138)
);

AOI31xp67_ASAP7_75t_L g1139 ( 
.A1(n_1032),
.A2(n_926),
.A3(n_803),
.B(n_885),
.Y(n_1139)
);

INVxp67_ASAP7_75t_SL g1140 ( 
.A(n_980),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_950),
.B(n_803),
.Y(n_1141)
);

AO31x2_ASAP7_75t_L g1142 ( 
.A1(n_1053),
.A2(n_917),
.A3(n_931),
.B(n_918),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1072),
.A2(n_926),
.B(n_918),
.C(n_916),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_939),
.A2(n_918),
.B(n_916),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_994),
.B(n_931),
.Y(n_1145)
);

NAND3x1_ASAP7_75t_L g1146 ( 
.A(n_1026),
.B(n_2),
.C(n_6),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1041),
.Y(n_1147)
);

NAND2x1_ASAP7_75t_L g1148 ( 
.A(n_980),
.B(n_843),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_966),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_968),
.A2(n_916),
.B(n_917),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_954),
.B(n_931),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1076),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_971),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_950),
.B(n_843),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_1078),
.Y(n_1155)
);

O2A1O1Ixp5_ASAP7_75t_SL g1156 ( 
.A1(n_1074),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_984),
.A2(n_421),
.B(n_147),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_1028),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_942),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_949),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_993),
.B(n_1001),
.Y(n_1161)
);

AO31x2_ASAP7_75t_L g1162 ( 
.A1(n_1048),
.A2(n_421),
.A3(n_10),
.B(n_11),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1078),
.B(n_421),
.Y(n_1163)
);

AOI21x1_ASAP7_75t_L g1164 ( 
.A1(n_999),
.A2(n_421),
.B(n_145),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_1058),
.Y(n_1165)
);

AOI21x1_ASAP7_75t_SL g1166 ( 
.A1(n_987),
.A2(n_8),
.B(n_11),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1078),
.B(n_421),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_SL g1168 ( 
.A(n_1012),
.B(n_13),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1004),
.B(n_421),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_958),
.A2(n_137),
.B(n_132),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1060),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1036),
.A2(n_20),
.B(n_21),
.C(n_23),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_995),
.A2(n_130),
.B(n_126),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_940),
.B(n_123),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_995),
.A2(n_119),
.B(n_112),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1001),
.B(n_24),
.Y(n_1176)
);

AOI21x1_ASAP7_75t_SL g1177 ( 
.A1(n_1073),
.A2(n_1011),
.B(n_1042),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_957),
.B(n_26),
.Y(n_1178)
);

OA22x2_ASAP7_75t_L g1179 ( 
.A1(n_1035),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1033),
.A2(n_32),
.B(n_33),
.C(n_36),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_998),
.A2(n_55),
.B(n_95),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_SL g1182 ( 
.A1(n_1020),
.A2(n_110),
.B(n_93),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_998),
.A2(n_87),
.B(n_81),
.Y(n_1183)
);

AOI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1002),
.A2(n_58),
.B(n_38),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_SL g1185 ( 
.A1(n_1048),
.A2(n_33),
.B(n_39),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1002),
.A2(n_40),
.B(n_41),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1014),
.A2(n_40),
.B(n_42),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1033),
.A2(n_1018),
.B(n_1037),
.C(n_1040),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1000),
.A2(n_1005),
.B(n_1006),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_975),
.Y(n_1190)
);

OR2x2_ASAP7_75t_L g1191 ( 
.A(n_1018),
.B(n_1030),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_952),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_SL g1193 ( 
.A1(n_1020),
.A2(n_1012),
.B(n_1055),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1027),
.B(n_1024),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1014),
.A2(n_1038),
.B(n_1046),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1064),
.A2(n_1061),
.B(n_1044),
.Y(n_1196)
);

AOI21xp33_ASAP7_75t_L g1197 ( 
.A1(n_1047),
.A2(n_1074),
.B(n_1049),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1052),
.A2(n_1069),
.B(n_1043),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_978),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1045),
.A2(n_981),
.B(n_1079),
.Y(n_1200)
);

OA21x2_ASAP7_75t_L g1201 ( 
.A1(n_1067),
.A2(n_1047),
.B(n_1050),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_952),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_992),
.Y(n_1203)
);

INVx4_ASAP7_75t_L g1204 ( 
.A(n_1055),
.Y(n_1204)
);

OR2x6_ASAP7_75t_L g1205 ( 
.A(n_970),
.B(n_952),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_997),
.A2(n_1025),
.B1(n_1023),
.B2(n_1065),
.Y(n_1206)
);

OAI22x1_ASAP7_75t_L g1207 ( 
.A1(n_1070),
.A2(n_962),
.B1(n_973),
.B2(n_1056),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1031),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_981),
.A2(n_1031),
.B(n_1009),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_981),
.A2(n_1009),
.B(n_1077),
.Y(n_1210)
);

AO21x2_ASAP7_75t_L g1211 ( 
.A1(n_1057),
.A2(n_990),
.B(n_1056),
.Y(n_1211)
);

O2A1O1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_953),
.A2(n_963),
.B(n_941),
.C(n_990),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_953),
.A2(n_963),
.B(n_1081),
.Y(n_1213)
);

AO22x2_ASAP7_75t_L g1214 ( 
.A1(n_1056),
.A2(n_990),
.B1(n_941),
.B2(n_1017),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1081),
.B(n_967),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1071),
.A2(n_996),
.B(n_960),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_972),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_980),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_946),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1022),
.B(n_610),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_SL g1221 ( 
.A1(n_991),
.A2(n_818),
.B(n_861),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_946),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1071),
.A2(n_996),
.B(n_960),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1148),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1119),
.Y(n_1225)
);

AO31x2_ASAP7_75t_L g1226 ( 
.A1(n_1124),
.A2(n_1207),
.A3(n_1208),
.B(n_1116),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1135),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1107),
.A2(n_1183),
.B(n_1220),
.C(n_1221),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_1100),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1147),
.Y(n_1230)
);

BUFx4f_ASAP7_75t_L g1231 ( 
.A(n_1085),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1152),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1092),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1106),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1221),
.A2(n_1200),
.B(n_1138),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1131),
.Y(n_1236)
);

BUFx8_ASAP7_75t_L g1237 ( 
.A(n_1155),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1123),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_SL g1239 ( 
.A1(n_1212),
.A2(n_1185),
.B(n_1102),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1104),
.B(n_1099),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1216),
.A2(n_1223),
.B(n_1082),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1198),
.A2(n_1093),
.B(n_1189),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_SL g1243 ( 
.A1(n_1171),
.A2(n_1122),
.B1(n_1149),
.B2(n_1165),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_1083),
.B(n_1096),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1179),
.A2(n_1098),
.B1(n_1178),
.B2(n_1197),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1120),
.A2(n_1217),
.B1(n_1151),
.B2(n_1165),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1219),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1099),
.B(n_1161),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1088),
.A2(n_1130),
.B(n_1086),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1101),
.A2(n_1090),
.B1(n_1174),
.B2(n_1168),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1100),
.Y(n_1251)
);

OAI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1168),
.A2(n_1183),
.B1(n_1094),
.B2(n_1118),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1217),
.B(n_1084),
.Y(n_1253)
);

AO21x2_ASAP7_75t_L g1254 ( 
.A1(n_1209),
.A2(n_1144),
.B(n_1195),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1164),
.A2(n_1170),
.B(n_1150),
.Y(n_1255)
);

OAI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1098),
.A2(n_1125),
.B(n_1188),
.Y(n_1256)
);

O2A1O1Ixp33_ASAP7_75t_SL g1257 ( 
.A1(n_1180),
.A2(n_1172),
.B(n_1197),
.C(n_1126),
.Y(n_1257)
);

OR2x6_ASAP7_75t_L g1258 ( 
.A(n_1193),
.B(n_1210),
.Y(n_1258)
);

AO21x2_ASAP7_75t_L g1259 ( 
.A1(n_1094),
.A2(n_1095),
.B(n_1143),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1155),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1153),
.Y(n_1261)
);

AOI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1121),
.A2(n_1116),
.B(n_1095),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1222),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1157),
.A2(n_1181),
.B(n_1177),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1086),
.A2(n_1196),
.B(n_1108),
.Y(n_1265)
);

INVxp33_ASAP7_75t_L g1266 ( 
.A(n_1114),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1173),
.A2(n_1175),
.B(n_1169),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1169),
.A2(n_1184),
.B(n_1141),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1214),
.A2(n_1125),
.B1(n_1211),
.B2(n_1087),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1100),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_SL g1271 ( 
.A1(n_1111),
.A2(n_1105),
.B(n_1141),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1214),
.A2(n_1211),
.B1(n_1160),
.B2(n_1199),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1103),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1186),
.A2(n_1187),
.B(n_1132),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1203),
.Y(n_1275)
);

A2O1A1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1133),
.A2(n_1174),
.B(n_1134),
.C(n_1194),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1166),
.A2(n_1134),
.B(n_1154),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1154),
.A2(n_1201),
.B(n_1108),
.Y(n_1278)
);

OR2x2_ASAP7_75t_L g1279 ( 
.A(n_1137),
.B(n_1158),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1110),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1127),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1129),
.A2(n_1213),
.B(n_1206),
.Y(n_1282)
);

AO31x2_ASAP7_75t_L g1283 ( 
.A1(n_1139),
.A2(n_1206),
.A3(n_1115),
.B(n_1176),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1156),
.A2(n_1109),
.B(n_1113),
.Y(n_1284)
);

AO31x2_ASAP7_75t_L g1285 ( 
.A1(n_1115),
.A2(n_1091),
.A3(n_1103),
.B(n_1097),
.Y(n_1285)
);

A2O1A1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1159),
.A2(n_1190),
.B(n_1191),
.C(n_1145),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1146),
.A2(n_1167),
.B(n_1163),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1202),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1083),
.A2(n_1096),
.B1(n_1205),
.B2(n_1089),
.Y(n_1289)
);

AOI21xp33_ASAP7_75t_L g1290 ( 
.A1(n_1128),
.A2(n_1091),
.B(n_1205),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1202),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1182),
.A2(n_1218),
.B(n_1097),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1112),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1097),
.Y(n_1294)
);

OR2x6_ASAP7_75t_L g1295 ( 
.A(n_1083),
.B(n_1096),
.Y(n_1295)
);

HB1xp67_ASAP7_75t_L g1296 ( 
.A(n_1103),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_SL g1297 ( 
.A(n_1204),
.B(n_1215),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1192),
.B(n_1205),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1215),
.A2(n_1140),
.B(n_1218),
.C(n_1128),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1115),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1162),
.Y(n_1301)
);

O2A1O1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1162),
.A2(n_1089),
.B(n_1142),
.C(n_1204),
.Y(n_1302)
);

AOI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1142),
.A2(n_481),
.B1(n_311),
.B2(n_338),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1119),
.Y(n_1304)
);

OA21x2_ASAP7_75t_L g1305 ( 
.A1(n_1124),
.A2(n_1195),
.B(n_1216),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1082),
.A2(n_1216),
.B(n_1223),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1220),
.B(n_605),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1119),
.Y(n_1308)
);

OA21x2_ASAP7_75t_L g1309 ( 
.A1(n_1124),
.A2(n_1195),
.B(n_1216),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1208),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1082),
.A2(n_1216),
.B(n_1223),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1119),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1153),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1119),
.Y(n_1314)
);

AO21x2_ASAP7_75t_L g1315 ( 
.A1(n_1136),
.A2(n_1130),
.B(n_1209),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1148),
.Y(n_1316)
);

AOI221xp5_ASAP7_75t_L g1317 ( 
.A1(n_1221),
.A2(n_682),
.B1(n_650),
.B2(n_649),
.C(n_547),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1119),
.Y(n_1318)
);

AOI21xp33_ASAP7_75t_L g1319 ( 
.A1(n_1221),
.A2(n_899),
.B(n_650),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1220),
.A2(n_899),
.B1(n_1085),
.B2(n_629),
.Y(n_1320)
);

NOR2x1_ASAP7_75t_L g1321 ( 
.A(n_1204),
.B(n_988),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1220),
.A2(n_899),
.B1(n_1085),
.B2(n_629),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1082),
.A2(n_1216),
.B(n_1223),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1083),
.B(n_1096),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1216),
.A2(n_1223),
.B(n_1082),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1220),
.B(n_605),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1119),
.Y(n_1327)
);

NOR2xp67_ASAP7_75t_L g1328 ( 
.A(n_1110),
.B(n_799),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1119),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1208),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1107),
.A2(n_815),
.B(n_814),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1171),
.A2(n_930),
.B1(n_899),
.B2(n_612),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1216),
.A2(n_1223),
.B(n_1082),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1119),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1107),
.A2(n_815),
.B(n_814),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1216),
.A2(n_1223),
.B(n_1082),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1101),
.B(n_1015),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1208),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1119),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1155),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1107),
.A2(n_815),
.B(n_814),
.Y(n_1341)
);

OAI221xp5_ASAP7_75t_L g1342 ( 
.A1(n_1221),
.A2(n_815),
.B1(n_814),
.B2(n_650),
.C(n_649),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1148),
.Y(n_1343)
);

AOI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1144),
.A2(n_1124),
.B(n_1117),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1119),
.Y(n_1345)
);

INVx4_ASAP7_75t_L g1346 ( 
.A(n_1155),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1083),
.B(n_1096),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1155),
.Y(n_1348)
);

OAI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1168),
.A2(n_1220),
.B1(n_514),
.B2(n_629),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1082),
.A2(n_1216),
.B(n_1223),
.Y(n_1350)
);

AO21x2_ASAP7_75t_L g1351 ( 
.A1(n_1136),
.A2(n_1130),
.B(n_1209),
.Y(n_1351)
);

AO21x2_ASAP7_75t_L g1352 ( 
.A1(n_1136),
.A2(n_1130),
.B(n_1209),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1119),
.Y(n_1353)
);

NOR2x1_ASAP7_75t_L g1354 ( 
.A(n_1321),
.B(n_1331),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1233),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1231),
.A2(n_1245),
.B1(n_1317),
.B2(n_1250),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1310),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1244),
.B(n_1324),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1265),
.A2(n_1228),
.B(n_1249),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1229),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1253),
.B(n_1279),
.Y(n_1361)
);

OA21x2_ASAP7_75t_L g1362 ( 
.A1(n_1235),
.A2(n_1311),
.B(n_1306),
.Y(n_1362)
);

OA21x2_ASAP7_75t_L g1363 ( 
.A1(n_1306),
.A2(n_1323),
.B(n_1311),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1323),
.A2(n_1350),
.B(n_1267),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1231),
.A2(n_1245),
.B1(n_1342),
.B2(n_1303),
.Y(n_1365)
);

INVxp67_ASAP7_75t_L g1366 ( 
.A(n_1261),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1229),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1233),
.Y(n_1368)
);

OA21x2_ASAP7_75t_L g1369 ( 
.A1(n_1350),
.A2(n_1242),
.B(n_1241),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1247),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1280),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1247),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1240),
.B(n_1248),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1307),
.B(n_1326),
.Y(n_1374)
);

BUFx2_ASAP7_75t_L g1375 ( 
.A(n_1313),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1298),
.B(n_1266),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1325),
.A2(n_1336),
.B(n_1333),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1244),
.B(n_1324),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1332),
.A2(n_1349),
.B1(n_1320),
.B2(n_1322),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_SL g1380 ( 
.A1(n_1276),
.A2(n_1335),
.B(n_1341),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1268),
.A2(n_1278),
.B(n_1274),
.Y(n_1381)
);

INVxp67_ASAP7_75t_L g1382 ( 
.A(n_1238),
.Y(n_1382)
);

O2A1O1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1349),
.A2(n_1257),
.B(n_1252),
.C(n_1256),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1246),
.B(n_1266),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1332),
.A2(n_1243),
.B1(n_1295),
.B2(n_1276),
.Y(n_1385)
);

O2A1O1Ixp5_ASAP7_75t_L g1386 ( 
.A1(n_1262),
.A2(n_1290),
.B(n_1287),
.C(n_1344),
.Y(n_1386)
);

A2O1A1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1286),
.A2(n_1347),
.B(n_1302),
.C(n_1277),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1275),
.B(n_1234),
.Y(n_1388)
);

O2A1O1Ixp5_ASAP7_75t_L g1389 ( 
.A1(n_1286),
.A2(n_1270),
.B(n_1294),
.C(n_1301),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1347),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1225),
.B(n_1227),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1238),
.Y(n_1392)
);

CKINVDCx20_ASAP7_75t_R g1393 ( 
.A(n_1280),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1237),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_SL g1395 ( 
.A1(n_1295),
.A2(n_1258),
.B(n_1299),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1347),
.B(n_1295),
.Y(n_1396)
);

AOI21x1_ASAP7_75t_SL g1397 ( 
.A1(n_1251),
.A2(n_1296),
.B(n_1273),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1328),
.A2(n_1289),
.B1(n_1293),
.B2(n_1269),
.Y(n_1398)
);

O2A1O1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1257),
.A2(n_1239),
.B(n_1271),
.C(n_1263),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1230),
.B(n_1353),
.Y(n_1400)
);

O2A1O1Ixp5_ASAP7_75t_L g1401 ( 
.A1(n_1300),
.A2(n_1224),
.B(n_1316),
.C(n_1343),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1275),
.B(n_1236),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1293),
.A2(n_1269),
.B1(n_1327),
.B2(n_1232),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_SL g1404 ( 
.A1(n_1258),
.A2(n_1259),
.B(n_1346),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1304),
.B(n_1318),
.Y(n_1405)
);

O2A1O1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1308),
.A2(n_1314),
.B(n_1345),
.C(n_1339),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1226),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1312),
.A2(n_1334),
.B1(n_1329),
.B2(n_1272),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1330),
.Y(n_1409)
);

INVxp67_ASAP7_75t_L g1410 ( 
.A(n_1288),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1278),
.A2(n_1277),
.B(n_1264),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1226),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1272),
.A2(n_1224),
.B1(n_1343),
.B2(n_1281),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1259),
.B(n_1291),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1338),
.Y(n_1415)
);

O2A1O1Ixp33_ASAP7_75t_L g1416 ( 
.A1(n_1297),
.A2(n_1281),
.B(n_1352),
.C(n_1351),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1346),
.A2(n_1260),
.B1(n_1348),
.B2(n_1340),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1338),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_SL g1419 ( 
.A1(n_1260),
.A2(n_1340),
.B(n_1348),
.Y(n_1419)
);

OAI22x1_ASAP7_75t_L g1420 ( 
.A1(n_1305),
.A2(n_1309),
.B1(n_1226),
.B2(n_1292),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1260),
.B(n_1348),
.Y(n_1421)
);

AOI211xp5_ASAP7_75t_L g1422 ( 
.A1(n_1264),
.A2(n_1284),
.B(n_1292),
.C(n_1282),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1260),
.A2(n_1340),
.B1(n_1348),
.B2(n_1305),
.Y(n_1423)
);

AND2x2_ASAP7_75t_SL g1424 ( 
.A(n_1305),
.B(n_1309),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1285),
.Y(n_1425)
);

O2A1O1Ixp5_ASAP7_75t_L g1426 ( 
.A1(n_1283),
.A2(n_1285),
.B(n_1255),
.C(n_1315),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1283),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1285),
.B(n_1254),
.Y(n_1428)
);

O2A1O1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1319),
.A2(n_1342),
.B(n_1317),
.C(n_1221),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1298),
.B(n_1337),
.Y(n_1430)
);

AOI31xp33_ASAP7_75t_L g1431 ( 
.A1(n_1317),
.A2(n_1319),
.A3(n_1245),
.B(n_1256),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1298),
.B(n_1337),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1244),
.B(n_1324),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_1280),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1231),
.A2(n_1245),
.B1(n_1085),
.B2(n_1317),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1298),
.B(n_1337),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1240),
.B(n_1248),
.Y(n_1437)
);

O2A1O1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1319),
.A2(n_1342),
.B(n_1317),
.C(n_1221),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1310),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_SL g1440 ( 
.A1(n_1228),
.A2(n_1107),
.B(n_1220),
.Y(n_1440)
);

OAI31xp33_ASAP7_75t_L g1441 ( 
.A1(n_1342),
.A2(n_1319),
.A3(n_1349),
.B(n_1221),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1317),
.A2(n_1349),
.B1(n_1322),
.B2(n_1320),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_SL g1443 ( 
.A1(n_1228),
.A2(n_1107),
.B(n_1220),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1233),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1298),
.B(n_1337),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1298),
.B(n_1337),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1298),
.B(n_1337),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1261),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_1260),
.Y(n_1449)
);

INVx3_ASAP7_75t_L g1450 ( 
.A(n_1411),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_SL g1451 ( 
.A1(n_1383),
.A2(n_1438),
.B(n_1429),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1414),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1407),
.B(n_1412),
.Y(n_1453)
);

INVx2_ASAP7_75t_SL g1454 ( 
.A(n_1388),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1396),
.Y(n_1455)
);

BUFx12f_ASAP7_75t_L g1456 ( 
.A(n_1371),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_SL g1457 ( 
.A(n_1354),
.B(n_1365),
.Y(n_1457)
);

OA21x2_ASAP7_75t_L g1458 ( 
.A1(n_1426),
.A2(n_1386),
.B(n_1359),
.Y(n_1458)
);

NOR2xp67_ASAP7_75t_L g1459 ( 
.A(n_1355),
.B(n_1368),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1373),
.B(n_1437),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1360),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1387),
.B(n_1396),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1357),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1370),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1372),
.Y(n_1465)
);

OA21x2_ASAP7_75t_L g1466 ( 
.A1(n_1389),
.A2(n_1425),
.B(n_1427),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1444),
.Y(n_1467)
);

AO21x2_ASAP7_75t_L g1468 ( 
.A1(n_1387),
.A2(n_1416),
.B(n_1380),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1407),
.B(n_1412),
.Y(n_1469)
);

INVxp67_ASAP7_75t_SL g1470 ( 
.A(n_1367),
.Y(n_1470)
);

INVxp67_ASAP7_75t_SL g1471 ( 
.A(n_1367),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1361),
.B(n_1384),
.Y(n_1472)
);

AO21x2_ASAP7_75t_L g1473 ( 
.A1(n_1431),
.A2(n_1442),
.B(n_1428),
.Y(n_1473)
);

AOI222xp33_ASAP7_75t_L g1474 ( 
.A1(n_1379),
.A2(n_1356),
.B1(n_1435),
.B2(n_1385),
.C1(n_1374),
.C2(n_1398),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1402),
.Y(n_1475)
);

NOR2x1_ASAP7_75t_L g1476 ( 
.A(n_1395),
.B(n_1404),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1415),
.B(n_1418),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1428),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1396),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1390),
.B(n_1378),
.Y(n_1480)
);

OR2x6_ASAP7_75t_L g1481 ( 
.A(n_1440),
.B(n_1443),
.Y(n_1481)
);

INVxp67_ASAP7_75t_L g1482 ( 
.A(n_1376),
.Y(n_1482)
);

OA21x2_ASAP7_75t_L g1483 ( 
.A1(n_1401),
.A2(n_1428),
.B(n_1409),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1390),
.B(n_1378),
.Y(n_1484)
);

INVxp67_ASAP7_75t_L g1485 ( 
.A(n_1375),
.Y(n_1485)
);

OR2x6_ASAP7_75t_L g1486 ( 
.A(n_1399),
.B(n_1420),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_1405),
.Y(n_1487)
);

OAI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1441),
.A2(n_1403),
.B(n_1406),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1381),
.B(n_1408),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1358),
.B(n_1378),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1363),
.A2(n_1364),
.B(n_1381),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_SL g1492 ( 
.A1(n_1394),
.A2(n_1413),
.B(n_1417),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1362),
.B(n_1358),
.Y(n_1493)
);

INVx3_ASAP7_75t_L g1494 ( 
.A(n_1381),
.Y(n_1494)
);

OAI211xp5_ASAP7_75t_L g1495 ( 
.A1(n_1366),
.A2(n_1382),
.B(n_1448),
.C(n_1392),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1423),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1410),
.Y(n_1497)
);

OA21x2_ASAP7_75t_L g1498 ( 
.A1(n_1439),
.A2(n_1400),
.B(n_1424),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1424),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1391),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1393),
.Y(n_1501)
);

INVx4_ASAP7_75t_R g1502 ( 
.A(n_1454),
.Y(n_1502)
);

OAI221xp5_ASAP7_75t_SL g1503 ( 
.A1(n_1451),
.A2(n_1430),
.B1(n_1447),
.B2(n_1446),
.C(n_1445),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1499),
.B(n_1493),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1493),
.B(n_1422),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1452),
.B(n_1436),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1493),
.B(n_1498),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1461),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1493),
.B(n_1377),
.Y(n_1509)
);

AND2x4_ASAP7_75t_L g1510 ( 
.A(n_1493),
.B(n_1433),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1498),
.B(n_1452),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1478),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1454),
.B(n_1432),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1472),
.B(n_1434),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1494),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1466),
.B(n_1450),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1466),
.B(n_1450),
.Y(n_1517)
);

AOI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1481),
.A2(n_1419),
.B(n_1369),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1489),
.B(n_1475),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1481),
.A2(n_1434),
.B1(n_1393),
.B2(n_1449),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1487),
.B(n_1421),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1463),
.Y(n_1522)
);

AO21x2_ASAP7_75t_L g1523 ( 
.A1(n_1491),
.A2(n_1397),
.B(n_1369),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1472),
.B(n_1460),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1463),
.Y(n_1525)
);

INVxp67_ASAP7_75t_L g1526 ( 
.A(n_1500),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1481),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1487),
.B(n_1449),
.Y(n_1528)
);

INVxp67_ASAP7_75t_L g1529 ( 
.A(n_1497),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1483),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1504),
.B(n_1496),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1519),
.B(n_1489),
.Y(n_1532)
);

OAI211xp5_ASAP7_75t_L g1533 ( 
.A1(n_1503),
.A2(n_1451),
.B(n_1474),
.C(n_1488),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1504),
.B(n_1496),
.Y(n_1534)
);

AOI221xp5_ASAP7_75t_L g1535 ( 
.A1(n_1529),
.A2(n_1488),
.B1(n_1457),
.B2(n_1460),
.C(n_1482),
.Y(n_1535)
);

AOI222xp33_ASAP7_75t_L g1536 ( 
.A1(n_1529),
.A2(n_1474),
.B1(n_1524),
.B2(n_1514),
.C1(n_1485),
.C2(n_1526),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1519),
.B(n_1466),
.Y(n_1537)
);

OAI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1518),
.A2(n_1481),
.B(n_1476),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1512),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_R g1540 ( 
.A(n_1520),
.B(n_1501),
.Y(n_1540)
);

NAND3xp33_ASAP7_75t_L g1541 ( 
.A(n_1503),
.B(n_1481),
.C(n_1495),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1508),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1512),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1511),
.B(n_1470),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_1521),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1522),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_SL g1547 ( 
.A1(n_1527),
.A2(n_1468),
.B1(n_1473),
.B2(n_1462),
.Y(n_1547)
);

NAND3xp33_ASAP7_75t_SL g1548 ( 
.A(n_1518),
.B(n_1495),
.C(n_1477),
.Y(n_1548)
);

NAND3xp33_ASAP7_75t_L g1549 ( 
.A(n_1527),
.B(n_1476),
.C(n_1458),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1507),
.B(n_1462),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1527),
.A2(n_1468),
.B1(n_1473),
.B2(n_1462),
.Y(n_1551)
);

NAND4xp25_ASAP7_75t_L g1552 ( 
.A(n_1528),
.B(n_1492),
.C(n_1459),
.D(n_1477),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1511),
.B(n_1471),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1527),
.A2(n_1492),
.B1(n_1486),
.B2(n_1479),
.Y(n_1554)
);

OAI221xp5_ASAP7_75t_L g1555 ( 
.A1(n_1527),
.A2(n_1486),
.B1(n_1455),
.B2(n_1479),
.C(n_1459),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1522),
.Y(n_1556)
);

INVx2_ASAP7_75t_SL g1557 ( 
.A(n_1502),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1525),
.Y(n_1558)
);

OAI31xp33_ASAP7_75t_SL g1559 ( 
.A1(n_1505),
.A2(n_1490),
.A3(n_1480),
.B(n_1484),
.Y(n_1559)
);

AOI33xp33_ASAP7_75t_L g1560 ( 
.A1(n_1505),
.A2(n_1465),
.A3(n_1467),
.B1(n_1464),
.B2(n_1469),
.B3(n_1453),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1507),
.B(n_1469),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1527),
.A2(n_1486),
.B1(n_1455),
.B2(n_1480),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1515),
.Y(n_1563)
);

INVx1_ASAP7_75t_SL g1564 ( 
.A(n_1513),
.Y(n_1564)
);

AO21x2_ASAP7_75t_L g1565 ( 
.A1(n_1523),
.A2(n_1530),
.B(n_1517),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1565),
.Y(n_1566)
);

AOI21x1_ASAP7_75t_L g1567 ( 
.A1(n_1549),
.A2(n_1530),
.B(n_1517),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1546),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1565),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1565),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1546),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1556),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_1539),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1539),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_1557),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1558),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1544),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1544),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1553),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1553),
.Y(n_1580)
);

OR2x6_ASAP7_75t_L g1581 ( 
.A(n_1538),
.B(n_1527),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1533),
.B(n_1506),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1550),
.B(n_1507),
.Y(n_1583)
);

INVxp67_ASAP7_75t_L g1584 ( 
.A(n_1548),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1532),
.Y(n_1585)
);

OA21x2_ASAP7_75t_L g1586 ( 
.A1(n_1549),
.A2(n_1509),
.B(n_1516),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1543),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1550),
.Y(n_1588)
);

INVx1_ASAP7_75t_SL g1589 ( 
.A(n_1542),
.Y(n_1589)
);

OA21x2_ASAP7_75t_L g1590 ( 
.A1(n_1551),
.A2(n_1509),
.B(n_1516),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_SL g1591 ( 
.A1(n_1541),
.A2(n_1473),
.B(n_1486),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1588),
.B(n_1531),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_R g1593 ( 
.A(n_1584),
.B(n_1456),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1588),
.B(n_1590),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1577),
.B(n_1537),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1577),
.B(n_1532),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1579),
.B(n_1564),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1575),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1588),
.B(n_1531),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1590),
.B(n_1534),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1582),
.B(n_1536),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1572),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1582),
.B(n_1545),
.Y(n_1603)
);

NAND2x1p5_ASAP7_75t_L g1604 ( 
.A(n_1574),
.B(n_1551),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1586),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1584),
.B(n_1545),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1575),
.B(n_1557),
.Y(n_1607)
);

AOI31xp33_ASAP7_75t_L g1608 ( 
.A1(n_1589),
.A2(n_1535),
.A3(n_1547),
.B(n_1554),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1572),
.Y(n_1609)
);

OAI221xp5_ASAP7_75t_L g1610 ( 
.A1(n_1591),
.A2(n_1552),
.B1(n_1559),
.B2(n_1555),
.C(n_1562),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1590),
.B(n_1534),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1572),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1575),
.B(n_1505),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1574),
.Y(n_1614)
);

INVx1_ASAP7_75t_SL g1615 ( 
.A(n_1589),
.Y(n_1615)
);

NOR2x1_ASAP7_75t_L g1616 ( 
.A(n_1575),
.B(n_1563),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1576),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1580),
.B(n_1560),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1576),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1576),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1568),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1574),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1573),
.Y(n_1623)
);

BUFx2_ASAP7_75t_L g1624 ( 
.A(n_1581),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1590),
.B(n_1561),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1568),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1583),
.B(n_1510),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1590),
.B(n_1561),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1580),
.B(n_1528),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1571),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1571),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1587),
.B(n_1506),
.Y(n_1632)
);

OAI21xp33_ASAP7_75t_L g1633 ( 
.A1(n_1601),
.A2(n_1581),
.B(n_1585),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1618),
.B(n_1585),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1602),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1609),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1615),
.B(n_1587),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1592),
.B(n_1599),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1612),
.Y(n_1639)
);

INVxp33_ASAP7_75t_L g1640 ( 
.A(n_1593),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1617),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1619),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1620),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1621),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1592),
.B(n_1583),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1596),
.B(n_1585),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1598),
.B(n_1583),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1626),
.Y(n_1648)
);

NOR2xp67_ASAP7_75t_SL g1649 ( 
.A(n_1610),
.B(n_1456),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1630),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1598),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1623),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1622),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1631),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1614),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1623),
.B(n_1603),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1599),
.B(n_1583),
.Y(n_1657)
);

INVx1_ASAP7_75t_SL g1658 ( 
.A(n_1606),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1614),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1613),
.B(n_1583),
.Y(n_1660)
);

OAI21xp33_ASAP7_75t_L g1661 ( 
.A1(n_1608),
.A2(n_1581),
.B(n_1567),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1607),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1597),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1597),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1629),
.Y(n_1665)
);

NAND2xp67_ASAP7_75t_L g1666 ( 
.A(n_1594),
.B(n_1456),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1616),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1653),
.Y(n_1668)
);

AO22x1_ASAP7_75t_L g1669 ( 
.A1(n_1640),
.A2(n_1652),
.B1(n_1658),
.B2(n_1667),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1652),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1662),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1662),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1646),
.B(n_1596),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1646),
.B(n_1595),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1643),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1640),
.B(n_1632),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1645),
.Y(n_1677)
);

CKINVDCx14_ASAP7_75t_R g1678 ( 
.A(n_1656),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1638),
.Y(n_1679)
);

NOR2x1_ASAP7_75t_L g1680 ( 
.A(n_1637),
.B(n_1607),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1643),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1634),
.B(n_1595),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_1651),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1663),
.B(n_1573),
.Y(n_1684)
);

AND2x4_ASAP7_75t_L g1685 ( 
.A(n_1651),
.B(n_1638),
.Y(n_1685)
);

AO21x2_ASAP7_75t_L g1686 ( 
.A1(n_1661),
.A2(n_1594),
.B(n_1570),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1649),
.A2(n_1581),
.B1(n_1604),
.B2(n_1624),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1647),
.B(n_1627),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1645),
.Y(n_1689)
);

AOI22x1_ASAP7_75t_L g1690 ( 
.A1(n_1667),
.A2(n_1604),
.B1(n_1624),
.B2(n_1605),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1644),
.Y(n_1691)
);

OAI21xp33_ASAP7_75t_L g1692 ( 
.A1(n_1633),
.A2(n_1604),
.B(n_1581),
.Y(n_1692)
);

OAI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1692),
.A2(n_1649),
.B1(n_1664),
.B2(n_1634),
.C(n_1665),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1685),
.B(n_1657),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1678),
.B(n_1666),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1685),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1679),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1680),
.A2(n_1659),
.B(n_1655),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1673),
.Y(n_1699)
);

OAI211xp5_ASAP7_75t_SL g1700 ( 
.A1(n_1670),
.A2(n_1648),
.B(n_1654),
.C(n_1650),
.Y(n_1700)
);

AOI221xp5_ASAP7_75t_L g1701 ( 
.A1(n_1669),
.A2(n_1605),
.B1(n_1644),
.B2(n_1600),
.C(n_1611),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1685),
.B(n_1657),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1687),
.A2(n_1581),
.B1(n_1613),
.B2(n_1647),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1683),
.A2(n_1690),
.B1(n_1581),
.B2(n_1676),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1688),
.B(n_1660),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1688),
.Y(n_1706)
);

INVxp67_ASAP7_75t_SL g1707 ( 
.A(n_1669),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1688),
.B(n_1677),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1673),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1668),
.B(n_1666),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_SL g1711 ( 
.A(n_1690),
.B(n_1647),
.Y(n_1711)
);

NOR2x1_ASAP7_75t_L g1712 ( 
.A(n_1696),
.B(n_1668),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1694),
.B(n_1702),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1699),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1694),
.B(n_1702),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1708),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1705),
.B(n_1671),
.Y(n_1717)
);

NOR2xp67_ASAP7_75t_L g1718 ( 
.A(n_1711),
.B(n_1683),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1696),
.B(n_1671),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1709),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1707),
.B(n_1672),
.Y(n_1721)
);

HB1xp67_ASAP7_75t_L g1722 ( 
.A(n_1706),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1716),
.B(n_1697),
.Y(n_1723)
);

AOI21xp33_ASAP7_75t_SL g1724 ( 
.A1(n_1721),
.A2(n_1695),
.B(n_1704),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1722),
.B(n_1684),
.Y(n_1725)
);

AOI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1714),
.A2(n_1701),
.B1(n_1700),
.B2(n_1698),
.C(n_1693),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1718),
.A2(n_1705),
.B1(n_1686),
.B2(n_1703),
.Y(n_1727)
);

AOI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1712),
.A2(n_1711),
.B(n_1686),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1720),
.B(n_1710),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1713),
.A2(n_1686),
.B1(n_1708),
.B2(n_1706),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1719),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1713),
.A2(n_1689),
.B1(n_1677),
.B2(n_1672),
.Y(n_1732)
);

OAI211xp5_ASAP7_75t_L g1733 ( 
.A1(n_1717),
.A2(n_1691),
.B(n_1681),
.C(n_1675),
.Y(n_1733)
);

AOI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1726),
.A2(n_1715),
.B1(n_1717),
.B2(n_1727),
.Y(n_1734)
);

INVxp67_ASAP7_75t_L g1735 ( 
.A(n_1731),
.Y(n_1735)
);

AOI221x1_ASAP7_75t_L g1736 ( 
.A1(n_1728),
.A2(n_1724),
.B1(n_1729),
.B2(n_1719),
.C(n_1715),
.Y(n_1736)
);

XNOR2xp5_ASAP7_75t_L g1737 ( 
.A(n_1732),
.B(n_1719),
.Y(n_1737)
);

AOI221xp5_ASAP7_75t_L g1738 ( 
.A1(n_1733),
.A2(n_1675),
.B1(n_1689),
.B2(n_1605),
.C(n_1682),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1737),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1734),
.B(n_1735),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1736),
.B(n_1723),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1738),
.B(n_1725),
.Y(n_1742)
);

NAND3xp33_ASAP7_75t_L g1743 ( 
.A(n_1736),
.B(n_1730),
.C(n_1682),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1737),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_R g1745 ( 
.A(n_1739),
.B(n_1674),
.Y(n_1745)
);

OAI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1741),
.A2(n_1743),
.B1(n_1740),
.B2(n_1744),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1742),
.A2(n_1639),
.B(n_1635),
.Y(n_1747)
);

AOI31xp33_ASAP7_75t_L g1748 ( 
.A1(n_1741),
.A2(n_1674),
.A3(n_1660),
.B(n_1641),
.Y(n_1748)
);

OAI211xp5_ASAP7_75t_L g1749 ( 
.A1(n_1741),
.A2(n_1642),
.B(n_1636),
.C(n_1586),
.Y(n_1749)
);

INVxp67_ASAP7_75t_SL g1750 ( 
.A(n_1746),
.Y(n_1750)
);

AOI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1748),
.A2(n_1600),
.B1(n_1611),
.B2(n_1570),
.C(n_1566),
.Y(n_1751)
);

OAI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1749),
.A2(n_1747),
.B1(n_1607),
.B2(n_1613),
.Y(n_1752)
);

XNOR2xp5_ASAP7_75t_L g1753 ( 
.A(n_1750),
.B(n_1745),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1753),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1754),
.B(n_1752),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1755),
.A2(n_1751),
.B(n_1570),
.Y(n_1756)
);

OAI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1756),
.A2(n_1629),
.B1(n_1625),
.B2(n_1628),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1757),
.A2(n_1569),
.B1(n_1570),
.B2(n_1566),
.Y(n_1758)
);

AOI22xp5_ASAP7_75t_SL g1759 ( 
.A1(n_1758),
.A2(n_1628),
.B1(n_1625),
.B2(n_1586),
.Y(n_1759)
);

OA21x2_ASAP7_75t_L g1760 ( 
.A1(n_1759),
.A2(n_1569),
.B(n_1566),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1759),
.B(n_1627),
.Y(n_1761)
);

INVxp67_ASAP7_75t_L g1762 ( 
.A(n_1761),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1762),
.A2(n_1760),
.B1(n_1569),
.B2(n_1566),
.Y(n_1763)
);

AOI211xp5_ASAP7_75t_L g1764 ( 
.A1(n_1763),
.A2(n_1569),
.B(n_1578),
.C(n_1540),
.Y(n_1764)
);


endmodule