module fake_ariane_2376_n_2849 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_502, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_297, n_503, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_231, n_366, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_514, n_418, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_2849);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_502;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_297;
input n_503;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_514;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;

output n_2849;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_2818;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_1837;
wire n_817;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_2461;
wire n_2207;
wire n_1706;
wire n_2702;
wire n_524;
wire n_2731;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_737;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_520;
wire n_870;
wire n_2547;
wire n_1453;
wire n_958;
wire n_945;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_557;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_559;
wire n_2233;
wire n_2663;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_533;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_612;
wire n_2739;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_2703;
wire n_696;
wire n_1442;
wire n_2620;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_762;
wire n_2791;
wire n_555;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2693;
wire n_2745;
wire n_2087;
wire n_669;
wire n_1491;
wire n_931;
wire n_2628;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_615;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_1932;
wire n_749;
wire n_1780;
wire n_2825;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_564;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_552;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_1592;
wire n_637;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_2811;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1053;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_529;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2783;
wire n_2599;
wire n_727;
wire n_590;
wire n_699;
wire n_2075;
wire n_1726;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_545;
wire n_2496;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_536;
wire n_2031;
wire n_2418;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2780;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_1402;
wire n_957;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_527;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_551;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_1373;
wire n_1081;
wire n_742;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_2119;
wire n_1719;
wire n_1540;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_2785;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_2772;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_1191;
wire n_618;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_602;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_1318;
wire n_854;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_1856;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_640;
wire n_2016;
wire n_2667;
wire n_2723;
wire n_2725;
wire n_1118;
wire n_943;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_1561;
wire n_649;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_1201;
wire n_1288;
wire n_2605;
wire n_858;
wire n_2796;
wire n_1185;
wire n_2475;
wire n_2804;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_2747;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2820;
wire n_2613;
wire n_1165;
wire n_1641;
wire n_538;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_2647;
wire n_588;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_623;
wire n_2608;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_2767;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_540;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_2828;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_1893;
wire n_932;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_2843;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_556;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_541;
wire n_2604;
wire n_1775;
wire n_788;
wire n_908;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_2630;
wire n_591;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_2395;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_898;
wire n_857;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_2583;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_1459;
wire n_840;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_614;
wire n_2775;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_2206;
wire n_635;
wire n_2784;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_2429;
wire n_684;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_723;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_2846;
wire n_1781;
wire n_709;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1983;
wire n_1273;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_1043;
wire n_1923;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_537;
wire n_1063;
wire n_991;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_1474;
wire n_937;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_1871;
wire n_803;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_548;
wire n_2336;
wire n_523;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_1308;
wire n_573;
wire n_796;
wire n_2823;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

BUFx10_ASAP7_75t_L g520 ( 
.A(n_14),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_229),
.Y(n_521)
);

CKINVDCx16_ASAP7_75t_R g522 ( 
.A(n_349),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_215),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_239),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_374),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_508),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_460),
.Y(n_527)
);

HB1xp67_ASAP7_75t_SL g528 ( 
.A(n_272),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_470),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_487),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_163),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_1),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_217),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_127),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_95),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_478),
.Y(n_536)
);

BUFx10_ASAP7_75t_L g537 ( 
.A(n_435),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_232),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_112),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_51),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_366),
.Y(n_541)
);

INVxp67_ASAP7_75t_SL g542 ( 
.A(n_90),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_324),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_308),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_328),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_19),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_169),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_375),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_493),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_32),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_231),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_183),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_418),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_263),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_18),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_61),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_342),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_425),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_311),
.Y(n_559)
);

CKINVDCx16_ASAP7_75t_R g560 ( 
.A(n_16),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_391),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_261),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_419),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_359),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_296),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_484),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_102),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_276),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_153),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_297),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_129),
.Y(n_571)
);

BUFx10_ASAP7_75t_L g572 ( 
.A(n_316),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_385),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_383),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_505),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_404),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_439),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_496),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_233),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_101),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_118),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_31),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_393),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_495),
.Y(n_584)
);

CKINVDCx14_ASAP7_75t_R g585 ( 
.A(n_75),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_384),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_238),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_344),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_364),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_372),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_218),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_428),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_302),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_377),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_517),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_283),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_349),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_205),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_473),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_33),
.Y(n_600)
);

INVx1_ASAP7_75t_SL g601 ( 
.A(n_257),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_464),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_326),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_456),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_414),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_499),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_463),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_331),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_451),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_343),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_241),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_440),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_324),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_20),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_65),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_200),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_518),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_162),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_191),
.Y(n_619)
);

BUFx5_ASAP7_75t_L g620 ( 
.A(n_152),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_480),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_406),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_396),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_431),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_420),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_475),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_256),
.Y(n_627)
);

BUFx10_ASAP7_75t_L g628 ( 
.A(n_119),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_483),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_442),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_56),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_179),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_386),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_157),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_416),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_126),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_502),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_135),
.Y(n_638)
);

INVx1_ASAP7_75t_SL g639 ( 
.A(n_507),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_78),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_330),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_491),
.Y(n_642)
);

CKINVDCx14_ASAP7_75t_R g643 ( 
.A(n_389),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_411),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_252),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_312),
.Y(n_646)
);

CKINVDCx16_ASAP7_75t_R g647 ( 
.A(n_271),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_54),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_246),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_397),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_116),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_202),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_226),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_231),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_270),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_187),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_466),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_271),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_106),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_492),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_207),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_494),
.Y(n_662)
);

BUFx10_ASAP7_75t_L g663 ( 
.A(n_58),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_285),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_145),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_287),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_122),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_405),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_89),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_413),
.Y(n_670)
);

BUFx5_ASAP7_75t_L g671 ( 
.A(n_253),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_253),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_196),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_376),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_408),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_387),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_403),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_258),
.Y(n_678)
);

CKINVDCx16_ASAP7_75t_R g679 ( 
.A(n_327),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_42),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_292),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_497),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_373),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_415),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_37),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_407),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_26),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_519),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_102),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_343),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_432),
.Y(n_691)
);

CKINVDCx14_ASAP7_75t_R g692 ( 
.A(n_122),
.Y(n_692)
);

BUFx5_ASAP7_75t_L g693 ( 
.A(n_433),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_210),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_516),
.Y(n_695)
);

BUFx10_ASAP7_75t_L g696 ( 
.A(n_305),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_230),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_203),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_121),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_14),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_474),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_322),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_513),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_436),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_370),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_208),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_509),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_424),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_237),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_200),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_143),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_395),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_500),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_421),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_39),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_217),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_449),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_335),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_29),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_211),
.Y(n_720)
);

CKINVDCx16_ASAP7_75t_R g721 ( 
.A(n_514),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_257),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_329),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_251),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_290),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_180),
.Y(n_726)
);

BUFx8_ASAP7_75t_SL g727 ( 
.A(n_114),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_168),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_126),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_201),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_104),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_363),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_319),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_444),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_380),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_454),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_379),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_141),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_186),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_378),
.Y(n_740)
);

BUFx2_ASAP7_75t_SL g741 ( 
.A(n_133),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_169),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_286),
.Y(n_743)
);

HB1xp67_ASAP7_75t_SL g744 ( 
.A(n_180),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_237),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_388),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_127),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_13),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_320),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_323),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_117),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_95),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_351),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_422),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_489),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_74),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_441),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_400),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_266),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_450),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_218),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_230),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_427),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_163),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_468),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_281),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_178),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_261),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_345),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_252),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_66),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_17),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_114),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_334),
.Y(n_774)
);

BUFx2_ASAP7_75t_SL g775 ( 
.A(n_430),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_448),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_34),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_515),
.Y(n_778)
);

BUFx2_ASAP7_75t_L g779 ( 
.A(n_212),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_486),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_381),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_128),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_73),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_477),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_394),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_447),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_115),
.Y(n_787)
);

BUFx10_ASAP7_75t_L g788 ( 
.A(n_246),
.Y(n_788)
);

CKINVDCx16_ASAP7_75t_R g789 ( 
.A(n_83),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_345),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_333),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_312),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_193),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_238),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_15),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_294),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_134),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_152),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_410),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_138),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_462),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_123),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_328),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_382),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_255),
.Y(n_805)
);

BUFx10_ASAP7_75t_L g806 ( 
.A(n_124),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_205),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_50),
.Y(n_808)
);

CKINVDCx16_ASAP7_75t_R g809 ( 
.A(n_251),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_401),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_282),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_390),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_121),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_453),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_248),
.Y(n_815)
);

CKINVDCx16_ASAP7_75t_R g816 ( 
.A(n_101),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_501),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_287),
.Y(n_818)
);

CKINVDCx20_ASAP7_75t_R g819 ( 
.A(n_267),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_334),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_503),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_308),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_465),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_361),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_455),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_319),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_467),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_112),
.Y(n_828)
);

BUFx2_ASAP7_75t_L g829 ( 
.A(n_144),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_279),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_336),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_457),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_438),
.Y(n_833)
);

BUFx5_ASAP7_75t_L g834 ( 
.A(n_320),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_471),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_307),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_183),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_459),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_512),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_235),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_476),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_48),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_443),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_458),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_197),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_446),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_71),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_248),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_452),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_194),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_244),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_11),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_402),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_42),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_323),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_219),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_35),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_429),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_294),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_423),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_233),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_62),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_511),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_232),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_269),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_105),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_196),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_365),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_322),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_12),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_479),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_398),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_5),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_288),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_333),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_437),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_417),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_70),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_124),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_207),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_188),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_469),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_58),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_243),
.Y(n_884)
);

BUFx10_ASAP7_75t_L g885 ( 
.A(n_249),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_187),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_116),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_138),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_434),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_461),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_179),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_12),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_202),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_445),
.Y(n_894)
);

INVx4_ASAP7_75t_R g895 ( 
.A(n_182),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_148),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_262),
.Y(n_897)
);

CKINVDCx20_ASAP7_75t_R g898 ( 
.A(n_426),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_276),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_113),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_318),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_360),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_306),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_219),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_250),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_412),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_103),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_361),
.Y(n_908)
);

INVx4_ASAP7_75t_R g909 ( 
.A(n_254),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_409),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_83),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_167),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_35),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_85),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_297),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_392),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_342),
.Y(n_917)
);

CKINVDCx14_ASAP7_75t_R g918 ( 
.A(n_488),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_175),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_485),
.Y(n_920)
);

BUFx10_ASAP7_75t_L g921 ( 
.A(n_249),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_109),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_216),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_130),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_270),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_371),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_49),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_67),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_131),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_125),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_490),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_472),
.Y(n_932)
);

INVx1_ASAP7_75t_SL g933 ( 
.A(n_498),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_94),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_177),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_482),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_296),
.Y(n_937)
);

INVx1_ASAP7_75t_SL g938 ( 
.A(n_265),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_254),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_481),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_115),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_504),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_111),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_245),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_92),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_399),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_70),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_225),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_132),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_506),
.Y(n_950)
);

INVx1_ASAP7_75t_SL g951 ( 
.A(n_172),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_134),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_213),
.Y(n_953)
);

BUFx10_ASAP7_75t_L g954 ( 
.A(n_304),
.Y(n_954)
);

BUFx10_ASAP7_75t_L g955 ( 
.A(n_510),
.Y(n_955)
);

INVxp67_ASAP7_75t_SL g956 ( 
.A(n_930),
.Y(n_956)
);

INVxp67_ASAP7_75t_SL g957 ( 
.A(n_930),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_930),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_585),
.Y(n_959)
);

CKINVDCx16_ASAP7_75t_R g960 ( 
.A(n_692),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_673),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_610),
.Y(n_962)
);

INVxp67_ASAP7_75t_SL g963 ( 
.A(n_673),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_535),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_620),
.Y(n_965)
);

CKINVDCx20_ASAP7_75t_R g966 ( 
.A(n_587),
.Y(n_966)
);

INVxp33_ASAP7_75t_L g967 ( 
.A(n_727),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_546),
.B(n_715),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_620),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_620),
.Y(n_970)
);

CKINVDCx16_ASAP7_75t_R g971 ( 
.A(n_522),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_620),
.Y(n_972)
);

INVxp33_ASAP7_75t_L g973 ( 
.A(n_727),
.Y(n_973)
);

INVxp33_ASAP7_75t_L g974 ( 
.A(n_779),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_620),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_721),
.Y(n_976)
);

INVxp67_ASAP7_75t_SL g977 ( 
.A(n_753),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_753),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_764),
.Y(n_979)
);

CKINVDCx16_ASAP7_75t_R g980 ( 
.A(n_560),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_620),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_764),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_770),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_770),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_772),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_772),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_797),
.Y(n_987)
);

INVxp67_ASAP7_75t_SL g988 ( 
.A(n_797),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_587),
.Y(n_989)
);

INVxp67_ASAP7_75t_SL g990 ( 
.A(n_851),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_851),
.Y(n_991)
);

INVxp33_ASAP7_75t_SL g992 ( 
.A(n_609),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_875),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_875),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_904),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_573),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_904),
.Y(n_997)
);

CKINVDCx20_ASAP7_75t_R g998 ( 
.A(n_661),
.Y(n_998)
);

CKINVDCx16_ASAP7_75t_R g999 ( 
.A(n_647),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_620),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_671),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_573),
.Y(n_1002)
);

CKINVDCx16_ASAP7_75t_R g1003 ( 
.A(n_679),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_661),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_594),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_671),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_671),
.Y(n_1007)
);

CKINVDCx16_ASAP7_75t_R g1008 ( 
.A(n_789),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_671),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_829),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_671),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_594),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_671),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_671),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_700),
.Y(n_1015)
);

INVxp33_ASAP7_75t_SL g1016 ( 
.A(n_712),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_834),
.Y(n_1017)
);

CKINVDCx20_ASAP7_75t_R g1018 ( 
.A(n_700),
.Y(n_1018)
);

INVxp67_ASAP7_75t_SL g1019 ( 
.A(n_535),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_834),
.Y(n_1020)
);

INVxp67_ASAP7_75t_SL g1021 ( 
.A(n_535),
.Y(n_1021)
);

INVxp67_ASAP7_75t_L g1022 ( 
.A(n_528),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_834),
.Y(n_1023)
);

INVxp67_ASAP7_75t_SL g1024 ( 
.A(n_535),
.Y(n_1024)
);

INVxp67_ASAP7_75t_SL g1025 ( 
.A(n_555),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_606),
.Y(n_1026)
);

INVxp33_ASAP7_75t_SL g1027 ( 
.A(n_812),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_834),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_834),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_834),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_992),
.A2(n_728),
.B1(n_739),
.B2(n_716),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_965),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_965),
.Y(n_1033)
);

OA21x2_ASAP7_75t_L g1034 ( 
.A1(n_1001),
.A2(n_575),
.B(n_525),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_972),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_963),
.B(n_643),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_972),
.Y(n_1037)
);

OA21x2_ASAP7_75t_L g1038 ( 
.A1(n_1006),
.A2(n_578),
.B(n_577),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_969),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_1007),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_969),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_975),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_970),
.A2(n_592),
.B(n_586),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_970),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_1009),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_981),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_956),
.B(n_595),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_981),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_1000),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_957),
.B(n_564),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_1000),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_964),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_964),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_1011),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_1013),
.Y(n_1055)
);

INVxp33_ASAP7_75t_SL g1056 ( 
.A(n_976),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_975),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_977),
.B(n_602),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1029),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1029),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_1022),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1014),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_964),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1030),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1030),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_1017),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_971),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_960),
.B(n_537),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_988),
.B(n_607),
.Y(n_1069)
);

CKINVDCx6p67_ASAP7_75t_R g1070 ( 
.A(n_980),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1020),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_1023),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_1028),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_958),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_1019),
.B(n_564),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_992),
.A2(n_809),
.B1(n_816),
.B2(n_744),
.Y(n_1076)
);

NAND2xp33_ASAP7_75t_L g1077 ( 
.A(n_976),
.B(n_959),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_1016),
.A2(n_794),
.B1(n_830),
.B2(n_739),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_1021),
.A2(n_642),
.B(n_623),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_961),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1024),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1025),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_1016),
.A2(n_728),
.B1(n_794),
.B2(n_716),
.Y(n_1083)
);

INVx2_ASAP7_75t_SL g1084 ( 
.A(n_959),
.Y(n_1084)
);

INVx4_ASAP7_75t_L g1085 ( 
.A(n_978),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_979),
.A2(n_657),
.B(n_650),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_990),
.B(n_913),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_982),
.A2(n_675),
.B(n_668),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_983),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_984),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_985),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_1027),
.B(n_918),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1089),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_1031),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_1070),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1089),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_1070),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_1040),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1074),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_1031),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_R g1101 ( 
.A(n_1077),
.B(n_996),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1091),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1091),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1091),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_1067),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_R g1106 ( 
.A(n_1084),
.B(n_996),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1082),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1082),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1051),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_1056),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_1061),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_1061),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_R g1113 ( 
.A(n_1084),
.B(n_1002),
.Y(n_1113)
);

INVxp67_ASAP7_75t_L g1114 ( 
.A(n_1092),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1051),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1051),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1036),
.B(n_974),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_1083),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_1078),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_1078),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_1076),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_1090),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_1090),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_1036),
.Y(n_1124)
);

CKINVDCx16_ASAP7_75t_R g1125 ( 
.A(n_1087),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_1090),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_1090),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1044),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_1087),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_1090),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1071),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1044),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_1068),
.Y(n_1133)
);

AOI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1032),
.A2(n_701),
.B(n_677),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_1090),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_1081),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1081),
.B(n_1027),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_1050),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1040),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1048),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1048),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1087),
.A2(n_695),
.B1(n_703),
.B2(n_606),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_1087),
.B(n_999),
.Y(n_1143)
);

CKINVDCx20_ASAP7_75t_R g1144 ( 
.A(n_1058),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1041),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_R g1146 ( 
.A(n_1080),
.B(n_1002),
.Y(n_1146)
);

OAI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_1047),
.A2(n_1003),
.B1(n_1008),
.B2(n_818),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1071),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1080),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1129),
.B(n_1050),
.Y(n_1150)
);

NAND3xp33_ASAP7_75t_L g1151 ( 
.A(n_1114),
.B(n_1085),
.C(n_1012),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1117),
.B(n_1005),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1128),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1128),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1109),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1138),
.B(n_1050),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_1110),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1136),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_1136),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1109),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_1125),
.B(n_1005),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1132),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1138),
.B(n_1050),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1131),
.Y(n_1164)
);

BUFx3_ASAP7_75t_L g1165 ( 
.A(n_1105),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1143),
.B(n_1085),
.Y(n_1166)
);

AND2x6_ASAP7_75t_L g1167 ( 
.A(n_1098),
.B(n_1080),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1115),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_1098),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_1095),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_1095),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1146),
.B(n_1075),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_1098),
.Y(n_1173)
);

NAND2xp33_ASAP7_75t_SL g1174 ( 
.A(n_1106),
.B(n_695),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1111),
.B(n_1012),
.Y(n_1175)
);

AND2x6_ASAP7_75t_L g1176 ( 
.A(n_1139),
.B(n_1115),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1124),
.B(n_1085),
.Y(n_1177)
);

AND2x6_ASAP7_75t_L g1178 ( 
.A(n_1139),
.B(n_1080),
.Y(n_1178)
);

BUFx4f_ASAP7_75t_L g1179 ( 
.A(n_1107),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1116),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_1139),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_1116),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1097),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1137),
.B(n_1075),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1108),
.B(n_1075),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1112),
.B(n_1026),
.Y(n_1186)
);

BUFx4f_ASAP7_75t_L g1187 ( 
.A(n_1148),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_1145),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1118),
.A2(n_1034),
.B1(n_1038),
.B2(n_968),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1132),
.Y(n_1190)
);

NAND3x1_ASAP7_75t_L g1191 ( 
.A(n_1142),
.B(n_968),
.C(n_966),
.Y(n_1191)
);

INVx1_ASAP7_75t_SL g1192 ( 
.A(n_1113),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1093),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1144),
.B(n_1026),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1140),
.Y(n_1195)
);

AO22x2_ASAP7_75t_L g1196 ( 
.A1(n_1094),
.A2(n_989),
.B1(n_998),
.B2(n_966),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1096),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_1145),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1140),
.Y(n_1199)
);

INVx4_ASAP7_75t_L g1200 ( 
.A(n_1135),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_1141),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1144),
.B(n_967),
.Y(n_1202)
);

INVx5_ASAP7_75t_L g1203 ( 
.A(n_1141),
.Y(n_1203)
);

CKINVDCx16_ASAP7_75t_R g1204 ( 
.A(n_1101),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1099),
.B(n_1040),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_1149),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1102),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1124),
.B(n_1069),
.Y(n_1208)
);

AO22x2_ASAP7_75t_L g1209 ( 
.A1(n_1094),
.A2(n_998),
.B1(n_1004),
.B2(n_989),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1121),
.B(n_973),
.Y(n_1210)
);

OAI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1118),
.A2(n_819),
.B1(n_830),
.B2(n_818),
.Y(n_1211)
);

INVxp67_ASAP7_75t_SL g1212 ( 
.A(n_1103),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1104),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1147),
.B(n_1085),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1133),
.B(n_1045),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1097),
.Y(n_1216)
);

AND2x6_ASAP7_75t_L g1217 ( 
.A(n_1134),
.B(n_574),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1135),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1119),
.B(n_1010),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1133),
.B(n_986),
.Y(n_1220)
);

INVx1_ASAP7_75t_SL g1221 ( 
.A(n_1100),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1122),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1123),
.B(n_1045),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1126),
.Y(n_1224)
);

INVx5_ASAP7_75t_L g1225 ( 
.A(n_1127),
.Y(n_1225)
);

OR2x6_ASAP7_75t_L g1226 ( 
.A(n_1120),
.B(n_741),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1165),
.B(n_962),
.Y(n_1227)
);

INVxp67_ASAP7_75t_L g1228 ( 
.A(n_1215),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1153),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1150),
.B(n_1100),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1153),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1201),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1184),
.B(n_1130),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1186),
.B(n_1004),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1164),
.Y(n_1235)
);

AND2x6_ASAP7_75t_L g1236 ( 
.A(n_1150),
.B(n_574),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1185),
.B(n_1045),
.Y(n_1237)
);

NAND2x1p5_ASAP7_75t_L g1238 ( 
.A(n_1171),
.B(n_1041),
.Y(n_1238)
);

AO22x2_ASAP7_75t_L g1239 ( 
.A1(n_1221),
.A2(n_1018),
.B1(n_1015),
.B2(n_837),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_1159),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1159),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1193),
.Y(n_1242)
);

NAND3xp33_ASAP7_75t_L g1243 ( 
.A(n_1194),
.B(n_1018),
.C(n_1015),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1197),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1201),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1154),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1158),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1213),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1207),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1154),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1162),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1162),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1219),
.B(n_987),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1190),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1190),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1175),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1199),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1152),
.B(n_991),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1199),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_1157),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1205),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1177),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1161),
.B(n_993),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1214),
.B(n_1055),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1155),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1160),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1195),
.Y(n_1267)
);

AO22x2_ASAP7_75t_L g1268 ( 
.A1(n_1196),
.A2(n_837),
.B1(n_934),
.B2(n_819),
.Y(n_1268)
);

NAND2x1p5_ASAP7_75t_L g1269 ( 
.A(n_1216),
.B(n_1041),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1177),
.B(n_994),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1168),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_1204),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1211),
.A2(n_833),
.B1(n_765),
.B2(n_737),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1210),
.B(n_995),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1159),
.Y(n_1275)
);

NAND2x1p5_ASAP7_75t_L g1276 ( 
.A(n_1192),
.B(n_1041),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1208),
.B(n_997),
.Y(n_1277)
);

INVx8_ASAP7_75t_L g1278 ( 
.A(n_1170),
.Y(n_1278)
);

AO22x2_ASAP7_75t_L g1279 ( 
.A1(n_1196),
.A2(n_939),
.B1(n_934),
.B2(n_521),
.Y(n_1279)
);

AO22x2_ASAP7_75t_L g1280 ( 
.A1(n_1209),
.A2(n_1191),
.B1(n_1220),
.B2(n_1172),
.Y(n_1280)
);

INVxp67_ASAP7_75t_L g1281 ( 
.A(n_1220),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1179),
.B(n_703),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1218),
.B(n_1222),
.Y(n_1283)
);

INVx4_ASAP7_75t_L g1284 ( 
.A(n_1225),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1180),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_1183),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1226),
.Y(n_1287)
);

NOR2xp67_ASAP7_75t_L g1288 ( 
.A(n_1151),
.B(n_1063),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1182),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1206),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1166),
.B(n_737),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_1202),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1156),
.B(n_939),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1206),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1166),
.Y(n_1295)
);

AO22x2_ASAP7_75t_L g1296 ( 
.A1(n_1209),
.A2(n_601),
.B1(n_689),
.B2(n_634),
.Y(n_1296)
);

INVxp67_ASAP7_75t_L g1297 ( 
.A(n_1226),
.Y(n_1297)
);

NAND3xp33_ASAP7_75t_L g1298 ( 
.A(n_1222),
.B(n_1224),
.C(n_1174),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_1187),
.Y(n_1299)
);

CKINVDCx14_ASAP7_75t_R g1300 ( 
.A(n_1225),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1212),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1163),
.B(n_765),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1225),
.B(n_780),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1173),
.Y(n_1304)
);

NAND2x1p5_ASAP7_75t_L g1305 ( 
.A(n_1187),
.B(n_1046),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1182),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1224),
.B(n_1055),
.Y(n_1307)
);

OAI221xp5_ASAP7_75t_L g1308 ( 
.A1(n_1179),
.A2(n_542),
.B1(n_774),
.B2(n_912),
.C(n_711),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_1200),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1200),
.B(n_780),
.Y(n_1310)
);

OAI221xp5_ASAP7_75t_L g1311 ( 
.A1(n_1189),
.A2(n_951),
.B1(n_945),
.B2(n_938),
.C(n_551),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1182),
.Y(n_1312)
);

AO22x2_ASAP7_75t_L g1313 ( 
.A1(n_1169),
.A2(n_913),
.B1(n_568),
.B2(n_569),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1173),
.Y(n_1314)
);

AO22x2_ASAP7_75t_L g1315 ( 
.A1(n_1181),
.A2(n_568),
.B1(n_569),
.B2(n_547),
.Y(n_1315)
);

O2A1O1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1181),
.A2(n_1033),
.B(n_1035),
.C(n_1032),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1173),
.B(n_833),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1188),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1188),
.Y(n_1319)
);

INVxp67_ASAP7_75t_L g1320 ( 
.A(n_1188),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1198),
.B(n_520),
.Y(n_1321)
);

NAND2x1p5_ASAP7_75t_L g1322 ( 
.A(n_1203),
.B(n_1046),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1198),
.Y(n_1323)
);

BUFx8_ASAP7_75t_L g1324 ( 
.A(n_1167),
.Y(n_1324)
);

NAND2xp33_ASAP7_75t_SL g1325 ( 
.A(n_1223),
.B(n_898),
.Y(n_1325)
);

AOI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1167),
.A2(n_841),
.B1(n_898),
.B2(n_889),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1198),
.B(n_841),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1264),
.A2(n_1203),
.B(n_1035),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1235),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1228),
.B(n_1167),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1242),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1233),
.A2(n_1203),
.B(n_1037),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1244),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1301),
.A2(n_936),
.B1(n_889),
.B2(n_551),
.Y(n_1334)
);

AOI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1237),
.A2(n_1043),
.B(n_1079),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1274),
.B(n_1167),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1234),
.B(n_936),
.Y(n_1337)
);

BUFx12f_ASAP7_75t_L g1338 ( 
.A(n_1260),
.Y(n_1338)
);

O2A1O1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1292),
.A2(n_524),
.B(n_540),
.C(n_534),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1262),
.B(n_1178),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1316),
.A2(n_1057),
.B(n_1042),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1326),
.B(n_1042),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1317),
.B(n_1178),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1255),
.Y(n_1344)
);

A2O1A1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1298),
.A2(n_1088),
.B(n_1086),
.C(n_1079),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1299),
.B(n_1178),
.Y(n_1346)
);

O2A1O1Ixp33_ASAP7_75t_SL g1347 ( 
.A1(n_1283),
.A2(n_1057),
.B(n_1060),
.C(n_1059),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1261),
.A2(n_1060),
.B(n_1059),
.Y(n_1348)
);

A2O1A1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1325),
.A2(n_1086),
.B(n_1088),
.C(n_1043),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1293),
.B(n_1064),
.Y(n_1350)
);

AND2x2_ASAP7_75t_SL g1351 ( 
.A(n_1273),
.B(n_547),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1295),
.B(n_1178),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1307),
.A2(n_1065),
.B(n_1064),
.Y(n_1353)
);

INVx5_ASAP7_75t_L g1354 ( 
.A(n_1278),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1270),
.B(n_1176),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1270),
.B(n_1176),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1229),
.A2(n_1065),
.B(n_1066),
.Y(n_1357)
);

INVxp67_ASAP7_75t_SL g1358 ( 
.A(n_1324),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1229),
.A2(n_1066),
.B(n_1062),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1290),
.A2(n_552),
.B1(n_556),
.B2(n_550),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1231),
.A2(n_1066),
.B(n_1062),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1303),
.B(n_553),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1231),
.A2(n_1062),
.B(n_1054),
.Y(n_1363)
);

A2O1A1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1294),
.A2(n_1054),
.B(n_1046),
.C(n_846),
.Y(n_1364)
);

O2A1O1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1308),
.A2(n_544),
.B(n_559),
.C(n_554),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1253),
.B(n_1176),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1246),
.A2(n_1054),
.B(n_1176),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1324),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1248),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1246),
.A2(n_1073),
.B(n_1072),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1321),
.B(n_1046),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1263),
.B(n_1063),
.Y(n_1372)
);

A2O1A1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1311),
.A2(n_590),
.B(n_846),
.C(n_757),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_1278),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1258),
.B(n_1063),
.Y(n_1375)
);

OAI321xp33_ASAP7_75t_L g1376 ( 
.A1(n_1243),
.A2(n_588),
.A3(n_596),
.B1(n_608),
.B2(n_597),
.C(n_571),
.Y(n_1376)
);

CKINVDCx11_ASAP7_75t_R g1377 ( 
.A(n_1272),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_SL g1378 ( 
.A(n_1303),
.B(n_553),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1250),
.A2(n_1073),
.B(n_1072),
.Y(n_1379)
);

CKINVDCx10_ASAP7_75t_R g1380 ( 
.A(n_1286),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1309),
.A2(n_552),
.B1(n_556),
.B2(n_550),
.Y(n_1381)
);

O2A1O1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1310),
.A2(n_614),
.B(n_616),
.C(n_611),
.Y(n_1382)
);

NAND3xp33_ASAP7_75t_L g1383 ( 
.A(n_1256),
.B(n_531),
.C(n_523),
.Y(n_1383)
);

INVx1_ASAP7_75t_SL g1384 ( 
.A(n_1227),
.Y(n_1384)
);

BUFx4f_ASAP7_75t_L g1385 ( 
.A(n_1230),
.Y(n_1385)
);

AO22x1_ASAP7_75t_L g1386 ( 
.A1(n_1230),
.A2(n_562),
.B1(n_565),
.B2(n_557),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1251),
.A2(n_1073),
.B(n_1072),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1252),
.A2(n_1259),
.B(n_1254),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1314),
.A2(n_1073),
.B(n_1072),
.Y(n_1389)
);

OAI321xp33_ASAP7_75t_L g1390 ( 
.A1(n_1282),
.A2(n_685),
.A3(n_653),
.B1(n_694),
.B2(n_664),
.C(n_645),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1257),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1291),
.B(n_1302),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1300),
.Y(n_1393)
);

AOI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1302),
.A2(n_1217),
.B1(n_532),
.B2(n_538),
.Y(n_1394)
);

AO22x1_ASAP7_75t_L g1395 ( 
.A1(n_1291),
.A2(n_567),
.B1(n_579),
.B2(n_570),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1314),
.A2(n_1073),
.B(n_1072),
.Y(n_1396)
);

INVx4_ASAP7_75t_L g1397 ( 
.A(n_1284),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1241),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1249),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1236),
.B(n_1063),
.Y(n_1400)
);

A2O1A1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1288),
.A2(n_757),
.B(n_590),
.C(n_714),
.Y(n_1401)
);

O2A1O1Ixp5_ASAP7_75t_SL g1402 ( 
.A1(n_1327),
.A2(n_699),
.B(n_710),
.C(n_698),
.Y(n_1402)
);

A2O1A1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1232),
.A2(n_732),
.B(n_735),
.C(n_704),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1245),
.A2(n_1217),
.B(n_1038),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1236),
.B(n_1217),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1304),
.A2(n_1038),
.B(n_1034),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1304),
.A2(n_1038),
.B(n_1034),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1236),
.B(n_1313),
.Y(n_1408)
);

INVxp67_ASAP7_75t_L g1409 ( 
.A(n_1277),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1284),
.B(n_558),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1281),
.B(n_520),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1241),
.B(n_558),
.Y(n_1412)
);

BUFx8_ASAP7_75t_L g1413 ( 
.A(n_1287),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1304),
.A2(n_1034),
.B(n_1039),
.Y(n_1414)
);

NOR2xp67_ASAP7_75t_L g1415 ( 
.A(n_1297),
.B(n_1052),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1268),
.B(n_520),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_1241),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1323),
.A2(n_1049),
.B(n_1039),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1236),
.B(n_1217),
.Y(n_1419)
);

A2O1A1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1247),
.A2(n_740),
.B(n_746),
.C(n_736),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1280),
.B(n_565),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1238),
.A2(n_724),
.B(n_726),
.C(n_719),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1337),
.B(n_1350),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1328),
.A2(n_1318),
.B(n_1315),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1344),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1334),
.B(n_1269),
.Y(n_1426)
);

NOR2x1_ASAP7_75t_L g1427 ( 
.A(n_1368),
.B(n_1240),
.Y(n_1427)
);

OR2x6_ASAP7_75t_SL g1428 ( 
.A(n_1381),
.B(n_567),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1391),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1342),
.A2(n_1276),
.B(n_1320),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1393),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1332),
.A2(n_1315),
.B(n_1322),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1329),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1336),
.A2(n_1305),
.B1(n_1280),
.B2(n_1268),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1384),
.B(n_1240),
.Y(n_1435)
);

BUFx12f_ASAP7_75t_L g1436 ( 
.A(n_1377),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1399),
.Y(n_1437)
);

A2O1A1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1365),
.A2(n_1319),
.B(n_1289),
.C(n_1312),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1409),
.B(n_1275),
.Y(n_1439)
);

BUFx2_ASAP7_75t_SL g1440 ( 
.A(n_1354),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1330),
.A2(n_1279),
.B1(n_1296),
.B2(n_1275),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1351),
.A2(n_1279),
.B1(n_1239),
.B2(n_1296),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1392),
.B(n_1275),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1343),
.A2(n_878),
.B1(n_579),
.B2(n_865),
.Y(n_1444)
);

O2A1O1Ixp33_ASAP7_75t_L g1445 ( 
.A1(n_1339),
.A2(n_1373),
.B(n_1347),
.C(n_1422),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1394),
.A2(n_947),
.B1(n_879),
.B2(n_865),
.Y(n_1446)
);

O2A1O1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1382),
.A2(n_742),
.B(n_745),
.C(n_738),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1416),
.A2(n_1239),
.B1(n_1267),
.B2(n_1266),
.Y(n_1448)
);

AOI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1335),
.A2(n_1306),
.B(n_1271),
.Y(n_1449)
);

OR2x6_ASAP7_75t_L g1450 ( 
.A(n_1340),
.B(n_1265),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1395),
.B(n_1285),
.Y(n_1451)
);

NAND2xp33_ASAP7_75t_SL g1452 ( 
.A(n_1374),
.B(n_570),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1385),
.B(n_576),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1367),
.A2(n_839),
.B(n_705),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1366),
.A2(n_947),
.B1(n_879),
.B2(n_867),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1414),
.A2(n_916),
.B(n_910),
.Y(n_1456)
);

A2O1A1Ixp33_ASAP7_75t_SL g1457 ( 
.A1(n_1353),
.A2(n_761),
.B(n_767),
.C(n_751),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1331),
.B(n_866),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1333),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1411),
.Y(n_1460)
);

O2A1O1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1420),
.A2(n_777),
.B(n_782),
.C(n_773),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1369),
.B(n_1052),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1386),
.B(n_866),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1405),
.A2(n_1419),
.B(n_1346),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1398),
.Y(n_1465)
);

A2O1A1Ixp33_ASAP7_75t_L g1466 ( 
.A1(n_1390),
.A2(n_561),
.B(n_717),
.C(n_660),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_SL g1467 ( 
.A(n_1385),
.B(n_563),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1340),
.B(n_1355),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_SL g1469 ( 
.A(n_1356),
.B(n_563),
.Y(n_1469)
);

NOR3xp33_ASAP7_75t_SL g1470 ( 
.A(n_1383),
.B(n_874),
.C(n_867),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1370),
.A2(n_916),
.B(n_910),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1398),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1388),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1375),
.Y(n_1474)
);

INVx8_ASAP7_75t_L g1475 ( 
.A(n_1354),
.Y(n_1475)
);

CKINVDCx8_ASAP7_75t_R g1476 ( 
.A(n_1380),
.Y(n_1476)
);

AO22x1_ASAP7_75t_L g1477 ( 
.A1(n_1358),
.A2(n_878),
.B1(n_900),
.B2(n_874),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1346),
.B(n_1053),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1371),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1357),
.A2(n_1049),
.B(n_1039),
.Y(n_1480)
);

AOI22x1_ASAP7_75t_L g1481 ( 
.A1(n_1341),
.A2(n_901),
.B1(n_948),
.B2(n_900),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1372),
.B(n_901),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1348),
.A2(n_1049),
.B(n_1039),
.Y(n_1483)
);

OR2x6_ASAP7_75t_L g1484 ( 
.A(n_1368),
.B(n_775),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1354),
.A2(n_1352),
.B1(n_1397),
.B2(n_1412),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1362),
.B(n_1378),
.Y(n_1486)
);

CKINVDCx20_ASAP7_75t_R g1487 ( 
.A(n_1413),
.Y(n_1487)
);

O2A1O1Ixp5_ASAP7_75t_L g1488 ( 
.A1(n_1410),
.A2(n_791),
.B(n_802),
.C(n_783),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1421),
.B(n_948),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1398),
.B(n_946),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1417),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1338),
.Y(n_1492)
);

INVx6_ASAP7_75t_L g1493 ( 
.A(n_1413),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1417),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1397),
.B(n_533),
.Y(n_1495)
);

NOR3xp33_ASAP7_75t_SL g1496 ( 
.A(n_1360),
.B(n_543),
.C(n_539),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1415),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1417),
.B(n_572),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1400),
.Y(n_1499)
);

NAND2xp33_ASAP7_75t_SL g1500 ( 
.A(n_1408),
.B(n_545),
.Y(n_1500)
);

OAI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1359),
.A2(n_763),
.B(n_754),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1361),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1403),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1379),
.A2(n_1049),
.B(n_1039),
.Y(n_1504)
);

AOI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1387),
.A2(n_1049),
.B(n_1039),
.Y(n_1505)
);

AO21x1_ASAP7_75t_L g1506 ( 
.A1(n_1404),
.A2(n_801),
.B(n_778),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1402),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1376),
.B(n_946),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_R g1509 ( 
.A(n_1401),
.B(n_576),
.Y(n_1509)
);

O2A1O1Ixp33_ASAP7_75t_SL g1510 ( 
.A1(n_1364),
.A2(n_813),
.B(n_820),
.C(n_808),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1349),
.B(n_572),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1363),
.B(n_581),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1389),
.B(n_582),
.Y(n_1513)
);

O2A1O1Ixp33_ASAP7_75t_L g1514 ( 
.A1(n_1345),
.A2(n_847),
.B(n_855),
.C(n_845),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_SL g1515 ( 
.A(n_1396),
.B(n_776),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_1418),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1406),
.Y(n_1517)
);

AOI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1407),
.A2(n_821),
.B(n_810),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1350),
.B(n_776),
.Y(n_1519)
);

BUFx2_ASAP7_75t_L g1520 ( 
.A(n_1393),
.Y(n_1520)
);

INVx1_ASAP7_75t_SL g1521 ( 
.A(n_1384),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1475),
.Y(n_1522)
);

INVx2_ASAP7_75t_SL g1523 ( 
.A(n_1493),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_L g1524 ( 
.A(n_1475),
.Y(n_1524)
);

BUFx12f_ASAP7_75t_L g1525 ( 
.A(n_1436),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_SL g1526 ( 
.A(n_1423),
.B(n_876),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1475),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1484),
.Y(n_1528)
);

CKINVDCx16_ASAP7_75t_R g1529 ( 
.A(n_1487),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1459),
.Y(n_1530)
);

BUFx12f_ASAP7_75t_L g1531 ( 
.A(n_1493),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1484),
.Y(n_1532)
);

INVx4_ASAP7_75t_L g1533 ( 
.A(n_1465),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1437),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1431),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1474),
.B(n_1053),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1435),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1449),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1433),
.Y(n_1539)
);

BUFx6f_ASAP7_75t_L g1540 ( 
.A(n_1450),
.Y(n_1540)
);

INVx2_ASAP7_75t_SL g1541 ( 
.A(n_1520),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1425),
.Y(n_1542)
);

INVx5_ASAP7_75t_SL g1543 ( 
.A(n_1484),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1465),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1519),
.A2(n_572),
.B1(n_663),
.B2(n_628),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1429),
.Y(n_1546)
);

BUFx3_ASAP7_75t_L g1547 ( 
.A(n_1443),
.Y(n_1547)
);

BUFx12f_ASAP7_75t_L g1548 ( 
.A(n_1492),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1478),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1442),
.A2(n_1448),
.B1(n_1503),
.B2(n_1511),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1439),
.Y(n_1551)
);

NAND2x1p5_ASAP7_75t_L g1552 ( 
.A(n_1494),
.B(n_717),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_1450),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1473),
.Y(n_1554)
);

INVx5_ASAP7_75t_L g1555 ( 
.A(n_1450),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1472),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1517),
.Y(n_1557)
);

INVx5_ASAP7_75t_L g1558 ( 
.A(n_1516),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1478),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1462),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1498),
.B(n_628),
.Y(n_1561)
);

BUFx6f_ASAP7_75t_L g1562 ( 
.A(n_1468),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1494),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1499),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1521),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1479),
.Y(n_1566)
);

BUFx8_ASAP7_75t_L g1567 ( 
.A(n_1476),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1491),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1451),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1521),
.Y(n_1570)
);

INVx6_ASAP7_75t_SL g1571 ( 
.A(n_1440),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1497),
.Y(n_1572)
);

INVx5_ASAP7_75t_L g1573 ( 
.A(n_1516),
.Y(n_1573)
);

INVx6_ASAP7_75t_L g1574 ( 
.A(n_1516),
.Y(n_1574)
);

INVx1_ASAP7_75t_SL g1575 ( 
.A(n_1427),
.Y(n_1575)
);

NAND2x1p5_ASAP7_75t_L g1576 ( 
.A(n_1453),
.B(n_784),
.Y(n_1576)
);

BUFx2_ASAP7_75t_SL g1577 ( 
.A(n_1467),
.Y(n_1577)
);

INVx5_ASAP7_75t_L g1578 ( 
.A(n_1507),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1460),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1502),
.Y(n_1580)
);

BUFx6f_ASAP7_75t_L g1581 ( 
.A(n_1426),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_1469),
.Y(n_1582)
);

AOI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1452),
.A2(n_663),
.B1(n_696),
.B2(n_628),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1428),
.B(n_954),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1441),
.Y(n_1585)
);

CKINVDCx16_ASAP7_75t_R g1586 ( 
.A(n_1509),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1434),
.Y(n_1587)
);

INVx2_ASAP7_75t_SL g1588 ( 
.A(n_1486),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1512),
.Y(n_1589)
);

BUFx3_ASAP7_75t_L g1590 ( 
.A(n_1485),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_1495),
.Y(n_1591)
);

INVx3_ASAP7_75t_L g1592 ( 
.A(n_1458),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1500),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1438),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1514),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1463),
.B(n_954),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1430),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1482),
.Y(n_1598)
);

BUFx2_ASAP7_75t_SL g1599 ( 
.A(n_1490),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1506),
.Y(n_1600)
);

INVx5_ASAP7_75t_L g1601 ( 
.A(n_1464),
.Y(n_1601)
);

INVx3_ASAP7_75t_SL g1602 ( 
.A(n_1515),
.Y(n_1602)
);

INVx1_ASAP7_75t_SL g1603 ( 
.A(n_1432),
.Y(n_1603)
);

INVx6_ASAP7_75t_SL g1604 ( 
.A(n_1477),
.Y(n_1604)
);

OA21x2_ASAP7_75t_L g1605 ( 
.A1(n_1538),
.A2(n_1424),
.B(n_1456),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1601),
.A2(n_1501),
.B(n_1518),
.Y(n_1606)
);

AOI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1586),
.A2(n_1508),
.B1(n_1496),
.B2(n_1446),
.Y(n_1607)
);

OAI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1538),
.A2(n_1505),
.B(n_1504),
.Y(n_1608)
);

OA21x2_ASAP7_75t_L g1609 ( 
.A1(n_1603),
.A2(n_1454),
.B(n_1471),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1554),
.Y(n_1610)
);

AOI22x1_ASAP7_75t_L g1611 ( 
.A1(n_1533),
.A2(n_1593),
.B1(n_1599),
.B2(n_1589),
.Y(n_1611)
);

OAI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1526),
.A2(n_1445),
.B(n_1466),
.Y(n_1612)
);

OAI22x1_ASAP7_75t_L g1613 ( 
.A1(n_1587),
.A2(n_1481),
.B1(n_1489),
.B2(n_1513),
.Y(n_1613)
);

OAI21x1_ASAP7_75t_L g1614 ( 
.A1(n_1580),
.A2(n_1480),
.B(n_1483),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1567),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1570),
.B(n_1535),
.Y(n_1616)
);

BUFx2_ASAP7_75t_L g1617 ( 
.A(n_1535),
.Y(n_1617)
);

OAI21x1_ASAP7_75t_L g1618 ( 
.A1(n_1580),
.A2(n_1501),
.B(n_1488),
.Y(n_1618)
);

OAI21x1_ASAP7_75t_L g1619 ( 
.A1(n_1594),
.A2(n_1461),
.B(n_1447),
.Y(n_1619)
);

OAI21x1_ASAP7_75t_L g1620 ( 
.A1(n_1557),
.A2(n_1600),
.B(n_1589),
.Y(n_1620)
);

OAI21x1_ASAP7_75t_L g1621 ( 
.A1(n_1557),
.A2(n_1455),
.B(n_1444),
.Y(n_1621)
);

AO221x2_ASAP7_75t_L g1622 ( 
.A1(n_1597),
.A2(n_923),
.B1(n_869),
.B2(n_870),
.C(n_873),
.Y(n_1622)
);

OAI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1526),
.A2(n_1470),
.B(n_1510),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1583),
.A2(n_1457),
.B(n_883),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1539),
.Y(n_1625)
);

AO21x2_ASAP7_75t_L g1626 ( 
.A1(n_1600),
.A2(n_827),
.B(n_825),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_1574),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1570),
.B(n_859),
.Y(n_1628)
);

NAND2x1_ASAP7_75t_L g1629 ( 
.A(n_1574),
.B(n_1581),
.Y(n_1629)
);

OAI21x1_ASAP7_75t_L g1630 ( 
.A1(n_1536),
.A2(n_863),
.B(n_853),
.Y(n_1630)
);

AO21x2_ASAP7_75t_L g1631 ( 
.A1(n_1569),
.A2(n_872),
.B(n_871),
.Y(n_1631)
);

BUFx2_ASAP7_75t_L g1632 ( 
.A(n_1571),
.Y(n_1632)
);

INVx4_ASAP7_75t_L g1633 ( 
.A(n_1581),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1565),
.Y(n_1634)
);

OAI21x1_ASAP7_75t_L g1635 ( 
.A1(n_1536),
.A2(n_890),
.B(n_882),
.Y(n_1635)
);

OA21x2_ASAP7_75t_L g1636 ( 
.A1(n_1603),
.A2(n_906),
.B(n_894),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1564),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1571),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1572),
.A2(n_920),
.B(n_886),
.Y(n_1639)
);

BUFx2_ASAP7_75t_SL g1640 ( 
.A(n_1523),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1565),
.B(n_884),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1601),
.B(n_784),
.Y(n_1642)
);

OA21x2_ASAP7_75t_L g1643 ( 
.A1(n_1585),
.A2(n_902),
.B(n_897),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1550),
.A2(n_1595),
.B1(n_1598),
.B2(n_1592),
.Y(n_1644)
);

OAI21x1_ASAP7_75t_L g1645 ( 
.A1(n_1564),
.A2(n_917),
.B(n_914),
.Y(n_1645)
);

AO222x2_ASAP7_75t_L g1646 ( 
.A1(n_1584),
.A2(n_806),
.B1(n_696),
.B2(n_885),
.C1(n_788),
.C2(n_663),
.Y(n_1646)
);

BUFx6f_ASAP7_75t_L g1647 ( 
.A(n_1524),
.Y(n_1647)
);

OA21x2_ASAP7_75t_L g1648 ( 
.A1(n_1530),
.A2(n_937),
.B(n_919),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1556),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1534),
.Y(n_1650)
);

OAI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1545),
.A2(n_949),
.B(n_943),
.Y(n_1651)
);

INVx2_ASAP7_75t_SL g1652 ( 
.A(n_1574),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1566),
.Y(n_1653)
);

OAI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1552),
.A2(n_648),
.B(n_618),
.Y(n_1654)
);

CKINVDCx16_ASAP7_75t_R g1655 ( 
.A(n_1529),
.Y(n_1655)
);

OAI21x1_ASAP7_75t_L g1656 ( 
.A1(n_1552),
.A2(n_648),
.B(n_618),
.Y(n_1656)
);

OAI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1592),
.A2(n_680),
.B(n_658),
.Y(n_1657)
);

NOR2xp67_ASAP7_75t_L g1658 ( 
.A(n_1601),
.B(n_0),
.Y(n_1658)
);

OAI21x1_ASAP7_75t_L g1659 ( 
.A1(n_1542),
.A2(n_680),
.B(n_658),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1546),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1578),
.Y(n_1661)
);

OAI21x1_ASAP7_75t_L g1662 ( 
.A1(n_1560),
.A2(n_756),
.B(n_697),
.Y(n_1662)
);

OAI21x1_ASAP7_75t_SL g1663 ( 
.A1(n_1541),
.A2(n_756),
.B(n_697),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1622),
.A2(n_1550),
.B1(n_1598),
.B2(n_1596),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1661),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1637),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1634),
.B(n_1581),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1625),
.Y(n_1668)
);

OAI21x1_ASAP7_75t_L g1669 ( 
.A1(n_1608),
.A2(n_1559),
.B(n_1549),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1637),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1610),
.Y(n_1671)
);

INVx3_ASAP7_75t_L g1672 ( 
.A(n_1661),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1649),
.Y(n_1673)
);

INVx3_ASAP7_75t_L g1674 ( 
.A(n_1627),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1610),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1615),
.Y(n_1676)
);

HB1xp67_ASAP7_75t_L g1677 ( 
.A(n_1617),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1650),
.Y(n_1678)
);

NOR2x1_ASAP7_75t_L g1679 ( 
.A(n_1633),
.B(n_1590),
.Y(n_1679)
);

NAND2x1p5_ASAP7_75t_L g1680 ( 
.A(n_1636),
.B(n_1601),
.Y(n_1680)
);

INVx2_ASAP7_75t_SL g1681 ( 
.A(n_1616),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1627),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_SL g1683 ( 
.A1(n_1622),
.A2(n_1590),
.B1(n_1543),
.B2(n_1593),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1653),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1620),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1620),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1660),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1660),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_1629),
.Y(n_1689)
);

AO21x2_ASAP7_75t_L g1690 ( 
.A1(n_1626),
.A2(n_1608),
.B(n_1614),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1643),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1605),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1605),
.Y(n_1693)
);

OA21x2_ASAP7_75t_L g1694 ( 
.A1(n_1614),
.A2(n_1563),
.B(n_1568),
.Y(n_1694)
);

INVx4_ASAP7_75t_SL g1695 ( 
.A(n_1642),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1643),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1643),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1652),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1605),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1662),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1636),
.Y(n_1701)
);

OAI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1607),
.A2(n_1591),
.B1(n_1604),
.B2(n_1602),
.Y(n_1702)
);

BUFx6f_ASAP7_75t_L g1703 ( 
.A(n_1647),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1636),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1662),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1659),
.Y(n_1706)
);

INVxp67_ASAP7_75t_L g1707 ( 
.A(n_1628),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1645),
.Y(n_1708)
);

NAND2x1p5_ASAP7_75t_L g1709 ( 
.A(n_1633),
.B(n_1555),
.Y(n_1709)
);

AOI21x1_ASAP7_75t_L g1710 ( 
.A1(n_1613),
.A2(n_1532),
.B(n_1528),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1659),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_1615),
.Y(n_1712)
);

NAND2xp33_ASAP7_75t_SL g1713 ( 
.A(n_1676),
.B(n_1647),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1673),
.B(n_1641),
.Y(n_1714)
);

NAND2xp33_ASAP7_75t_R g1715 ( 
.A(n_1694),
.B(n_1648),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1681),
.B(n_1655),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1681),
.B(n_1640),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1677),
.B(n_1633),
.Y(n_1718)
);

NOR2x1_ASAP7_75t_SL g1719 ( 
.A(n_1710),
.B(n_1531),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1668),
.B(n_1579),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_R g1721 ( 
.A(n_1676),
.B(n_1567),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1674),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1698),
.B(n_1652),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1668),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_R g1725 ( 
.A(n_1712),
.B(n_1525),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1666),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1666),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1670),
.Y(n_1728)
);

BUFx4f_ASAP7_75t_SL g1729 ( 
.A(n_1703),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1670),
.Y(n_1730)
);

NAND2xp33_ASAP7_75t_R g1731 ( 
.A(n_1694),
.B(n_1648),
.Y(n_1731)
);

AO31x2_ASAP7_75t_L g1732 ( 
.A1(n_1691),
.A2(n_1613),
.A3(n_1606),
.B(n_1533),
.Y(n_1732)
);

BUFx6f_ASAP7_75t_L g1733 ( 
.A(n_1703),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_SL g1734 ( 
.A1(n_1680),
.A2(n_1622),
.B1(n_1646),
.B2(n_1648),
.Y(n_1734)
);

INVx3_ASAP7_75t_L g1735 ( 
.A(n_1674),
.Y(n_1735)
);

OAI21x1_ASAP7_75t_L g1736 ( 
.A1(n_1710),
.A2(n_1611),
.B(n_1639),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1712),
.Y(n_1737)
);

CKINVDCx16_ASAP7_75t_R g1738 ( 
.A(n_1667),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1678),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1665),
.B(n_1627),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1678),
.B(n_1578),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1679),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1684),
.Y(n_1743)
);

CKINVDCx20_ASAP7_75t_R g1744 ( 
.A(n_1707),
.Y(n_1744)
);

NAND3xp33_ASAP7_75t_SL g1745 ( 
.A(n_1683),
.B(n_1644),
.C(n_1612),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1684),
.B(n_1588),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1687),
.Y(n_1747)
);

BUFx6f_ASAP7_75t_L g1748 ( 
.A(n_1703),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_L g1749 ( 
.A(n_1703),
.Y(n_1749)
);

NOR3xp33_ASAP7_75t_SL g1750 ( 
.A(n_1702),
.B(n_1623),
.C(n_593),
.Y(n_1750)
);

BUFx4f_ASAP7_75t_SL g1751 ( 
.A(n_1703),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1687),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1688),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1665),
.B(n_1632),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1665),
.B(n_1578),
.Y(n_1755)
);

CKINVDCx16_ASAP7_75t_R g1756 ( 
.A(n_1689),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1672),
.B(n_1638),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1672),
.B(n_1578),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1694),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_R g1760 ( 
.A(n_1674),
.B(n_1548),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_1689),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1672),
.B(n_1647),
.Y(n_1762)
);

O2A1O1Ixp33_ASAP7_75t_SL g1763 ( 
.A1(n_1682),
.A2(n_1646),
.B(n_880),
.C(n_907),
.Y(n_1763)
);

CKINVDCx20_ASAP7_75t_R g1764 ( 
.A(n_1689),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1688),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1671),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1754),
.B(n_1682),
.Y(n_1767)
);

INVxp67_ASAP7_75t_L g1768 ( 
.A(n_1714),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1737),
.B(n_1591),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1723),
.B(n_1682),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1718),
.B(n_1694),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1759),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1724),
.Y(n_1773)
);

AND2x4_ASAP7_75t_L g1774 ( 
.A(n_1742),
.B(n_1695),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1724),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1761),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1759),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_SL g1778 ( 
.A1(n_1734),
.A2(n_1626),
.B1(n_1631),
.B2(n_1543),
.Y(n_1778)
);

AND2x4_ASAP7_75t_L g1779 ( 
.A(n_1757),
.B(n_1695),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1720),
.B(n_1685),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1766),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1739),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1746),
.B(n_1685),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1747),
.Y(n_1784)
);

INVxp67_ASAP7_75t_L g1785 ( 
.A(n_1717),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1716),
.B(n_1686),
.Y(n_1786)
);

BUFx2_ASAP7_75t_L g1787 ( 
.A(n_1722),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1752),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1726),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1753),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1765),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1743),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1738),
.B(n_1686),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1741),
.B(n_1689),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1741),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1727),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1757),
.B(n_1690),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1740),
.B(n_1689),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1795),
.B(n_1732),
.Y(n_1799)
);

AOI21xp33_ASAP7_75t_L g1800 ( 
.A1(n_1795),
.A2(n_1731),
.B(n_1715),
.Y(n_1800)
);

AND2x6_ASAP7_75t_L g1801 ( 
.A(n_1774),
.B(n_1543),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1772),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1773),
.Y(n_1803)
);

AO21x2_ASAP7_75t_L g1804 ( 
.A1(n_1772),
.A2(n_1745),
.B(n_1763),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1771),
.B(n_1756),
.Y(n_1805)
);

OAI221xp5_ASAP7_75t_L g1806 ( 
.A1(n_1778),
.A2(n_1734),
.B1(n_1745),
.B2(n_1750),
.C(n_1731),
.Y(n_1806)
);

INVx5_ASAP7_75t_L g1807 ( 
.A(n_1774),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1777),
.Y(n_1808)
);

AOI21xp33_ASAP7_75t_L g1809 ( 
.A1(n_1777),
.A2(n_1715),
.B(n_1755),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1782),
.Y(n_1810)
);

AOI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1793),
.A2(n_1750),
.B1(n_1664),
.B2(n_1644),
.Y(n_1811)
);

OAI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1768),
.A2(n_1736),
.B(n_1744),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1792),
.Y(n_1813)
);

OAI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1773),
.A2(n_1658),
.B(n_1755),
.Y(n_1814)
);

BUFx2_ASAP7_75t_L g1815 ( 
.A(n_1776),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1781),
.Y(n_1816)
);

NAND2x1_ASAP7_75t_L g1817 ( 
.A(n_1787),
.B(n_1722),
.Y(n_1817)
);

OAI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1775),
.A2(n_1758),
.B(n_1713),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1781),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_SL g1820 ( 
.A1(n_1771),
.A2(n_1719),
.B1(n_1631),
.B2(n_1764),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1785),
.A2(n_1751),
.B1(n_1729),
.B2(n_1758),
.Y(n_1821)
);

A2O1A1Ixp33_ASAP7_75t_L g1822 ( 
.A1(n_1793),
.A2(n_1624),
.B(n_1651),
.C(n_1774),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1784),
.Y(n_1823)
);

INVx3_ASAP7_75t_L g1824 ( 
.A(n_1779),
.Y(n_1824)
);

BUFx6f_ASAP7_75t_SL g1825 ( 
.A(n_1779),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1789),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1783),
.B(n_1732),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1784),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1789),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1802),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1823),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1807),
.B(n_1776),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1807),
.B(n_1779),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1807),
.B(n_1786),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1810),
.B(n_1775),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1813),
.B(n_1788),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1807),
.B(n_1786),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1824),
.B(n_1815),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1802),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1828),
.Y(n_1840)
);

OAI211xp5_ASAP7_75t_L g1841 ( 
.A1(n_1812),
.A2(n_1721),
.B(n_1760),
.C(n_1787),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1824),
.B(n_1770),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1824),
.B(n_1770),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1805),
.B(n_1767),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1808),
.Y(n_1845)
);

OAI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1822),
.A2(n_1806),
.B1(n_1811),
.B2(n_1820),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1803),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1805),
.B(n_1767),
.Y(n_1848)
);

OAI221xp5_ASAP7_75t_L g1849 ( 
.A1(n_1800),
.A2(n_1794),
.B1(n_1780),
.B2(n_1797),
.C(n_1591),
.Y(n_1849)
);

OAI221xp5_ASAP7_75t_L g1850 ( 
.A1(n_1822),
.A2(n_1780),
.B1(n_1797),
.B2(n_1791),
.C(n_1790),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1803),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1808),
.B(n_1788),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1818),
.B(n_1798),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1804),
.B(n_1790),
.Y(n_1854)
);

AO21x2_ASAP7_75t_L g1855 ( 
.A1(n_1809),
.A2(n_1663),
.B(n_1657),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1816),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1816),
.Y(n_1857)
);

BUFx6f_ASAP7_75t_SL g1858 ( 
.A(n_1801),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1799),
.B(n_1791),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1817),
.B(n_1769),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1827),
.B(n_1732),
.Y(n_1861)
);

AO21x2_ASAP7_75t_L g1862 ( 
.A1(n_1804),
.A2(n_1639),
.B(n_1635),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1847),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1852),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1833),
.B(n_1821),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1833),
.B(n_1832),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1852),
.Y(n_1867)
);

INVxp67_ASAP7_75t_SL g1868 ( 
.A(n_1854),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1830),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1846),
.A2(n_1850),
.B1(n_1855),
.B2(n_1862),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1833),
.B(n_1814),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1838),
.B(n_1732),
.Y(n_1872)
);

INVx1_ASAP7_75t_SL g1873 ( 
.A(n_1832),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1847),
.Y(n_1874)
);

INVx1_ASAP7_75t_SL g1875 ( 
.A(n_1838),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1842),
.B(n_1801),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1851),
.B(n_1819),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1831),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1840),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_1834),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1835),
.Y(n_1881)
);

INVx3_ASAP7_75t_L g1882 ( 
.A(n_1834),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1844),
.B(n_1735),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1860),
.B(n_1725),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1844),
.B(n_1735),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1835),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1836),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1848),
.B(n_1860),
.Y(n_1888)
);

INVxp33_ASAP7_75t_L g1889 ( 
.A(n_1837),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1842),
.B(n_1843),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1859),
.B(n_1819),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1843),
.B(n_1801),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1848),
.B(n_1801),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1875),
.B(n_1859),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1881),
.B(n_1830),
.Y(n_1895)
);

OR2x6_ASAP7_75t_L g1896 ( 
.A(n_1866),
.B(n_1871),
.Y(n_1896)
);

INVxp67_ASAP7_75t_SL g1897 ( 
.A(n_1868),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1888),
.B(n_1853),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1888),
.B(n_1853),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1866),
.B(n_1837),
.Y(n_1900)
);

NAND2xp67_ASAP7_75t_L g1901 ( 
.A(n_1864),
.B(n_1839),
.Y(n_1901)
);

AND2x4_ASAP7_75t_L g1902 ( 
.A(n_1884),
.B(n_1801),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1863),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1863),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1893),
.B(n_1841),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1893),
.B(n_1855),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1865),
.B(n_1855),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1874),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1880),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1890),
.B(n_1861),
.Y(n_1910)
);

INVxp67_ASAP7_75t_SL g1911 ( 
.A(n_1870),
.Y(n_1911)
);

NOR2x1_ASAP7_75t_L g1912 ( 
.A(n_1874),
.B(n_1845),
.Y(n_1912)
);

INVxp67_ASAP7_75t_SL g1913 ( 
.A(n_1880),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1881),
.B(n_1839),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1865),
.B(n_1845),
.Y(n_1915)
);

INVx2_ASAP7_75t_SL g1916 ( 
.A(n_1880),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1878),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1878),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1879),
.Y(n_1919)
);

BUFx2_ASAP7_75t_L g1920 ( 
.A(n_1882),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1873),
.B(n_1887),
.Y(n_1921)
);

INVx2_ASAP7_75t_SL g1922 ( 
.A(n_1882),
.Y(n_1922)
);

AOI21xp33_ASAP7_75t_L g1923 ( 
.A1(n_1873),
.A2(n_1861),
.B(n_1862),
.Y(n_1923)
);

AOI211xp5_ASAP7_75t_SL g1924 ( 
.A1(n_1882),
.A2(n_1849),
.B(n_1604),
.C(n_1858),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1864),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1867),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1886),
.A2(n_1862),
.B(n_1856),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1883),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1876),
.B(n_1740),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1879),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1886),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1867),
.Y(n_1932)
);

INVxp67_ASAP7_75t_L g1933 ( 
.A(n_1877),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1887),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1871),
.A2(n_1858),
.B1(n_1857),
.B2(n_1856),
.Y(n_1935)
);

INVx2_ASAP7_75t_SL g1936 ( 
.A(n_1876),
.Y(n_1936)
);

NAND2x1_ASAP7_75t_L g1937 ( 
.A(n_1876),
.B(n_1825),
.Y(n_1937)
);

CKINVDCx16_ASAP7_75t_R g1938 ( 
.A(n_1896),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1897),
.B(n_1891),
.Y(n_1939)
);

BUFx6f_ASAP7_75t_L g1940 ( 
.A(n_1920),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1894),
.B(n_1889),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1913),
.Y(n_1942)
);

BUFx2_ASAP7_75t_L g1943 ( 
.A(n_1896),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1913),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1896),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1898),
.B(n_1876),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1925),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1897),
.B(n_1891),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1925),
.Y(n_1949)
);

BUFx3_ASAP7_75t_L g1950 ( 
.A(n_1936),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1911),
.B(n_1869),
.Y(n_1951)
);

AND2x4_ASAP7_75t_L g1952 ( 
.A(n_1915),
.B(n_1871),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1899),
.B(n_1883),
.Y(n_1953)
);

OAI33xp33_ASAP7_75t_L g1954 ( 
.A1(n_1931),
.A2(n_1872),
.A3(n_1869),
.B1(n_1892),
.B2(n_603),
.B3(n_598),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1900),
.B(n_1885),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1926),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1911),
.B(n_1885),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_L g1958 ( 
.A(n_1933),
.B(n_1871),
.Y(n_1958)
);

INVxp67_ASAP7_75t_L g1959 ( 
.A(n_1909),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1905),
.B(n_1733),
.Y(n_1960)
);

CKINVDCx5p33_ASAP7_75t_R g1961 ( 
.A(n_1902),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1926),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1932),
.Y(n_1963)
);

INVx4_ASAP7_75t_L g1964 ( 
.A(n_1909),
.Y(n_1964)
);

INVx1_ASAP7_75t_SL g1965 ( 
.A(n_1937),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1929),
.B(n_1733),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1928),
.B(n_1733),
.Y(n_1967)
);

HB1xp67_ASAP7_75t_L g1968 ( 
.A(n_1912),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1902),
.B(n_1748),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1932),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1903),
.Y(n_1971)
);

AO21x2_ASAP7_75t_L g1972 ( 
.A1(n_1927),
.A2(n_880),
.B(n_793),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1901),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1933),
.B(n_793),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1916),
.B(n_1748),
.Y(n_1975)
);

NOR2x1_ASAP7_75t_L g1976 ( 
.A(n_1921),
.B(n_907),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1934),
.B(n_1826),
.Y(n_1977)
);

BUFx2_ASAP7_75t_L g1978 ( 
.A(n_1922),
.Y(n_1978)
);

AOI22xp33_ASAP7_75t_L g1979 ( 
.A1(n_1907),
.A2(n_1858),
.B1(n_1577),
.B2(n_788),
.Y(n_1979)
);

NOR2x1_ASAP7_75t_L g1980 ( 
.A(n_1917),
.B(n_1918),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1904),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1910),
.B(n_1748),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1906),
.Y(n_1983)
);

INVx1_ASAP7_75t_SL g1984 ( 
.A(n_1895),
.Y(n_1984)
);

AOI22xp33_ASAP7_75t_L g1985 ( 
.A1(n_1923),
.A2(n_788),
.B1(n_806),
.B2(n_696),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1908),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1919),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1930),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1895),
.Y(n_1989)
);

INVx1_ASAP7_75t_SL g1990 ( 
.A(n_1914),
.Y(n_1990)
);

OAI21x1_ASAP7_75t_L g1991 ( 
.A1(n_1927),
.A2(n_1829),
.B(n_1826),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1914),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1935),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1924),
.B(n_1749),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1923),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1924),
.B(n_1829),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1907),
.B(n_555),
.Y(n_1997)
);

INVx1_ASAP7_75t_SL g1998 ( 
.A(n_1896),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1913),
.Y(n_1999)
);

HB1xp67_ASAP7_75t_L g2000 ( 
.A(n_1897),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1896),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1946),
.B(n_1825),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_2000),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_2000),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1942),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1940),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1953),
.B(n_1825),
.Y(n_2007)
);

CKINVDCx16_ASAP7_75t_R g2008 ( 
.A(n_1938),
.Y(n_2008)
);

NOR2x1p5_ASAP7_75t_SL g2009 ( 
.A(n_1945),
.B(n_2001),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1944),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1999),
.Y(n_2011)
);

AND2x4_ASAP7_75t_L g2012 ( 
.A(n_1950),
.B(n_1561),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1968),
.B(n_1980),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1940),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1968),
.B(n_591),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1939),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1955),
.B(n_1749),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1943),
.B(n_1749),
.Y(n_2018)
);

INVxp67_ASAP7_75t_L g2019 ( 
.A(n_1940),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1958),
.B(n_600),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_L g2021 ( 
.A(n_1961),
.B(n_806),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1960),
.B(n_1762),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1952),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1958),
.B(n_613),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1939),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1965),
.B(n_1522),
.Y(n_2026)
);

INVx1_ASAP7_75t_SL g2027 ( 
.A(n_1998),
.Y(n_2027)
);

INVx1_ASAP7_75t_SL g2028 ( 
.A(n_1978),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1969),
.B(n_1522),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1948),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1948),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1984),
.B(n_615),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1990),
.B(n_619),
.Y(n_2033)
);

NOR2xp33_ASAP7_75t_L g2034 ( 
.A(n_1954),
.B(n_885),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1952),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1995),
.B(n_627),
.Y(n_2036)
);

AND3x1_ASAP7_75t_L g2037 ( 
.A(n_1957),
.B(n_921),
.C(n_885),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1974),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1983),
.B(n_1964),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1964),
.Y(n_2040)
);

HB1xp67_ASAP7_75t_L g2041 ( 
.A(n_1959),
.Y(n_2041)
);

INVx2_ASAP7_75t_SL g2042 ( 
.A(n_1941),
.Y(n_2042)
);

CKINVDCx20_ASAP7_75t_R g2043 ( 
.A(n_1993),
.Y(n_2043)
);

INVx2_ASAP7_75t_SL g2044 ( 
.A(n_1966),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1982),
.B(n_1527),
.Y(n_2045)
);

OR2x2_ASAP7_75t_L g2046 ( 
.A(n_1957),
.B(n_1959),
.Y(n_2046)
);

NOR2xp33_ASAP7_75t_L g2047 ( 
.A(n_1954),
.B(n_921),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1974),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1967),
.B(n_1527),
.Y(n_2049)
);

INVx1_ASAP7_75t_SL g2050 ( 
.A(n_1951),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1991),
.Y(n_2051)
);

AND2x4_ASAP7_75t_L g2052 ( 
.A(n_1988),
.B(n_1524),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1947),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1989),
.B(n_631),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1976),
.Y(n_2055)
);

NAND2x1p5_ASAP7_75t_L g2056 ( 
.A(n_1997),
.B(n_1949),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1973),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1956),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1992),
.B(n_632),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_1987),
.B(n_1971),
.Y(n_2060)
);

NOR3xp33_ASAP7_75t_SL g2061 ( 
.A(n_1981),
.B(n_638),
.C(n_636),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1962),
.Y(n_2062)
);

INVxp67_ASAP7_75t_L g2063 ( 
.A(n_1951),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1975),
.B(n_640),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1986),
.B(n_641),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1994),
.B(n_646),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1972),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1972),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1963),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_1979),
.B(n_649),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1970),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1977),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1985),
.B(n_651),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_1979),
.B(n_652),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1985),
.B(n_654),
.Y(n_2075)
);

INVxp67_ASAP7_75t_L g2076 ( 
.A(n_1997),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1977),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1996),
.B(n_655),
.Y(n_2078)
);

OR2x2_ASAP7_75t_L g2079 ( 
.A(n_1996),
.B(n_0),
.Y(n_2079)
);

AOI31xp33_ASAP7_75t_L g2080 ( 
.A1(n_2000),
.A2(n_1576),
.A3(n_665),
.B(n_666),
.Y(n_2080)
);

OAI21xp33_ASAP7_75t_L g2081 ( 
.A1(n_1968),
.A2(n_667),
.B(n_656),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1946),
.B(n_669),
.Y(n_2082)
);

INVx2_ASAP7_75t_SL g2083 ( 
.A(n_1952),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2000),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1946),
.B(n_672),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1958),
.B(n_678),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1940),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2000),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2041),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2046),
.Y(n_2090)
);

AND2x4_ASAP7_75t_L g2091 ( 
.A(n_2083),
.B(n_1524),
.Y(n_2091)
);

NAND3xp33_ASAP7_75t_L g2092 ( 
.A(n_2063),
.B(n_2013),
.C(n_2008),
.Y(n_2092)
);

AOI22xp5_ASAP7_75t_L g2093 ( 
.A1(n_2050),
.A2(n_1642),
.B1(n_1602),
.B2(n_1582),
.Y(n_2093)
);

NAND2x1_ASAP7_75t_SL g2094 ( 
.A(n_2006),
.B(n_2014),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2027),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2002),
.B(n_681),
.Y(n_2096)
);

HB1xp67_ASAP7_75t_L g2097 ( 
.A(n_2050),
.Y(n_2097)
);

AOI32xp33_ASAP7_75t_L g2098 ( 
.A1(n_2037),
.A2(n_1642),
.A3(n_702),
.B1(n_706),
.B2(n_690),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2028),
.B(n_687),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2027),
.Y(n_2100)
);

OR2x2_ASAP7_75t_L g2101 ( 
.A(n_2028),
.B(n_1),
.Y(n_2101)
);

NAND3xp33_ASAP7_75t_L g2102 ( 
.A(n_2013),
.B(n_580),
.C(n_555),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_2021),
.B(n_709),
.Y(n_2103)
);

OAI322xp33_ASAP7_75t_L g2104 ( 
.A1(n_2016),
.A2(n_720),
.A3(n_722),
.B1(n_725),
.B2(n_729),
.C1(n_723),
.C2(n_718),
.Y(n_2104)
);

INVxp67_ASAP7_75t_L g2105 ( 
.A(n_2037),
.Y(n_2105)
);

AND2x2_ASAP7_75t_SL g2106 ( 
.A(n_2023),
.B(n_1647),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2003),
.Y(n_2107)
);

INVxp67_ASAP7_75t_SL g2108 ( 
.A(n_2019),
.Y(n_2108)
);

OAI21xp33_ASAP7_75t_L g2109 ( 
.A1(n_2042),
.A2(n_731),
.B(n_730),
.Y(n_2109)
);

AOI22xp33_ASAP7_75t_L g2110 ( 
.A1(n_2057),
.A2(n_1691),
.B1(n_1697),
.B2(n_1696),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2004),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2084),
.Y(n_2112)
);

AOI22xp5_ASAP7_75t_L g2113 ( 
.A1(n_2051),
.A2(n_1582),
.B1(n_954),
.B2(n_921),
.Y(n_2113)
);

NOR2xp33_ASAP7_75t_L g2114 ( 
.A(n_2044),
.B(n_743),
.Y(n_2114)
);

NOR3xp33_ASAP7_75t_SL g2115 ( 
.A(n_2039),
.B(n_748),
.C(n_747),
.Y(n_2115)
);

OAI22xp5_ASAP7_75t_L g2116 ( 
.A1(n_2035),
.A2(n_1751),
.B1(n_1729),
.B2(n_750),
.Y(n_2116)
);

AOI22xp5_ASAP7_75t_L g2117 ( 
.A1(n_2043),
.A2(n_1582),
.B1(n_1576),
.B2(n_1575),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2088),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2079),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2082),
.B(n_749),
.Y(n_2120)
);

OAI22xp33_ASAP7_75t_L g2121 ( 
.A1(n_2025),
.A2(n_1582),
.B1(n_1680),
.B2(n_1796),
.Y(n_2121)
);

AOI21xp5_ASAP7_75t_L g2122 ( 
.A1(n_2015),
.A2(n_759),
.B(n_752),
.Y(n_2122)
);

INVx1_ASAP7_75t_SL g2123 ( 
.A(n_2085),
.Y(n_2123)
);

OAI22xp5_ASAP7_75t_L g2124 ( 
.A1(n_2030),
.A2(n_766),
.B1(n_768),
.B2(n_762),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2012),
.B(n_2087),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2031),
.B(n_2),
.Y(n_2126)
);

OR2x2_ASAP7_75t_L g2127 ( 
.A(n_2020),
.B(n_2),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2007),
.B(n_769),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2012),
.B(n_771),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_2056),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2065),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_2040),
.B(n_787),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2060),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2064),
.B(n_790),
.Y(n_2134)
);

INVx3_ASAP7_75t_L g2135 ( 
.A(n_2052),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_2056),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2005),
.Y(n_2137)
);

OAI221xp5_ASAP7_75t_L g2138 ( 
.A1(n_2078),
.A2(n_796),
.B1(n_800),
.B2(n_795),
.C(n_792),
.Y(n_2138)
);

OAI21xp5_ASAP7_75t_L g2139 ( 
.A1(n_2018),
.A2(n_805),
.B(n_803),
.Y(n_2139)
);

OAI21xp5_ASAP7_75t_SL g2140 ( 
.A1(n_2026),
.A2(n_580),
.B(n_555),
.Y(n_2140)
);

AOI21xp5_ASAP7_75t_L g2141 ( 
.A1(n_2015),
.A2(n_811),
.B(n_807),
.Y(n_2141)
);

OR2x2_ASAP7_75t_L g2142 ( 
.A(n_2024),
.B(n_2086),
.Y(n_2142)
);

AOI22xp5_ASAP7_75t_L g2143 ( 
.A1(n_2034),
.A2(n_2047),
.B1(n_2078),
.B2(n_2066),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_2061),
.B(n_815),
.Y(n_2144)
);

OAI22xp33_ASAP7_75t_L g2145 ( 
.A1(n_2080),
.A2(n_1680),
.B1(n_1796),
.B2(n_1697),
.Y(n_2145)
);

OAI21xp33_ASAP7_75t_L g2146 ( 
.A1(n_2017),
.A2(n_824),
.B(n_822),
.Y(n_2146)
);

OAI21xp5_ASAP7_75t_SL g2147 ( 
.A1(n_2010),
.A2(n_659),
.B(n_580),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2011),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2072),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2081),
.B(n_826),
.Y(n_2150)
);

HB1xp67_ASAP7_75t_L g2151 ( 
.A(n_2071),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2077),
.Y(n_2152)
);

INVxp67_ASAP7_75t_L g2153 ( 
.A(n_2073),
.Y(n_2153)
);

OAI22xp33_ASAP7_75t_L g2154 ( 
.A1(n_2080),
.A2(n_1696),
.B1(n_1575),
.B2(n_1701),
.Y(n_2154)
);

AOI222xp33_ASAP7_75t_L g2155 ( 
.A1(n_2009),
.A2(n_836),
.B1(n_828),
.B2(n_842),
.C1(n_840),
.C2(n_831),
.Y(n_2155)
);

AOI222xp33_ASAP7_75t_L g2156 ( 
.A1(n_2036),
.A2(n_852),
.B1(n_848),
.B2(n_856),
.C1(n_854),
.C2(n_850),
.Y(n_2156)
);

OR2x2_ASAP7_75t_L g2157 ( 
.A(n_2032),
.B(n_3),
.Y(n_2157)
);

AOI31xp33_ASAP7_75t_L g2158 ( 
.A1(n_2081),
.A2(n_2053),
.A3(n_2062),
.B(n_2058),
.Y(n_2158)
);

AOI32xp33_ASAP7_75t_L g2159 ( 
.A1(n_2069),
.A2(n_861),
.A3(n_864),
.B1(n_862),
.B2(n_857),
.Y(n_2159)
);

A2O1A1Ixp33_ASAP7_75t_L g2160 ( 
.A1(n_2033),
.A2(n_887),
.B(n_888),
.C(n_881),
.Y(n_2160)
);

OAI21xp5_ASAP7_75t_L g2161 ( 
.A1(n_2052),
.A2(n_892),
.B(n_891),
.Y(n_2161)
);

OAI21xp33_ASAP7_75t_SL g2162 ( 
.A1(n_2036),
.A2(n_1621),
.B(n_1619),
.Y(n_2162)
);

AOI221xp5_ASAP7_75t_L g2163 ( 
.A1(n_2059),
.A2(n_899),
.B1(n_903),
.B2(n_896),
.C(n_893),
.Y(n_2163)
);

AOI22xp5_ASAP7_75t_L g2164 ( 
.A1(n_2073),
.A2(n_908),
.B1(n_911),
.B2(n_905),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2070),
.B(n_915),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2054),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2074),
.B(n_922),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2059),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2075),
.B(n_924),
.Y(n_2169)
);

AOI221xp5_ASAP7_75t_L g2170 ( 
.A1(n_2038),
.A2(n_2048),
.B1(n_2075),
.B2(n_2067),
.C(n_2068),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2076),
.Y(n_2171)
);

OAI22xp33_ASAP7_75t_L g2172 ( 
.A1(n_2055),
.A2(n_1701),
.B1(n_1704),
.B2(n_1709),
.Y(n_2172)
);

NAND2xp33_ASAP7_75t_SL g2173 ( 
.A(n_2045),
.B(n_925),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_2029),
.B(n_927),
.Y(n_2174)
);

AOI22xp33_ASAP7_75t_L g2175 ( 
.A1(n_2022),
.A2(n_1690),
.B1(n_1695),
.B2(n_1704),
.Y(n_2175)
);

AOI22xp33_ASAP7_75t_L g2176 ( 
.A1(n_2049),
.A2(n_1690),
.B1(n_1695),
.B2(n_955),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2041),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2008),
.B(n_928),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_2002),
.B(n_929),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2002),
.B(n_935),
.Y(n_2180)
);

OAI221xp5_ASAP7_75t_L g2181 ( 
.A1(n_2050),
.A2(n_953),
.B1(n_944),
.B2(n_580),
.C(n_798),
.Y(n_2181)
);

INVx1_ASAP7_75t_SL g2182 ( 
.A(n_2008),
.Y(n_2182)
);

INVx2_ASAP7_75t_SL g2183 ( 
.A(n_2002),
.Y(n_2183)
);

OAI22xp5_ASAP7_75t_L g2184 ( 
.A1(n_2050),
.A2(n_733),
.B1(n_798),
.B2(n_659),
.Y(n_2184)
);

A2O1A1Ixp33_ASAP7_75t_L g2185 ( 
.A1(n_2050),
.A2(n_1621),
.B(n_941),
.C(n_952),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2041),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2041),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_L g2188 ( 
.A(n_2008),
.B(n_3),
.Y(n_2188)
);

AOI322xp5_ASAP7_75t_L g2189 ( 
.A1(n_2050),
.A2(n_1537),
.A3(n_1693),
.B1(n_1692),
.B2(n_1699),
.C1(n_1551),
.C2(n_1728),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2008),
.B(n_659),
.Y(n_2190)
);

OAI22xp5_ASAP7_75t_L g2191 ( 
.A1(n_2050),
.A2(n_733),
.B1(n_798),
.B2(n_659),
.Y(n_2191)
);

OR2x2_ASAP7_75t_L g2192 ( 
.A(n_2046),
.B(n_4),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2041),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2041),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2041),
.Y(n_2195)
);

OAI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_2050),
.A2(n_798),
.B1(n_941),
.B2(n_733),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2041),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2041),
.Y(n_2198)
);

AOI22xp33_ASAP7_75t_SL g2199 ( 
.A1(n_2050),
.A2(n_733),
.B1(n_952),
.B2(n_941),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2002),
.B(n_4),
.Y(n_2200)
);

AOI22xp5_ASAP7_75t_L g2201 ( 
.A1(n_2008),
.A2(n_1547),
.B1(n_952),
.B2(n_941),
.Y(n_2201)
);

OAI21xp5_ASAP7_75t_L g2202 ( 
.A1(n_2063),
.A2(n_1619),
.B(n_1654),
.Y(n_2202)
);

AOI22xp5_ASAP7_75t_L g2203 ( 
.A1(n_2008),
.A2(n_1547),
.B1(n_952),
.B2(n_1562),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2041),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2008),
.Y(n_2205)
);

OAI32xp33_ASAP7_75t_L g2206 ( 
.A1(n_2050),
.A2(n_1709),
.A3(n_1544),
.B1(n_1559),
.B2(n_1549),
.Y(n_2206)
);

AOI21xp5_ASAP7_75t_L g2207 ( 
.A1(n_2013),
.A2(n_877),
.B(n_876),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2041),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_SL g2209 ( 
.A(n_2008),
.B(n_834),
.Y(n_2209)
);

OR2x2_ASAP7_75t_L g2210 ( 
.A(n_2046),
.B(n_5),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2041),
.Y(n_2211)
);

HB1xp67_ASAP7_75t_L g2212 ( 
.A(n_2050),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2041),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2002),
.B(n_6),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2008),
.B(n_6),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2041),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2008),
.B(n_7),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_SL g2218 ( 
.A(n_2008),
.B(n_1544),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2008),
.B(n_7),
.Y(n_2219)
);

OAI21xp5_ASAP7_75t_L g2220 ( 
.A1(n_2063),
.A2(n_1656),
.B(n_1654),
.Y(n_2220)
);

OAI211xp5_ASAP7_75t_SL g2221 ( 
.A1(n_2013),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2041),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2008),
.B(n_8),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2008),
.B(n_9),
.Y(n_2224)
);

INVx2_ASAP7_75t_SL g2225 ( 
.A(n_2002),
.Y(n_2225)
);

NOR2xp33_ASAP7_75t_SL g2226 ( 
.A(n_2008),
.B(n_1563),
.Y(n_2226)
);

NOR2xp33_ASAP7_75t_L g2227 ( 
.A(n_2008),
.B(n_10),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2002),
.B(n_11),
.Y(n_2228)
);

OAI21xp33_ASAP7_75t_L g2229 ( 
.A1(n_2027),
.A2(n_1669),
.B(n_1700),
.Y(n_2229)
);

HB1xp67_ASAP7_75t_L g2230 ( 
.A(n_2050),
.Y(n_2230)
);

OAI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_2050),
.A2(n_1709),
.B1(n_1730),
.B2(n_1693),
.Y(n_2231)
);

INVx1_ASAP7_75t_SL g2232 ( 
.A(n_2008),
.Y(n_2232)
);

NOR3xp33_ASAP7_75t_L g2233 ( 
.A(n_2008),
.B(n_1656),
.C(n_877),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2008),
.B(n_13),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2041),
.Y(n_2235)
);

OAI22xp5_ASAP7_75t_L g2236 ( 
.A1(n_2050),
.A2(n_1699),
.B1(n_1692),
.B2(n_1700),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2008),
.B(n_15),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2008),
.B(n_16),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2182),
.B(n_17),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_2232),
.B(n_18),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2205),
.B(n_19),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2097),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2212),
.Y(n_2243)
);

NAND3xp33_ASAP7_75t_L g2244 ( 
.A(n_2230),
.B(n_868),
.C(n_858),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2192),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2210),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2094),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2151),
.Y(n_2248)
);

XNOR2xp5_ASAP7_75t_L g2249 ( 
.A(n_2092),
.B(n_20),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2095),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2100),
.B(n_21),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2123),
.B(n_21),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2101),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_2188),
.B(n_22),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2215),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_2108),
.B(n_22),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2217),
.Y(n_2257)
);

OR2x2_ASAP7_75t_L g2258 ( 
.A(n_2090),
.B(n_2133),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2227),
.B(n_23),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2219),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2155),
.B(n_23),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_2129),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_SL g2263 ( 
.A(n_2130),
.B(n_537),
.Y(n_2263)
);

INVxp67_ASAP7_75t_L g2264 ( 
.A(n_2223),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2224),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2099),
.B(n_24),
.Y(n_2266)
);

AND2x4_ASAP7_75t_L g2267 ( 
.A(n_2183),
.B(n_24),
.Y(n_2267)
);

INVxp67_ASAP7_75t_L g2268 ( 
.A(n_2234),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2237),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2238),
.Y(n_2270)
);

BUFx2_ASAP7_75t_L g2271 ( 
.A(n_2200),
.Y(n_2271)
);

INVxp67_ASAP7_75t_SL g2272 ( 
.A(n_2178),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2126),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2119),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2127),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2131),
.B(n_2214),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2157),
.Y(n_2277)
);

NOR2xp33_ASAP7_75t_L g2278 ( 
.A(n_2221),
.B(n_25),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2132),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2228),
.B(n_25),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_SL g2281 ( 
.A(n_2136),
.B(n_537),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2135),
.B(n_26),
.Y(n_2282)
);

INVxp67_ASAP7_75t_L g2283 ( 
.A(n_2226),
.Y(n_2283)
);

NAND2xp33_ASAP7_75t_SL g2284 ( 
.A(n_2115),
.B(n_27),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2225),
.B(n_27),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2135),
.B(n_28),
.Y(n_2286)
);

OAI21xp5_ASAP7_75t_L g2287 ( 
.A1(n_2089),
.A2(n_1635),
.B(n_1630),
.Y(n_2287)
);

AND2x2_ASAP7_75t_L g2288 ( 
.A(n_2128),
.B(n_28),
.Y(n_2288)
);

NAND2x1_ASAP7_75t_L g2289 ( 
.A(n_2091),
.B(n_2158),
.Y(n_2289)
);

INVxp67_ASAP7_75t_L g2290 ( 
.A(n_2173),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2174),
.B(n_29),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2156),
.B(n_30),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2177),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_2106),
.Y(n_2294)
);

NAND2xp33_ASAP7_75t_L g2295 ( 
.A(n_2186),
.B(n_693),
.Y(n_2295)
);

INVxp67_ASAP7_75t_SL g2296 ( 
.A(n_2144),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2114),
.B(n_30),
.Y(n_2297)
);

INVxp67_ASAP7_75t_L g2298 ( 
.A(n_2125),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2187),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2193),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2194),
.Y(n_2301)
);

HB1xp67_ASAP7_75t_L g2302 ( 
.A(n_2195),
.Y(n_2302)
);

HB1xp67_ASAP7_75t_L g2303 ( 
.A(n_2197),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2096),
.B(n_31),
.Y(n_2304)
);

OR2x2_ASAP7_75t_L g2305 ( 
.A(n_2198),
.B(n_32),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2159),
.B(n_33),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2164),
.B(n_34),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2204),
.Y(n_2308)
);

NOR2xp33_ASAP7_75t_L g2309 ( 
.A(n_2104),
.B(n_36),
.Y(n_2309)
);

OA21x2_ASAP7_75t_SL g2310 ( 
.A1(n_2218),
.A2(n_36),
.B(n_37),
.Y(n_2310)
);

AOI22x1_ASAP7_75t_L g2311 ( 
.A1(n_2208),
.A2(n_2213),
.B1(n_2216),
.B2(n_2211),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2164),
.B(n_38),
.Y(n_2312)
);

NAND2xp33_ASAP7_75t_SL g2313 ( 
.A(n_2222),
.B(n_38),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2235),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2168),
.B(n_39),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2179),
.B(n_40),
.Y(n_2316)
);

HB1xp67_ASAP7_75t_L g2317 ( 
.A(n_2107),
.Y(n_2317)
);

OR2x2_ASAP7_75t_L g2318 ( 
.A(n_2171),
.B(n_40),
.Y(n_2318)
);

INVx1_ASAP7_75t_SL g2319 ( 
.A(n_2180),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2160),
.B(n_41),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2190),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2142),
.Y(n_2322)
);

CKINVDCx20_ASAP7_75t_R g2323 ( 
.A(n_2143),
.Y(n_2323)
);

INVx1_ASAP7_75t_SL g2324 ( 
.A(n_2120),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2091),
.B(n_41),
.Y(n_2325)
);

INVxp33_ASAP7_75t_L g2326 ( 
.A(n_2134),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2105),
.B(n_43),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2169),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_SL g2329 ( 
.A(n_2098),
.B(n_955),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2111),
.B(n_43),
.Y(n_2330)
);

INVxp67_ASAP7_75t_L g2331 ( 
.A(n_2150),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2149),
.B(n_44),
.Y(n_2332)
);

HB1xp67_ASAP7_75t_L g2333 ( 
.A(n_2112),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2165),
.Y(n_2334)
);

OR2x2_ASAP7_75t_L g2335 ( 
.A(n_2118),
.B(n_44),
.Y(n_2335)
);

NOR2xp67_ASAP7_75t_L g2336 ( 
.A(n_2137),
.B(n_45),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2152),
.B(n_45),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2167),
.Y(n_2338)
);

OR2x2_ASAP7_75t_L g2339 ( 
.A(n_2148),
.B(n_46),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2146),
.B(n_46),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2166),
.B(n_47),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2153),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2103),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2124),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2207),
.B(n_47),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2109),
.B(n_48),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2163),
.B(n_49),
.Y(n_2347)
);

INVxp67_ASAP7_75t_L g2348 ( 
.A(n_2138),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_SL g2349 ( 
.A(n_2116),
.B(n_2139),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2161),
.B(n_50),
.Y(n_2350)
);

AOI22xp33_ASAP7_75t_L g2351 ( 
.A1(n_2170),
.A2(n_955),
.B1(n_868),
.B2(n_858),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2209),
.B(n_51),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2122),
.B(n_52),
.Y(n_2353)
);

NOR2xp33_ASAP7_75t_L g2354 ( 
.A(n_2181),
.B(n_52),
.Y(n_2354)
);

AOI21xp5_ASAP7_75t_L g2355 ( 
.A1(n_2141),
.A2(n_909),
.B(n_895),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2113),
.Y(n_2356)
);

OAI21xp33_ASAP7_75t_L g2357 ( 
.A1(n_2147),
.A2(n_2201),
.B(n_2140),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2271),
.Y(n_2358)
);

OR2x2_ASAP7_75t_L g2359 ( 
.A(n_2258),
.B(n_2184),
.Y(n_2359)
);

AND2x2_ASAP7_75t_L g2360 ( 
.A(n_2247),
.B(n_2239),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2256),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2276),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2240),
.Y(n_2363)
);

OAI31xp33_ASAP7_75t_L g2364 ( 
.A1(n_2313),
.A2(n_2154),
.A3(n_2145),
.B(n_2185),
.Y(n_2364)
);

OR2x2_ASAP7_75t_L g2365 ( 
.A(n_2248),
.B(n_2191),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_SL g2366 ( 
.A(n_2267),
.B(n_2319),
.Y(n_2366)
);

NAND3xp33_ASAP7_75t_L g2367 ( 
.A(n_2311),
.B(n_2199),
.C(n_2102),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2267),
.B(n_2196),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2319),
.B(n_2203),
.Y(n_2369)
);

AND2x2_ASAP7_75t_L g2370 ( 
.A(n_2285),
.B(n_2093),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2322),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_2298),
.B(n_2229),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2280),
.Y(n_2373)
);

HB1xp67_ASAP7_75t_L g2374 ( 
.A(n_2289),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2288),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_SL g2376 ( 
.A(n_2242),
.B(n_2162),
.Y(n_2376)
);

NAND3xp33_ASAP7_75t_L g2377 ( 
.A(n_2317),
.B(n_2233),
.C(n_2176),
.Y(n_2377)
);

AND2x4_ASAP7_75t_L g2378 ( 
.A(n_2251),
.B(n_2117),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2304),
.B(n_2110),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2336),
.Y(n_2380)
);

INVxp67_ASAP7_75t_L g2381 ( 
.A(n_2284),
.Y(n_2381)
);

OAI22xp5_ASAP7_75t_L g2382 ( 
.A1(n_2243),
.A2(n_2175),
.B1(n_2231),
.B2(n_2236),
.Y(n_2382)
);

NOR2x1_ASAP7_75t_L g2383 ( 
.A(n_2249),
.B(n_2172),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2278),
.B(n_2162),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2245),
.B(n_2189),
.Y(n_2385)
);

OR2x2_ASAP7_75t_L g2386 ( 
.A(n_2302),
.B(n_2303),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2246),
.B(n_2206),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2318),
.Y(n_2388)
);

AOI31xp33_ASAP7_75t_L g2389 ( 
.A1(n_2250),
.A2(n_2274),
.A3(n_2333),
.B(n_2299),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2337),
.Y(n_2390)
);

AND2x2_ASAP7_75t_L g2391 ( 
.A(n_2293),
.B(n_2202),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2330),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_2339),
.Y(n_2393)
);

AND2x4_ASAP7_75t_L g2394 ( 
.A(n_2262),
.B(n_2220),
.Y(n_2394)
);

NAND2x1_ASAP7_75t_SL g2395 ( 
.A(n_2325),
.B(n_2121),
.Y(n_2395)
);

INVxp67_ASAP7_75t_L g2396 ( 
.A(n_2254),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_SL g2397 ( 
.A(n_2253),
.B(n_693),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2275),
.B(n_53),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_2300),
.B(n_53),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2252),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2335),
.Y(n_2401)
);

NOR2x1_ASAP7_75t_L g2402 ( 
.A(n_2305),
.B(n_54),
.Y(n_2402)
);

INVxp67_ASAP7_75t_L g2403 ( 
.A(n_2316),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2282),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2286),
.Y(n_2405)
);

NOR2xp33_ASAP7_75t_L g2406 ( 
.A(n_2326),
.B(n_55),
.Y(n_2406)
);

NAND3xp33_ASAP7_75t_L g2407 ( 
.A(n_2264),
.B(n_589),
.C(n_527),
.Y(n_2407)
);

NOR2xp33_ASAP7_75t_L g2408 ( 
.A(n_2268),
.B(n_55),
.Y(n_2408)
);

INVx2_ASAP7_75t_SL g2409 ( 
.A(n_2241),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2277),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2266),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2273),
.B(n_56),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2324),
.B(n_57),
.Y(n_2413)
);

INVxp33_ASAP7_75t_L g2414 ( 
.A(n_2259),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2324),
.B(n_57),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2353),
.Y(n_2416)
);

INVx3_ASAP7_75t_L g2417 ( 
.A(n_2255),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2315),
.Y(n_2418)
);

HB1xp67_ASAP7_75t_L g2419 ( 
.A(n_2283),
.Y(n_2419)
);

OR2x2_ASAP7_75t_L g2420 ( 
.A(n_2332),
.B(n_59),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2291),
.Y(n_2421)
);

NOR2xp33_ASAP7_75t_L g2422 ( 
.A(n_2257),
.B(n_59),
.Y(n_2422)
);

AOI22xp5_ASAP7_75t_L g2423 ( 
.A1(n_2296),
.A2(n_1562),
.B1(n_1708),
.B2(n_1630),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2350),
.B(n_2352),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2260),
.B(n_60),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2323),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_2301),
.B(n_60),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2341),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2307),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2265),
.B(n_61),
.Y(n_2430)
);

INVxp67_ASAP7_75t_L g2431 ( 
.A(n_2309),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2269),
.B(n_62),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2312),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2270),
.B(n_63),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2340),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2272),
.B(n_63),
.Y(n_2436)
);

AND2x2_ASAP7_75t_L g2437 ( 
.A(n_2308),
.B(n_2314),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2342),
.B(n_64),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2292),
.Y(n_2439)
);

AND2x2_ASAP7_75t_L g2440 ( 
.A(n_2279),
.B(n_64),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_SL g2441 ( 
.A(n_2294),
.B(n_693),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2334),
.B(n_65),
.Y(n_2442)
);

OAI22xp5_ASAP7_75t_L g2443 ( 
.A1(n_2306),
.A2(n_1705),
.B1(n_1562),
.B2(n_1708),
.Y(n_2443)
);

AND2x2_ASAP7_75t_L g2444 ( 
.A(n_2343),
.B(n_66),
.Y(n_2444)
);

AND2x2_ASAP7_75t_L g2445 ( 
.A(n_2344),
.B(n_67),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2345),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_2349),
.B(n_68),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_2348),
.B(n_68),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2327),
.Y(n_2449)
);

NOR2xp33_ASAP7_75t_L g2450 ( 
.A(n_2261),
.B(n_69),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2338),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2297),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_2328),
.B(n_69),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2354),
.B(n_2290),
.Y(n_2454)
);

INVx1_ASAP7_75t_SL g2455 ( 
.A(n_2320),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2347),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2346),
.Y(n_2457)
);

HB1xp67_ASAP7_75t_L g2458 ( 
.A(n_2321),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_2331),
.B(n_71),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2355),
.B(n_72),
.Y(n_2460)
);

NOR2xp33_ASAP7_75t_L g2461 ( 
.A(n_2329),
.B(n_72),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2244),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2244),
.Y(n_2463)
);

INVxp67_ASAP7_75t_L g2464 ( 
.A(n_2263),
.Y(n_2464)
);

AND2x2_ASAP7_75t_L g2465 ( 
.A(n_2356),
.B(n_73),
.Y(n_2465)
);

INVxp67_ASAP7_75t_L g2466 ( 
.A(n_2281),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2295),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2357),
.Y(n_2468)
);

NOR2xp33_ASAP7_75t_L g2469 ( 
.A(n_2357),
.B(n_74),
.Y(n_2469)
);

INVx1_ASAP7_75t_SL g2470 ( 
.A(n_2310),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2351),
.B(n_75),
.Y(n_2471)
);

INVx3_ASAP7_75t_L g2472 ( 
.A(n_2287),
.Y(n_2472)
);

OR2x2_ASAP7_75t_L g2473 ( 
.A(n_2258),
.B(n_76),
.Y(n_2473)
);

NOR2x1_ASAP7_75t_L g2474 ( 
.A(n_2247),
.B(n_76),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2271),
.Y(n_2475)
);

OAI21xp5_ASAP7_75t_SL g2476 ( 
.A1(n_2247),
.A2(n_77),
.B(n_78),
.Y(n_2476)
);

AND2x2_ASAP7_75t_L g2477 ( 
.A(n_2247),
.B(n_77),
.Y(n_2477)
);

NOR2xp33_ASAP7_75t_L g2478 ( 
.A(n_2271),
.B(n_79),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2271),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2271),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2271),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2271),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2271),
.B(n_79),
.Y(n_2483)
);

INVx1_ASAP7_75t_SL g2484 ( 
.A(n_2271),
.Y(n_2484)
);

INVxp67_ASAP7_75t_L g2485 ( 
.A(n_2271),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2271),
.B(n_80),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2271),
.B(n_80),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_2247),
.B(n_81),
.Y(n_2488)
);

OR2x2_ASAP7_75t_L g2489 ( 
.A(n_2258),
.B(n_81),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2271),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2271),
.B(n_82),
.Y(n_2491)
);

INVx1_ASAP7_75t_SL g2492 ( 
.A(n_2271),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2271),
.B(n_82),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2271),
.B(n_84),
.Y(n_2494)
);

AND2x2_ASAP7_75t_L g2495 ( 
.A(n_2247),
.B(n_84),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2271),
.Y(n_2496)
);

NOR2xp33_ASAP7_75t_L g2497 ( 
.A(n_2271),
.B(n_85),
.Y(n_2497)
);

INVx2_ASAP7_75t_SL g2498 ( 
.A(n_2267),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2271),
.B(n_86),
.Y(n_2499)
);

OAI22xp5_ASAP7_75t_L g2500 ( 
.A1(n_2247),
.A2(n_1705),
.B1(n_1558),
.B2(n_1573),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2271),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2271),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2271),
.Y(n_2503)
);

AND2x2_ASAP7_75t_L g2504 ( 
.A(n_2247),
.B(n_86),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2271),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2247),
.B(n_87),
.Y(n_2506)
);

AOI221xp5_ASAP7_75t_L g2507 ( 
.A1(n_2376),
.A2(n_639),
.B1(n_933),
.B2(n_566),
.C(n_548),
.Y(n_2507)
);

CKINVDCx20_ASAP7_75t_R g2508 ( 
.A(n_2419),
.Y(n_2508)
);

NOR4xp25_ASAP7_75t_L g2509 ( 
.A(n_2484),
.B(n_89),
.C(n_87),
.D(n_88),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_2470),
.B(n_88),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2386),
.Y(n_2511)
);

AOI321xp33_ASAP7_75t_L g2512 ( 
.A1(n_2383),
.A2(n_2426),
.A3(n_2382),
.B1(n_2366),
.B2(n_2360),
.C(n_2372),
.Y(n_2512)
);

AOI211x1_ASAP7_75t_L g2513 ( 
.A1(n_2389),
.A2(n_92),
.B(n_90),
.C(n_91),
.Y(n_2513)
);

AND2x2_ASAP7_75t_L g2514 ( 
.A(n_2492),
.B(n_91),
.Y(n_2514)
);

NOR4xp25_ASAP7_75t_L g2515 ( 
.A(n_2485),
.B(n_96),
.C(n_93),
.D(n_94),
.Y(n_2515)
);

NAND4xp25_ASAP7_75t_L g2516 ( 
.A(n_2358),
.B(n_97),
.C(n_93),
.D(n_96),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2498),
.B(n_97),
.Y(n_2517)
);

NAND4xp75_ASAP7_75t_L g2518 ( 
.A(n_2474),
.B(n_100),
.C(n_98),
.D(n_99),
.Y(n_2518)
);

NAND2x1p5_ASAP7_75t_L g2519 ( 
.A(n_2474),
.B(n_98),
.Y(n_2519)
);

AOI21xp5_ASAP7_75t_SL g2520 ( 
.A1(n_2475),
.A2(n_2480),
.B(n_2479),
.Y(n_2520)
);

OAI21xp33_ASAP7_75t_L g2521 ( 
.A1(n_2468),
.A2(n_1669),
.B(n_1711),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_L g2522 ( 
.A(n_2478),
.B(n_99),
.Y(n_2522)
);

AOI21xp5_ASAP7_75t_L g2523 ( 
.A1(n_2374),
.A2(n_100),
.B(n_103),
.Y(n_2523)
);

NOR2x1_ASAP7_75t_L g2524 ( 
.A(n_2481),
.B(n_104),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2402),
.Y(n_2525)
);

OR2x2_ASAP7_75t_L g2526 ( 
.A(n_2482),
.B(n_105),
.Y(n_2526)
);

NAND3xp33_ASAP7_75t_SL g2527 ( 
.A(n_2490),
.B(n_2501),
.C(n_2496),
.Y(n_2527)
);

BUFx2_ASAP7_75t_SL g2528 ( 
.A(n_2502),
.Y(n_2528)
);

NAND3xp33_ASAP7_75t_L g2529 ( 
.A(n_2497),
.B(n_2367),
.C(n_2503),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2444),
.B(n_106),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2402),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_SL g2532 ( 
.A(n_2505),
.B(n_693),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2453),
.B(n_107),
.Y(n_2533)
);

NAND5xp2_ASAP7_75t_L g2534 ( 
.A(n_2363),
.B(n_109),
.C(n_107),
.D(n_108),
.E(n_110),
.Y(n_2534)
);

NOR3xp33_ASAP7_75t_L g2535 ( 
.A(n_2483),
.B(n_529),
.C(n_526),
.Y(n_2535)
);

NAND5xp2_ASAP7_75t_L g2536 ( 
.A(n_2362),
.B(n_111),
.C(n_108),
.D(n_110),
.E(n_113),
.Y(n_2536)
);

INVxp33_ASAP7_75t_L g2537 ( 
.A(n_2406),
.Y(n_2537)
);

AOI22xp5_ASAP7_75t_L g2538 ( 
.A1(n_2439),
.A2(n_1645),
.B1(n_1618),
.B2(n_1540),
.Y(n_2538)
);

NOR3xp33_ASAP7_75t_L g2539 ( 
.A(n_2486),
.B(n_536),
.C(n_530),
.Y(n_2539)
);

NAND3xp33_ASAP7_75t_L g2540 ( 
.A(n_2381),
.B(n_589),
.C(n_549),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2447),
.B(n_117),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2473),
.Y(n_2542)
);

NOR4xp25_ASAP7_75t_SL g2543 ( 
.A(n_2476),
.B(n_120),
.C(n_118),
.D(n_119),
.Y(n_2543)
);

NOR2xp33_ASAP7_75t_SL g2544 ( 
.A(n_2361),
.B(n_541),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2489),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2440),
.Y(n_2546)
);

HB1xp67_ASAP7_75t_L g2547 ( 
.A(n_2487),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2375),
.Y(n_2548)
);

NAND3xp33_ASAP7_75t_L g2549 ( 
.A(n_2422),
.B(n_589),
.C(n_584),
.Y(n_2549)
);

AOI221xp5_ASAP7_75t_L g2550 ( 
.A1(n_2384),
.A2(n_589),
.B1(n_599),
.B2(n_604),
.C(n_583),
.Y(n_2550)
);

NAND2xp33_ASAP7_75t_L g2551 ( 
.A(n_2458),
.B(n_693),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2413),
.Y(n_2552)
);

NOR2xp33_ASAP7_75t_L g2553 ( 
.A(n_2417),
.B(n_120),
.Y(n_2553)
);

NAND3xp33_ASAP7_75t_L g2554 ( 
.A(n_2469),
.B(n_612),
.C(n_605),
.Y(n_2554)
);

AOI22xp33_ASAP7_75t_L g2555 ( 
.A1(n_2380),
.A2(n_693),
.B1(n_1675),
.B2(n_1671),
.Y(n_2555)
);

XOR2x2_ASAP7_75t_L g2556 ( 
.A(n_2383),
.B(n_123),
.Y(n_2556)
);

AOI221xp5_ASAP7_75t_L g2557 ( 
.A1(n_2472),
.A2(n_2418),
.B1(n_2446),
.B2(n_2428),
.C(n_2416),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2415),
.Y(n_2558)
);

OAI221xp5_ASAP7_75t_L g2559 ( 
.A1(n_2387),
.A2(n_622),
.B1(n_624),
.B2(n_621),
.C(n_617),
.Y(n_2559)
);

BUFx2_ASAP7_75t_L g2560 ( 
.A(n_2417),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2491),
.Y(n_2561)
);

NOR2xp33_ASAP7_75t_L g2562 ( 
.A(n_2414),
.B(n_125),
.Y(n_2562)
);

HB1xp67_ASAP7_75t_L g2563 ( 
.A(n_2493),
.Y(n_2563)
);

OAI211xp5_ASAP7_75t_L g2564 ( 
.A1(n_2371),
.A2(n_130),
.B(n_128),
.C(n_129),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2494),
.Y(n_2565)
);

NOR2xp33_ASAP7_75t_R g2566 ( 
.A(n_2437),
.B(n_131),
.Y(n_2566)
);

NOR2xp33_ASAP7_75t_L g2567 ( 
.A(n_2499),
.B(n_132),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_SL g2568 ( 
.A(n_2451),
.B(n_2390),
.Y(n_2568)
);

NOR2xp33_ASAP7_75t_L g2569 ( 
.A(n_2392),
.B(n_133),
.Y(n_2569)
);

INVxp67_ASAP7_75t_SL g2570 ( 
.A(n_2368),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2399),
.B(n_135),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2427),
.Y(n_2572)
);

OAI211xp5_ASAP7_75t_L g2573 ( 
.A1(n_2410),
.A2(n_139),
.B(n_136),
.C(n_137),
.Y(n_2573)
);

INVxp67_ASAP7_75t_L g2574 ( 
.A(n_2424),
.Y(n_2574)
);

NOR4xp25_ASAP7_75t_L g2575 ( 
.A(n_2401),
.B(n_139),
.C(n_136),
.D(n_137),
.Y(n_2575)
);

AND2x2_ASAP7_75t_L g2576 ( 
.A(n_2477),
.B(n_140),
.Y(n_2576)
);

NAND4xp25_ASAP7_75t_L g2577 ( 
.A(n_2377),
.B(n_142),
.C(n_140),
.D(n_141),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_SL g2578 ( 
.A(n_2488),
.B(n_2495),
.Y(n_2578)
);

NAND3xp33_ASAP7_75t_L g2579 ( 
.A(n_2408),
.B(n_626),
.C(n_625),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2445),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2393),
.B(n_2409),
.Y(n_2581)
);

NAND4xp25_ASAP7_75t_SL g2582 ( 
.A(n_2391),
.B(n_2379),
.C(n_2506),
.D(n_2504),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2459),
.B(n_142),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_SL g2584 ( 
.A(n_2359),
.B(n_693),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2388),
.B(n_143),
.Y(n_2585)
);

NOR3xp33_ASAP7_75t_SL g2586 ( 
.A(n_2438),
.B(n_144),
.C(n_145),
.Y(n_2586)
);

OAI211xp5_ASAP7_75t_L g2587 ( 
.A1(n_2431),
.A2(n_148),
.B(n_146),
.C(n_147),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2420),
.Y(n_2588)
);

AND2x2_ASAP7_75t_L g2589 ( 
.A(n_2452),
.B(n_146),
.Y(n_2589)
);

INVx1_ASAP7_75t_SL g2590 ( 
.A(n_2436),
.Y(n_2590)
);

O2A1O1Ixp33_ASAP7_75t_L g2591 ( 
.A1(n_2398),
.A2(n_150),
.B(n_147),
.C(n_149),
.Y(n_2591)
);

NOR3xp33_ASAP7_75t_SL g2592 ( 
.A(n_2404),
.B(n_149),
.C(n_150),
.Y(n_2592)
);

NOR2xp33_ASAP7_75t_L g2593 ( 
.A(n_2373),
.B(n_151),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_SL g2594 ( 
.A(n_2364),
.B(n_629),
.Y(n_2594)
);

OAI22xp33_ASAP7_75t_L g2595 ( 
.A1(n_2508),
.A2(n_2412),
.B1(n_2430),
.B2(n_2425),
.Y(n_2595)
);

AOI221xp5_ASAP7_75t_L g2596 ( 
.A1(n_2507),
.A2(n_2472),
.B1(n_2400),
.B2(n_2405),
.C(n_2403),
.Y(n_2596)
);

AOI211xp5_ASAP7_75t_L g2597 ( 
.A1(n_2529),
.A2(n_2365),
.B(n_2434),
.C(n_2432),
.Y(n_2597)
);

OAI22xp5_ASAP7_75t_L g2598 ( 
.A1(n_2511),
.A2(n_2442),
.B1(n_2385),
.B2(n_2396),
.Y(n_2598)
);

O2A1O1Ixp33_ASAP7_75t_L g2599 ( 
.A1(n_2519),
.A2(n_2464),
.B(n_2466),
.C(n_2441),
.Y(n_2599)
);

AOI221xp5_ASAP7_75t_L g2600 ( 
.A1(n_2559),
.A2(n_2433),
.B1(n_2429),
.B2(n_2421),
.C(n_2456),
.Y(n_2600)
);

AND4x1_ASAP7_75t_L g2601 ( 
.A(n_2520),
.B(n_2450),
.C(n_2461),
.D(n_2449),
.Y(n_2601)
);

INVxp67_ASAP7_75t_L g2602 ( 
.A(n_2534),
.Y(n_2602)
);

OAI22xp5_ASAP7_75t_L g2603 ( 
.A1(n_2574),
.A2(n_2560),
.B1(n_2568),
.B2(n_2513),
.Y(n_2603)
);

OAI31xp33_ASAP7_75t_L g2604 ( 
.A1(n_2582),
.A2(n_2370),
.A3(n_2455),
.B(n_2411),
.Y(n_2604)
);

NOR3xp33_ASAP7_75t_L g2605 ( 
.A(n_2557),
.B(n_2407),
.C(n_2454),
.Y(n_2605)
);

OAI22xp33_ASAP7_75t_L g2606 ( 
.A1(n_2522),
.A2(n_2435),
.B1(n_2457),
.B2(n_2460),
.Y(n_2606)
);

INVxp67_ASAP7_75t_L g2607 ( 
.A(n_2536),
.Y(n_2607)
);

OAI22xp5_ASAP7_75t_L g2608 ( 
.A1(n_2548),
.A2(n_2467),
.B1(n_2369),
.B2(n_2448),
.Y(n_2608)
);

OAI21xp33_ASAP7_75t_SL g2609 ( 
.A1(n_2514),
.A2(n_2395),
.B(n_2397),
.Y(n_2609)
);

AOI221xp5_ASAP7_75t_L g2610 ( 
.A1(n_2509),
.A2(n_2394),
.B1(n_2443),
.B2(n_2378),
.C(n_2462),
.Y(n_2610)
);

OAI21xp5_ASAP7_75t_L g2611 ( 
.A1(n_2523),
.A2(n_2378),
.B(n_2465),
.Y(n_2611)
);

OAI22xp5_ASAP7_75t_SL g2612 ( 
.A1(n_2528),
.A2(n_2463),
.B1(n_2394),
.B2(n_2500),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2515),
.B(n_2471),
.Y(n_2613)
);

O2A1O1Ixp33_ASAP7_75t_SL g2614 ( 
.A1(n_2527),
.A2(n_2423),
.B(n_154),
.C(n_151),
.Y(n_2614)
);

NAND3xp33_ASAP7_75t_L g2615 ( 
.A(n_2512),
.B(n_2524),
.C(n_2525),
.Y(n_2615)
);

OAI21xp33_ASAP7_75t_L g2616 ( 
.A1(n_2581),
.A2(n_633),
.B(n_630),
.Y(n_2616)
);

OAI21xp5_ASAP7_75t_L g2617 ( 
.A1(n_2570),
.A2(n_1618),
.B(n_153),
.Y(n_2617)
);

AOI21xp33_ASAP7_75t_SL g2618 ( 
.A1(n_2519),
.A2(n_154),
.B(n_155),
.Y(n_2618)
);

OAI211xp5_ASAP7_75t_SL g2619 ( 
.A1(n_2561),
.A2(n_157),
.B(n_155),
.C(n_156),
.Y(n_2619)
);

O2A1O1Ixp33_ASAP7_75t_L g2620 ( 
.A1(n_2594),
.A2(n_159),
.B(n_156),
.C(n_158),
.Y(n_2620)
);

NOR2xp33_ASAP7_75t_L g2621 ( 
.A(n_2577),
.B(n_158),
.Y(n_2621)
);

OAI211xp5_ASAP7_75t_L g2622 ( 
.A1(n_2553),
.A2(n_161),
.B(n_159),
.C(n_160),
.Y(n_2622)
);

OA22x2_ASAP7_75t_L g2623 ( 
.A1(n_2531),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_2623)
);

OAI322xp33_ASAP7_75t_SL g2624 ( 
.A1(n_2572),
.A2(n_164),
.A3(n_165),
.B1(n_166),
.B2(n_167),
.C1(n_168),
.C2(n_170),
.Y(n_2624)
);

NAND3xp33_ASAP7_75t_L g2625 ( 
.A(n_2592),
.B(n_2562),
.C(n_2593),
.Y(n_2625)
);

OAI221xp5_ASAP7_75t_L g2626 ( 
.A1(n_2544),
.A2(n_644),
.B1(n_662),
.B2(n_637),
.C(n_635),
.Y(n_2626)
);

NOR2xp33_ASAP7_75t_L g2627 ( 
.A(n_2577),
.B(n_164),
.Y(n_2627)
);

OAI221xp5_ASAP7_75t_L g2628 ( 
.A1(n_2535),
.A2(n_676),
.B1(n_682),
.B2(n_674),
.C(n_670),
.Y(n_2628)
);

OAI22xp5_ASAP7_75t_L g2629 ( 
.A1(n_2526),
.A2(n_1573),
.B1(n_1558),
.B2(n_1555),
.Y(n_2629)
);

AOI221xp5_ASAP7_75t_L g2630 ( 
.A1(n_2565),
.A2(n_686),
.B1(n_688),
.B2(n_684),
.C(n_683),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_SL g2631 ( 
.A(n_2575),
.B(n_691),
.Y(n_2631)
);

NOR2xp33_ASAP7_75t_L g2632 ( 
.A(n_2518),
.B(n_165),
.Y(n_2632)
);

AND4x1_ASAP7_75t_L g2633 ( 
.A(n_2569),
.B(n_171),
.C(n_166),
.D(n_170),
.Y(n_2633)
);

AOI211xp5_ASAP7_75t_L g2634 ( 
.A1(n_2539),
.A2(n_173),
.B(n_171),
.C(n_172),
.Y(n_2634)
);

CKINVDCx5p33_ASAP7_75t_R g2635 ( 
.A(n_2566),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2576),
.B(n_173),
.Y(n_2636)
);

NOR2xp33_ASAP7_75t_L g2637 ( 
.A(n_2516),
.B(n_174),
.Y(n_2637)
);

OAI221xp5_ASAP7_75t_L g2638 ( 
.A1(n_2510),
.A2(n_713),
.B1(n_734),
.B2(n_708),
.C(n_707),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2556),
.Y(n_2639)
);

AOI311xp33_ASAP7_75t_L g2640 ( 
.A1(n_2542),
.A2(n_176),
.A3(n_174),
.B(n_175),
.C(n_177),
.Y(n_2640)
);

OAI221xp5_ASAP7_75t_L g2641 ( 
.A1(n_2585),
.A2(n_760),
.B1(n_781),
.B2(n_758),
.C(n_755),
.Y(n_2641)
);

XNOR2xp5_ASAP7_75t_L g2642 ( 
.A(n_2586),
.B(n_176),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2530),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2533),
.Y(n_2644)
);

AOI221xp5_ASAP7_75t_L g2645 ( 
.A1(n_2590),
.A2(n_799),
.B1(n_804),
.B2(n_786),
.C(n_785),
.Y(n_2645)
);

AND2x4_ASAP7_75t_L g2646 ( 
.A(n_2517),
.B(n_178),
.Y(n_2646)
);

NOR4xp25_ASAP7_75t_L g2647 ( 
.A(n_2545),
.B(n_184),
.C(n_181),
.D(n_182),
.Y(n_2647)
);

AOI21xp5_ASAP7_75t_L g2648 ( 
.A1(n_2564),
.A2(n_181),
.B(n_184),
.Y(n_2648)
);

OAI21xp5_ASAP7_75t_SL g2649 ( 
.A1(n_2537),
.A2(n_185),
.B(n_186),
.Y(n_2649)
);

AOI22xp33_ASAP7_75t_L g2650 ( 
.A1(n_2552),
.A2(n_1675),
.B1(n_1558),
.B2(n_1573),
.Y(n_2650)
);

AOI211x1_ASAP7_75t_L g2651 ( 
.A1(n_2573),
.A2(n_189),
.B(n_185),
.C(n_188),
.Y(n_2651)
);

OAI211xp5_ASAP7_75t_SL g2652 ( 
.A1(n_2578),
.A2(n_2546),
.B(n_2558),
.C(n_2580),
.Y(n_2652)
);

AOI21xp5_ASAP7_75t_L g2653 ( 
.A1(n_2615),
.A2(n_2541),
.B(n_2571),
.Y(n_2653)
);

AND2x2_ASAP7_75t_L g2654 ( 
.A(n_2640),
.B(n_2543),
.Y(n_2654)
);

OAI211xp5_ASAP7_75t_L g2655 ( 
.A1(n_2604),
.A2(n_2550),
.B(n_2563),
.C(n_2547),
.Y(n_2655)
);

OAI22xp5_ASAP7_75t_L g2656 ( 
.A1(n_2603),
.A2(n_2567),
.B1(n_2583),
.B2(n_2579),
.Y(n_2656)
);

NOR3xp33_ASAP7_75t_L g2657 ( 
.A(n_2652),
.B(n_2554),
.C(n_2588),
.Y(n_2657)
);

AOI22xp5_ASAP7_75t_L g2658 ( 
.A1(n_2595),
.A2(n_2589),
.B1(n_2587),
.B2(n_2521),
.Y(n_2658)
);

OAI321xp33_ASAP7_75t_L g2659 ( 
.A1(n_2611),
.A2(n_2584),
.A3(n_2555),
.B1(n_2532),
.B2(n_2540),
.C(n_2549),
.Y(n_2659)
);

AOI221xp5_ASAP7_75t_L g2660 ( 
.A1(n_2598),
.A2(n_2551),
.B1(n_2591),
.B2(n_2538),
.C(n_823),
.Y(n_2660)
);

XOR2x2_ASAP7_75t_L g2661 ( 
.A(n_2642),
.B(n_189),
.Y(n_2661)
);

OAI211xp5_ASAP7_75t_L g2662 ( 
.A1(n_2600),
.A2(n_192),
.B(n_190),
.C(n_191),
.Y(n_2662)
);

AOI221x1_ASAP7_75t_L g2663 ( 
.A1(n_2605),
.A2(n_193),
.B1(n_190),
.B2(n_192),
.C(n_194),
.Y(n_2663)
);

NOR2xp33_ASAP7_75t_R g2664 ( 
.A(n_2635),
.B(n_195),
.Y(n_2664)
);

AOI221x1_ASAP7_75t_L g2665 ( 
.A1(n_2608),
.A2(n_198),
.B1(n_195),
.B2(n_197),
.C(n_199),
.Y(n_2665)
);

OAI211xp5_ASAP7_75t_SL g2666 ( 
.A1(n_2597),
.A2(n_201),
.B(n_198),
.C(n_199),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2623),
.Y(n_2667)
);

AOI22xp33_ASAP7_75t_L g2668 ( 
.A1(n_2643),
.A2(n_1558),
.B1(n_1573),
.B2(n_1706),
.Y(n_2668)
);

AOI221xp5_ASAP7_75t_L g2669 ( 
.A1(n_2614),
.A2(n_832),
.B1(n_835),
.B2(n_817),
.C(n_814),
.Y(n_2669)
);

AOI22xp5_ASAP7_75t_L g2670 ( 
.A1(n_2602),
.A2(n_2607),
.B1(n_2639),
.B2(n_2644),
.Y(n_2670)
);

OAI221xp5_ASAP7_75t_SL g2671 ( 
.A1(n_2601),
.A2(n_206),
.B1(n_203),
.B2(n_204),
.C(n_208),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_SL g2672 ( 
.A(n_2647),
.B(n_838),
.Y(n_2672)
);

OAI211xp5_ASAP7_75t_L g2673 ( 
.A1(n_2609),
.A2(n_209),
.B(n_204),
.C(n_206),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_L g2674 ( 
.A(n_2651),
.B(n_209),
.Y(n_2674)
);

A2O1A1Ixp33_ASAP7_75t_L g2675 ( 
.A1(n_2621),
.A2(n_212),
.B(n_210),
.C(n_211),
.Y(n_2675)
);

BUFx6f_ASAP7_75t_L g2676 ( 
.A(n_2646),
.Y(n_2676)
);

BUFx2_ASAP7_75t_L g2677 ( 
.A(n_2623),
.Y(n_2677)
);

OAI22xp5_ASAP7_75t_L g2678 ( 
.A1(n_2612),
.A2(n_1540),
.B1(n_1555),
.B2(n_1706),
.Y(n_2678)
);

AOI211xp5_ASAP7_75t_SL g2679 ( 
.A1(n_2606),
.A2(n_2616),
.B(n_2596),
.C(n_2637),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_SL g2680 ( 
.A(n_2610),
.B(n_2618),
.Y(n_2680)
);

AOI22xp5_ASAP7_75t_L g2681 ( 
.A1(n_2627),
.A2(n_1609),
.B1(n_1540),
.B2(n_844),
.Y(n_2681)
);

NOR3xp33_ASAP7_75t_L g2682 ( 
.A(n_2641),
.B(n_849),
.C(n_843),
.Y(n_2682)
);

OAI221xp5_ASAP7_75t_SL g2683 ( 
.A1(n_2599),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.C(n_216),
.Y(n_2683)
);

OAI221xp5_ASAP7_75t_L g2684 ( 
.A1(n_2617),
.A2(n_860),
.B1(n_926),
.B2(n_931),
.C(n_932),
.Y(n_2684)
);

OAI211xp5_ASAP7_75t_SL g2685 ( 
.A1(n_2613),
.A2(n_221),
.B(n_214),
.C(n_220),
.Y(n_2685)
);

AOI21xp5_ASAP7_75t_L g2686 ( 
.A1(n_2624),
.A2(n_220),
.B(n_221),
.Y(n_2686)
);

AOI22xp5_ASAP7_75t_L g2687 ( 
.A1(n_2631),
.A2(n_2625),
.B1(n_2632),
.B2(n_2636),
.Y(n_2687)
);

OAI21xp5_ASAP7_75t_L g2688 ( 
.A1(n_2648),
.A2(n_942),
.B(n_940),
.Y(n_2688)
);

OAI221xp5_ASAP7_75t_L g2689 ( 
.A1(n_2669),
.A2(n_2649),
.B1(n_2620),
.B2(n_2638),
.C(n_2628),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2654),
.B(n_2677),
.Y(n_2690)
);

OAI211xp5_ASAP7_75t_SL g2691 ( 
.A1(n_2670),
.A2(n_2634),
.B(n_2630),
.C(n_2622),
.Y(n_2691)
);

INVx2_ASAP7_75t_SL g2692 ( 
.A(n_2664),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2676),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2676),
.Y(n_2694)
);

AOI21xp33_ASAP7_75t_SL g2695 ( 
.A1(n_2680),
.A2(n_2646),
.B(n_2626),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2667),
.B(n_2633),
.Y(n_2696)
);

OR2x2_ASAP7_75t_L g2697 ( 
.A(n_2674),
.B(n_2650),
.Y(n_2697)
);

INVx1_ASAP7_75t_SL g2698 ( 
.A(n_2661),
.Y(n_2698)
);

INVx2_ASAP7_75t_SL g2699 ( 
.A(n_2676),
.Y(n_2699)
);

AOI22xp33_ASAP7_75t_L g2700 ( 
.A1(n_2672),
.A2(n_2619),
.B1(n_2645),
.B2(n_2629),
.Y(n_2700)
);

AND2x2_ASAP7_75t_L g2701 ( 
.A(n_2657),
.B(n_222),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2665),
.B(n_222),
.Y(n_2702)
);

OAI32xp33_ASAP7_75t_L g2703 ( 
.A1(n_2685),
.A2(n_223),
.A3(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_2703)
);

INVx3_ASAP7_75t_L g2704 ( 
.A(n_2671),
.Y(n_2704)
);

OR2x2_ASAP7_75t_L g2705 ( 
.A(n_2683),
.B(n_223),
.Y(n_2705)
);

OAI22xp5_ASAP7_75t_L g2706 ( 
.A1(n_2684),
.A2(n_950),
.B1(n_1555),
.B2(n_1711),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2663),
.Y(n_2707)
);

AOI21xp5_ASAP7_75t_L g2708 ( 
.A1(n_2686),
.A2(n_224),
.B(n_227),
.Y(n_2708)
);

AOI221xp5_ASAP7_75t_L g2709 ( 
.A1(n_2707),
.A2(n_2656),
.B1(n_2653),
.B2(n_2660),
.C(n_2673),
.Y(n_2709)
);

NAND5xp2_ASAP7_75t_L g2710 ( 
.A(n_2708),
.B(n_2679),
.C(n_2655),
.D(n_2687),
.E(n_2658),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2699),
.B(n_2675),
.Y(n_2711)
);

AOI221xp5_ASAP7_75t_L g2712 ( 
.A1(n_2690),
.A2(n_2659),
.B1(n_2682),
.B2(n_2688),
.C(n_2666),
.Y(n_2712)
);

OAI211xp5_ASAP7_75t_SL g2713 ( 
.A1(n_2694),
.A2(n_2662),
.B(n_2681),
.C(n_2668),
.Y(n_2713)
);

CKINVDCx5p33_ASAP7_75t_R g2714 ( 
.A(n_2692),
.Y(n_2714)
);

CKINVDCx20_ASAP7_75t_R g2715 ( 
.A(n_2698),
.Y(n_2715)
);

NOR2x1_ASAP7_75t_L g2716 ( 
.A(n_2693),
.B(n_2678),
.Y(n_2716)
);

NAND3xp33_ASAP7_75t_L g2717 ( 
.A(n_2695),
.B(n_227),
.C(n_228),
.Y(n_2717)
);

NOR2x1_ASAP7_75t_L g2718 ( 
.A(n_2705),
.B(n_228),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2702),
.Y(n_2719)
);

AO22x2_ASAP7_75t_L g2720 ( 
.A1(n_2701),
.A2(n_235),
.B1(n_229),
.B2(n_234),
.Y(n_2720)
);

NAND4xp25_ASAP7_75t_L g2721 ( 
.A(n_2696),
.B(n_239),
.C(n_234),
.D(n_236),
.Y(n_2721)
);

NOR3xp33_ASAP7_75t_L g2722 ( 
.A(n_2691),
.B(n_236),
.C(n_240),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2704),
.B(n_240),
.Y(n_2723)
);

NOR3xp33_ASAP7_75t_L g2724 ( 
.A(n_2689),
.B(n_241),
.C(n_242),
.Y(n_2724)
);

AND2x2_ASAP7_75t_L g2725 ( 
.A(n_2700),
.B(n_242),
.Y(n_2725)
);

HB1xp67_ASAP7_75t_L g2726 ( 
.A(n_2720),
.Y(n_2726)
);

NOR2x1_ASAP7_75t_L g2727 ( 
.A(n_2715),
.B(n_2697),
.Y(n_2727)
);

CKINVDCx20_ASAP7_75t_R g2728 ( 
.A(n_2714),
.Y(n_2728)
);

BUFx6f_ASAP7_75t_L g2729 ( 
.A(n_2719),
.Y(n_2729)
);

CKINVDCx5p33_ASAP7_75t_R g2730 ( 
.A(n_2723),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_2722),
.B(n_2703),
.Y(n_2731)
);

INVxp67_ASAP7_75t_L g2732 ( 
.A(n_2710),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2720),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2725),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2711),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2718),
.Y(n_2736)
);

CKINVDCx5p33_ASAP7_75t_R g2737 ( 
.A(n_2717),
.Y(n_2737)
);

NAND2xp33_ASAP7_75t_R g2738 ( 
.A(n_2709),
.B(n_243),
.Y(n_2738)
);

CKINVDCx5p33_ASAP7_75t_R g2739 ( 
.A(n_2712),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2724),
.B(n_2706),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2716),
.Y(n_2741)
);

CKINVDCx5p33_ASAP7_75t_R g2742 ( 
.A(n_2721),
.Y(n_2742)
);

INVx1_ASAP7_75t_SL g2743 ( 
.A(n_2713),
.Y(n_2743)
);

CKINVDCx20_ASAP7_75t_R g2744 ( 
.A(n_2715),
.Y(n_2744)
);

OAI22x1_ASAP7_75t_L g2745 ( 
.A1(n_2741),
.A2(n_247),
.B1(n_244),
.B2(n_245),
.Y(n_2745)
);

HB1xp67_ASAP7_75t_L g2746 ( 
.A(n_2744),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2728),
.Y(n_2747)
);

OR2x2_ASAP7_75t_L g2748 ( 
.A(n_2732),
.B(n_247),
.Y(n_2748)
);

OA22x2_ASAP7_75t_L g2749 ( 
.A1(n_2743),
.A2(n_256),
.B1(n_250),
.B2(n_255),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2727),
.Y(n_2750)
);

CKINVDCx20_ASAP7_75t_R g2751 ( 
.A(n_2730),
.Y(n_2751)
);

AOI21xp5_ASAP7_75t_L g2752 ( 
.A1(n_2726),
.A2(n_258),
.B(n_259),
.Y(n_2752)
);

XNOR2x1_ASAP7_75t_L g2753 ( 
.A(n_2739),
.B(n_259),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2736),
.B(n_260),
.Y(n_2754)
);

AOI21xp5_ASAP7_75t_L g2755 ( 
.A1(n_2729),
.A2(n_260),
.B(n_262),
.Y(n_2755)
);

OAI22xp5_ASAP7_75t_L g2756 ( 
.A1(n_2729),
.A2(n_1609),
.B1(n_265),
.B2(n_263),
.Y(n_2756)
);

NOR2xp67_ASAP7_75t_L g2757 ( 
.A(n_2729),
.B(n_264),
.Y(n_2757)
);

AO22x2_ASAP7_75t_L g2758 ( 
.A1(n_2733),
.A2(n_267),
.B1(n_264),
.B2(n_266),
.Y(n_2758)
);

INVx1_ASAP7_75t_SL g2759 ( 
.A(n_2731),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_2735),
.Y(n_2760)
);

NOR2x1_ASAP7_75t_L g2761 ( 
.A(n_2734),
.B(n_268),
.Y(n_2761)
);

AOI22x1_ASAP7_75t_L g2762 ( 
.A1(n_2742),
.A2(n_2737),
.B1(n_2738),
.B2(n_2740),
.Y(n_2762)
);

AOI22xp5_ASAP7_75t_L g2763 ( 
.A1(n_2744),
.A2(n_1609),
.B1(n_272),
.B2(n_268),
.Y(n_2763)
);

OAI22xp5_ASAP7_75t_L g2764 ( 
.A1(n_2744),
.A2(n_274),
.B1(n_269),
.B2(n_273),
.Y(n_2764)
);

AOI22xp5_ASAP7_75t_L g2765 ( 
.A1(n_2750),
.A2(n_2746),
.B1(n_2751),
.B2(n_2747),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2758),
.Y(n_2766)
);

OAI22xp5_ASAP7_75t_L g2767 ( 
.A1(n_2759),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_2767)
);

OR2x6_ASAP7_75t_L g2768 ( 
.A(n_2760),
.B(n_275),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_2758),
.Y(n_2769)
);

AOI22xp33_ASAP7_75t_L g2770 ( 
.A1(n_2762),
.A2(n_2761),
.B1(n_2753),
.B2(n_2749),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2757),
.Y(n_2771)
);

OAI22xp33_ASAP7_75t_L g2772 ( 
.A1(n_2748),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.Y(n_2772)
);

OA22x2_ASAP7_75t_L g2773 ( 
.A1(n_2745),
.A2(n_280),
.B1(n_277),
.B2(n_278),
.Y(n_2773)
);

AOI22xp5_ASAP7_75t_L g2774 ( 
.A1(n_2763),
.A2(n_2754),
.B1(n_2756),
.B2(n_2764),
.Y(n_2774)
);

NOR2xp33_ASAP7_75t_L g2775 ( 
.A(n_2752),
.B(n_2755),
.Y(n_2775)
);

CKINVDCx20_ASAP7_75t_R g2776 ( 
.A(n_2746),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2746),
.Y(n_2777)
);

CKINVDCx20_ASAP7_75t_R g2778 ( 
.A(n_2746),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_SL g2779 ( 
.A(n_2746),
.B(n_280),
.Y(n_2779)
);

BUFx2_ASAP7_75t_L g2780 ( 
.A(n_2776),
.Y(n_2780)
);

HB1xp67_ASAP7_75t_L g2781 ( 
.A(n_2778),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2777),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2765),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2766),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2769),
.Y(n_2785)
);

INVx1_ASAP7_75t_SL g2786 ( 
.A(n_2768),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2768),
.Y(n_2787)
);

INVxp67_ASAP7_75t_L g2788 ( 
.A(n_2779),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2773),
.Y(n_2789)
);

HB1xp67_ASAP7_75t_L g2790 ( 
.A(n_2771),
.Y(n_2790)
);

HB1xp67_ASAP7_75t_L g2791 ( 
.A(n_2767),
.Y(n_2791)
);

INVx8_ASAP7_75t_L g2792 ( 
.A(n_2770),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2775),
.Y(n_2793)
);

OAI22xp5_ASAP7_75t_L g2794 ( 
.A1(n_2781),
.A2(n_2774),
.B1(n_2772),
.B2(n_283),
.Y(n_2794)
);

AOI21xp5_ASAP7_75t_L g2795 ( 
.A1(n_2780),
.A2(n_281),
.B(n_282),
.Y(n_2795)
);

OAI22x1_ASAP7_75t_L g2796 ( 
.A1(n_2783),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_2796)
);

AOI22xp5_ASAP7_75t_L g2797 ( 
.A1(n_2782),
.A2(n_289),
.B1(n_284),
.B2(n_288),
.Y(n_2797)
);

OAI22xp5_ASAP7_75t_L g2798 ( 
.A1(n_2793),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2792),
.B(n_291),
.Y(n_2799)
);

AND2x2_ASAP7_75t_L g2800 ( 
.A(n_2786),
.B(n_292),
.Y(n_2800)
);

OAI22xp5_ASAP7_75t_L g2801 ( 
.A1(n_2784),
.A2(n_293),
.B1(n_295),
.B2(n_298),
.Y(n_2801)
);

AOI21xp5_ASAP7_75t_L g2802 ( 
.A1(n_2792),
.A2(n_293),
.B(n_295),
.Y(n_2802)
);

NOR4xp25_ASAP7_75t_L g2803 ( 
.A(n_2785),
.B(n_298),
.C(n_299),
.D(n_300),
.Y(n_2803)
);

OAI22xp5_ASAP7_75t_L g2804 ( 
.A1(n_2789),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_2804)
);

CKINVDCx20_ASAP7_75t_R g2805 ( 
.A(n_2790),
.Y(n_2805)
);

CKINVDCx20_ASAP7_75t_R g2806 ( 
.A(n_2791),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2787),
.Y(n_2807)
);

XNOR2x1_ASAP7_75t_L g2808 ( 
.A(n_2788),
.B(n_301),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2805),
.B(n_302),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2806),
.Y(n_2810)
);

AOI21xp5_ASAP7_75t_L g2811 ( 
.A1(n_2799),
.A2(n_303),
.B(n_304),
.Y(n_2811)
);

AOI22xp5_ASAP7_75t_L g2812 ( 
.A1(n_2807),
.A2(n_303),
.B1(n_305),
.B2(n_306),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_SL g2813 ( 
.A(n_2803),
.B(n_307),
.Y(n_2813)
);

AOI22xp5_ASAP7_75t_L g2814 ( 
.A1(n_2808),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2800),
.Y(n_2815)
);

XNOR2xp5_ASAP7_75t_L g2816 ( 
.A(n_2794),
.B(n_309),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2796),
.Y(n_2817)
);

OAI22xp5_ASAP7_75t_L g2818 ( 
.A1(n_2797),
.A2(n_2802),
.B1(n_2795),
.B2(n_2804),
.Y(n_2818)
);

INVx1_ASAP7_75t_SL g2819 ( 
.A(n_2801),
.Y(n_2819)
);

NAND2xp33_ASAP7_75t_L g2820 ( 
.A(n_2798),
.B(n_310),
.Y(n_2820)
);

OAI22xp5_ASAP7_75t_L g2821 ( 
.A1(n_2810),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_2821)
);

XNOR2xp5_ASAP7_75t_L g2822 ( 
.A(n_2815),
.B(n_313),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2809),
.Y(n_2823)
);

INVx5_ASAP7_75t_L g2824 ( 
.A(n_2817),
.Y(n_2824)
);

OAI221xp5_ASAP7_75t_L g2825 ( 
.A1(n_2814),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.C(n_317),
.Y(n_2825)
);

OAI22xp5_ASAP7_75t_L g2826 ( 
.A1(n_2819),
.A2(n_317),
.B1(n_318),
.B2(n_321),
.Y(n_2826)
);

OAI221xp5_ASAP7_75t_L g2827 ( 
.A1(n_2816),
.A2(n_321),
.B1(n_325),
.B2(n_326),
.C(n_327),
.Y(n_2827)
);

AOI221x1_ASAP7_75t_L g2828 ( 
.A1(n_2818),
.A2(n_325),
.B1(n_329),
.B2(n_330),
.C(n_331),
.Y(n_2828)
);

OAI222xp33_ASAP7_75t_L g2829 ( 
.A1(n_2813),
.A2(n_2811),
.B1(n_2812),
.B2(n_2820),
.C1(n_337),
.C2(n_338),
.Y(n_2829)
);

OAI22xp5_ASAP7_75t_L g2830 ( 
.A1(n_2810),
.A2(n_332),
.B1(n_335),
.B2(n_336),
.Y(n_2830)
);

XNOR2x1_ASAP7_75t_L g2831 ( 
.A(n_2810),
.B(n_332),
.Y(n_2831)
);

AOI22xp33_ASAP7_75t_L g2832 ( 
.A1(n_2824),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_2832)
);

AOI22xp33_ASAP7_75t_SL g2833 ( 
.A1(n_2824),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.Y(n_2833)
);

OR2x2_ASAP7_75t_L g2834 ( 
.A(n_2823),
.B(n_340),
.Y(n_2834)
);

OAI22xp5_ASAP7_75t_SL g2835 ( 
.A1(n_2822),
.A2(n_341),
.B1(n_344),
.B2(n_346),
.Y(n_2835)
);

AOI221x1_ASAP7_75t_L g2836 ( 
.A1(n_2826),
.A2(n_346),
.B1(n_347),
.B2(n_348),
.C(n_350),
.Y(n_2836)
);

AOI222xp33_ASAP7_75t_L g2837 ( 
.A1(n_2829),
.A2(n_347),
.B1(n_348),
.B2(n_350),
.C1(n_351),
.C2(n_352),
.Y(n_2837)
);

AO21x1_ASAP7_75t_L g2838 ( 
.A1(n_2831),
.A2(n_352),
.B(n_353),
.Y(n_2838)
);

AOI222xp33_ASAP7_75t_L g2839 ( 
.A1(n_2825),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.C1(n_356),
.C2(n_357),
.Y(n_2839)
);

OAI221xp5_ASAP7_75t_L g2840 ( 
.A1(n_2827),
.A2(n_2830),
.B1(n_2821),
.B2(n_2828),
.C(n_357),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2824),
.Y(n_2841)
);

AOI22xp5_ASAP7_75t_L g2842 ( 
.A1(n_2841),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_2842)
);

AOI22xp33_ASAP7_75t_L g2843 ( 
.A1(n_2838),
.A2(n_358),
.B1(n_359),
.B2(n_360),
.Y(n_2843)
);

AOI22xp5_ASAP7_75t_L g2844 ( 
.A1(n_2835),
.A2(n_358),
.B1(n_362),
.B2(n_1553),
.Y(n_2844)
);

AOI22xp5_ASAP7_75t_L g2845 ( 
.A1(n_2837),
.A2(n_362),
.B1(n_1553),
.B2(n_367),
.Y(n_2845)
);

AOI22x1_ASAP7_75t_L g2846 ( 
.A1(n_2843),
.A2(n_2839),
.B1(n_2834),
.B2(n_2836),
.Y(n_2846)
);

OR2x2_ASAP7_75t_L g2847 ( 
.A(n_2844),
.B(n_2832),
.Y(n_2847)
);

AOI221xp5_ASAP7_75t_L g2848 ( 
.A1(n_2847),
.A2(n_2840),
.B1(n_2845),
.B2(n_2833),
.C(n_2842),
.Y(n_2848)
);

AOI211xp5_ASAP7_75t_L g2849 ( 
.A1(n_2848),
.A2(n_2846),
.B(n_368),
.C(n_369),
.Y(n_2849)
);


endmodule