module fake_jpeg_30707_n_536 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_536);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_536;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_53),
.B(n_55),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_56),
.Y(n_148)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_29),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_59),
.B(n_64),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_60),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_30),
.B(n_0),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_21),
.B(n_1),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_90),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_36),
.B(n_49),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_79),
.B(n_27),
.C(n_50),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_21),
.B(n_1),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_1),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_94),
.Y(n_124)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_45),
.B(n_34),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_19),
.B(n_2),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_99),
.B(n_20),
.Y(n_107)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_105),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_107),
.B(n_118),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_77),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_110),
.B(n_42),
.Y(n_206)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_56),
.A2(n_52),
.B1(n_38),
.B2(n_40),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_115),
.A2(n_126),
.B1(n_147),
.B2(n_156),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_66),
.A2(n_40),
.B1(n_38),
.B2(n_26),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_129),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_132),
.B(n_136),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_SL g136 ( 
.A1(n_64),
.A2(n_44),
.B(n_28),
.Y(n_136)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_101),
.A2(n_60),
.B1(n_103),
.B2(n_54),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_62),
.Y(n_153)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_59),
.A2(n_40),
.B1(n_38),
.B2(n_28),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_78),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_159),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_53),
.A2(n_43),
.B1(n_50),
.B2(n_47),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_163),
.A2(n_156),
.B1(n_138),
.B2(n_144),
.Y(n_195)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_79),
.Y(n_164)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_108),
.B(n_99),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_169),
.B(n_171),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_106),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_172),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_173),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_174),
.Y(n_234)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_175),
.Y(n_264)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_176),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_124),
.B(n_27),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_177),
.B(n_180),
.Y(n_245)
);

AO22x1_ASAP7_75t_SL g178 ( 
.A1(n_130),
.A2(n_70),
.B1(n_71),
.B2(n_87),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_178),
.A2(n_189),
.B1(n_126),
.B2(n_115),
.Y(n_243)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_47),
.Y(n_180)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_111),
.B(n_2),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_182),
.B(n_159),
.C(n_140),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_165),
.A2(n_89),
.B1(n_100),
.B2(n_105),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_183),
.A2(n_222),
.B1(n_170),
.B2(n_212),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_143),
.A2(n_43),
.B(n_34),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_184),
.Y(n_246)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_119),
.Y(n_185)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_185),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_55),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_186),
.B(n_198),
.Y(n_260)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_121),
.Y(n_187)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_187),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_109),
.A2(n_96),
.B1(n_44),
.B2(n_42),
.Y(n_189)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_191),
.Y(n_252)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_112),
.Y(n_192)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_192),
.Y(n_254)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_194),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_212),
.Y(n_242)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_125),
.Y(n_197)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_116),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_201),
.Y(n_267)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_203),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_139),
.B(n_42),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_204),
.B(n_205),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_117),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_206),
.B(n_209),
.Y(n_251)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_141),
.Y(n_207)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_207),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_208),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_134),
.B(n_42),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_123),
.Y(n_210)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_210),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_142),
.B(n_44),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_133),
.Y(n_213)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_213),
.Y(n_269)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_120),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_214),
.B(n_216),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_117),
.A2(n_96),
.B1(n_44),
.B2(n_4),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_215),
.A2(n_221),
.B1(n_225),
.B2(n_226),
.Y(n_248)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_137),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_149),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_217),
.B(n_218),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_153),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_158),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_219),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_160),
.A2(n_31),
.B1(n_51),
.B2(n_4),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_220),
.B(n_31),
.Y(n_275)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_114),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_151),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_223),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_166),
.B(n_31),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_224),
.Y(n_273)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_152),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_140),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_114),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_227),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_229),
.B(n_7),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_145),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_232),
.B(n_256),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_188),
.B(n_5),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_235),
.B(n_253),
.Y(n_276)
);

NAND2xp33_ASAP7_75t_SL g237 ( 
.A(n_181),
.B(n_178),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_237),
.A2(n_176),
.B(n_215),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_243),
.A2(n_249),
.B1(n_271),
.B2(n_173),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_190),
.A2(n_147),
.B1(n_148),
.B2(n_145),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_193),
.B(n_6),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_211),
.B(n_135),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_263),
.Y(n_285)
);

OR2x4_ASAP7_75t_L g263 ( 
.A(n_184),
.B(n_6),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_182),
.B(n_135),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_221),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_196),
.A2(n_148),
.B1(n_183),
.B2(n_223),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_274),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_275),
.Y(n_278)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_277),
.Y(n_319)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_279),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_217),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_280),
.B(n_284),
.Y(n_341)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_228),
.Y(n_281)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_281),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_232),
.B(n_168),
.C(n_197),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_282),
.B(n_283),
.C(n_293),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_189),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_245),
.B(n_210),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_273),
.A2(n_202),
.B1(n_226),
.B2(n_203),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_286),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_245),
.B(n_175),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_287),
.B(n_291),
.Y(n_342)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_228),
.Y(n_288)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_288),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_273),
.A2(n_179),
.B1(n_214),
.B2(n_191),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_289),
.A2(n_258),
.B(n_252),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_290),
.A2(n_311),
.B1(n_313),
.B2(n_268),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_187),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_242),
.B(n_185),
.C(n_208),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_255),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_294),
.B(n_295),
.Y(n_346)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_272),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_296),
.B(n_302),
.Y(n_325)
);

AO21x1_ASAP7_75t_L g349 ( 
.A1(n_297),
.A2(n_241),
.B(n_252),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_242),
.A2(n_227),
.B1(n_174),
.B2(n_51),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_298),
.A2(n_249),
.B1(n_243),
.B2(n_250),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_239),
.B(n_172),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_299),
.B(n_300),
.Y(n_351)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_231),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_265),
.B(n_6),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_231),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_303),
.B(n_304),
.Y(n_332)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_233),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_233),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_305),
.Y(n_320)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_254),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_306),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_242),
.A2(n_51),
.B1(n_172),
.B2(n_9),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_307),
.A2(n_259),
.B1(n_248),
.B2(n_275),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_240),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_308),
.Y(n_348)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_254),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_309),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_239),
.B(n_31),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_310),
.B(n_314),
.Y(n_333)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_261),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_312),
.B(n_264),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_238),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_246),
.B(n_7),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_270),
.B(n_8),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_316),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_270),
.B(n_8),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_266),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_317),
.A2(n_250),
.B1(n_238),
.B2(n_267),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_323),
.A2(n_331),
.B1(n_336),
.B2(n_337),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_326),
.A2(n_318),
.B(n_351),
.Y(n_382)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_327),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_328),
.A2(n_340),
.B1(n_345),
.B2(n_288),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_292),
.B(n_312),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_330),
.B(n_240),
.C(n_308),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_290),
.A2(n_237),
.B1(n_275),
.B2(n_251),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_297),
.A2(n_278),
.B(n_285),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_334),
.A2(n_339),
.B(n_317),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_292),
.A2(n_229),
.B1(n_263),
.B2(n_268),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_285),
.A2(n_258),
.B1(n_234),
.B2(n_235),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_278),
.A2(n_262),
.B(n_230),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_298),
.A2(n_269),
.B1(n_262),
.B2(n_253),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_285),
.A2(n_293),
.B1(n_296),
.B2(n_295),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_343),
.A2(n_352),
.B1(n_281),
.B2(n_236),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_344),
.A2(n_349),
.B(n_355),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_283),
.A2(n_269),
.B1(n_230),
.B2(n_257),
.Y(n_345)
);

XOR2x2_ASAP7_75t_SL g347 ( 
.A(n_282),
.B(n_257),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_347),
.B(n_350),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_301),
.A2(n_234),
.B1(n_240),
.B2(n_261),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_302),
.B(n_264),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_353),
.B(n_307),
.Y(n_357)
);

AO21x1_ASAP7_75t_L g355 ( 
.A1(n_315),
.A2(n_241),
.B(n_244),
.Y(n_355)
);

NAND3xp33_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_276),
.C(n_316),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_360),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_357),
.B(n_335),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_358),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_324),
.B(n_277),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_323),
.B(n_294),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_361),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_341),
.B(n_300),
.Y(n_362)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_362),
.Y(n_391)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_363),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_341),
.B(n_304),
.Y(n_364)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_364),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_334),
.A2(n_301),
.B(n_305),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_365),
.B(n_373),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_342),
.B(n_303),
.Y(n_366)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_366),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_346),
.B(n_279),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_368),
.B(n_369),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_346),
.B(n_244),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_330),
.B(n_311),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_370),
.B(n_384),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_332),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_383),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_372),
.A2(n_343),
.B1(n_337),
.B2(n_347),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_342),
.B(n_309),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_319),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_380),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_375),
.A2(n_388),
.B1(n_340),
.B2(n_328),
.Y(n_409)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_319),
.Y(n_376)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_376),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_326),
.B(n_236),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_377),
.A2(n_382),
.B(n_389),
.Y(n_417)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_329),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_378),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_325),
.B(n_306),
.Y(n_380)
);

OAI21xp33_ASAP7_75t_SL g381 ( 
.A1(n_339),
.A2(n_247),
.B(n_234),
.Y(n_381)
);

OAI21xp33_ASAP7_75t_SL g402 ( 
.A1(n_381),
.A2(n_349),
.B(n_344),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_351),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_329),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_386),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_325),
.B(n_308),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_331),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_347),
.A2(n_17),
.B(n_11),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_390),
.B(n_401),
.Y(n_436)
);

OA21x2_ASAP7_75t_L g396 ( 
.A1(n_379),
.A2(n_358),
.B(n_359),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_396),
.B(n_409),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_400),
.A2(n_410),
.B1(n_412),
.B2(n_367),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_387),
.B(n_350),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_402),
.A2(n_365),
.B(n_377),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_383),
.B(n_333),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_403),
.B(n_411),
.Y(n_421)
);

MAJx2_ASAP7_75t_L g404 ( 
.A(n_361),
.B(n_335),
.C(n_336),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_404),
.B(n_357),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_361),
.A2(n_349),
.B1(n_352),
.B2(n_353),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_373),
.B(n_324),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_372),
.A2(n_379),
.B1(n_359),
.B2(n_377),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_362),
.B(n_320),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_414),
.B(n_376),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_371),
.A2(n_345),
.B1(n_320),
.B2(n_354),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_418),
.B(n_420),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_367),
.A2(n_354),
.B1(n_348),
.B2(n_355),
.Y(n_419)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_419),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_364),
.B(n_321),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_394),
.B(n_370),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_422),
.B(n_430),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_423),
.A2(n_419),
.B1(n_409),
.B2(n_418),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_399),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_437),
.Y(n_448)
);

INVx13_ASAP7_75t_L g427 ( 
.A(n_406),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_427),
.B(n_435),
.Y(n_455)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_420),
.Y(n_428)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_428),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_394),
.B(n_387),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_431),
.B(n_440),
.C(n_441),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g432 ( 
.A1(n_391),
.A2(n_382),
.B1(n_407),
.B2(n_397),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_432),
.A2(n_434),
.B1(n_398),
.B2(n_396),
.Y(n_462)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_415),
.Y(n_433)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_433),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_413),
.A2(n_363),
.B1(n_389),
.B2(n_375),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_392),
.B(n_366),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_391),
.B(n_380),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_438),
.A2(n_442),
.B1(n_410),
.B2(n_395),
.Y(n_456)
);

OA21x2_ASAP7_75t_SL g439 ( 
.A1(n_405),
.A2(n_413),
.B(n_404),
.Y(n_439)
);

MAJx2_ASAP7_75t_L g460 ( 
.A(n_439),
.B(n_428),
.C(n_446),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_390),
.B(n_384),
.C(n_386),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_397),
.B(n_388),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_416),
.B(n_355),
.Y(n_443)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_443),
.Y(n_449)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_415),
.Y(n_444)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_444),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_407),
.B(n_374),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_445),
.Y(n_468)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_408),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_446),
.B(n_408),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_447),
.B(n_456),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_443),
.A2(n_405),
.B(n_416),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_451),
.A2(n_453),
.B(n_429),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_443),
.A2(n_412),
.B(n_417),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_441),
.B(n_400),
.C(n_401),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_440),
.C(n_431),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_425),
.A2(n_417),
.B1(n_395),
.B2(n_393),
.Y(n_459)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_459),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_460),
.Y(n_472)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_461),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_462),
.B(n_434),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_424),
.A2(n_396),
.B1(n_406),
.B2(n_398),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_463),
.B(n_464),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_424),
.A2(n_385),
.B1(n_378),
.B2(n_348),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_423),
.A2(n_322),
.B1(n_321),
.B2(n_338),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_465),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_430),
.A2(n_322),
.B1(n_338),
.B2(n_12),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_466),
.B(n_442),
.Y(n_481)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_469),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_479),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_471),
.B(n_480),
.Y(n_492)
);

INVxp33_ASAP7_75t_L g473 ( 
.A(n_455),
.Y(n_473)
);

INVx13_ASAP7_75t_L g498 ( 
.A(n_473),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_450),
.B(n_422),
.C(n_436),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_475),
.B(n_452),
.C(n_460),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_451),
.A2(n_429),
.B(n_426),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_477),
.A2(n_453),
.B(n_449),
.Y(n_490)
);

MAJx2_ASAP7_75t_L g479 ( 
.A(n_457),
.B(n_439),
.C(n_436),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_452),
.B(n_450),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_481),
.B(n_483),
.Y(n_493)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_458),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_448),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_485),
.A2(n_468),
.B1(n_454),
.B2(n_449),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_474),
.A2(n_448),
.B1(n_447),
.B2(n_463),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_487),
.B(n_488),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_489),
.B(n_495),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_490),
.B(n_494),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_480),
.B(n_462),
.C(n_465),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_491),
.B(n_478),
.C(n_472),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_471),
.B(n_426),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_SL g495 ( 
.A(n_479),
.B(n_427),
.C(n_421),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_470),
.B(n_464),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_496),
.B(n_500),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_482),
.B(n_445),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_473),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_475),
.B(n_466),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_497),
.A2(n_482),
.B1(n_472),
.B2(n_478),
.Y(n_505)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_505),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_509),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_507),
.B(n_508),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_491),
.A2(n_484),
.B1(n_468),
.B2(n_476),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_499),
.A2(n_458),
.B1(n_477),
.B2(n_467),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_493),
.A2(n_484),
.B1(n_438),
.B2(n_444),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_510),
.A2(n_512),
.B(n_509),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_498),
.B(n_469),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_511),
.B(n_494),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_492),
.B(n_433),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_515),
.A2(n_517),
.B1(n_520),
.B2(n_512),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_516),
.B(n_504),
.Y(n_522)
);

NOR2x1_ASAP7_75t_L g517 ( 
.A(n_505),
.B(n_486),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_501),
.A2(n_489),
.B(n_486),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_518),
.A2(n_503),
.B(n_496),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_SL g520 ( 
.A1(n_508),
.A2(n_498),
.B1(n_427),
.B2(n_500),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_521),
.B(n_522),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_523),
.A2(n_525),
.B(n_514),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_519),
.B(n_513),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_524),
.B(n_503),
.C(n_502),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_513),
.B(n_506),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_526),
.B(n_527),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_528),
.A2(n_521),
.B(n_492),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_530),
.B(n_10),
.C(n_11),
.Y(n_531)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_531),
.A2(n_529),
.B(n_12),
.Y(n_532)
);

AOI221xp5_ASAP7_75t_L g533 ( 
.A1(n_532),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.C(n_16),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_SL g534 ( 
.A1(n_533),
.A2(n_16),
.B1(n_10),
.B2(n_13),
.Y(n_534)
);

BUFx24_ASAP7_75t_SL g535 ( 
.A(n_534),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_13),
.Y(n_536)
);


endmodule