module fake_ariane_2242_n_756 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_756);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_756;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_670;
wire n_607;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_677;
wire n_614;
wire n_604;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_658;
wire n_705;
wire n_630;
wire n_616;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_697;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

INVx1_ASAP7_75t_L g154 ( 
.A(n_63),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_84),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_53),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_114),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_7),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_26),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_98),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_57),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_152),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_7),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_61),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_68),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_133),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_1),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_36),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_56),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_100),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_151),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_43),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_9),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_23),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_137),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_97),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_139),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_49),
.B(n_150),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_71),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_30),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_42),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_27),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_9),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_25),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_8),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_83),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_10),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_122),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_96),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_87),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_69),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_112),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_11),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_70),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_58),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_44),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_143),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_62),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_117),
.Y(n_206)
);

CKINVDCx6p67_ASAP7_75t_R g207 ( 
.A(n_167),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_183),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_174),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

OA21x2_ASAP7_75t_L g211 ( 
.A1(n_154),
.A2(n_0),
.B(n_1),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_155),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_0),
.Y(n_214)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

AND2x6_ASAP7_75t_L g221 ( 
.A(n_171),
.B(n_21),
.Y(n_221)
);

AND2x6_ASAP7_75t_L g222 ( 
.A(n_171),
.B(n_22),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_158),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_165),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_187),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_160),
.B(n_2),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_2),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_161),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_166),
.Y(n_229)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_176),
.B(n_3),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_169),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_178),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_186),
.Y(n_233)
);

AOI22x1_ASAP7_75t_SL g234 ( 
.A1(n_191),
.A2(n_198),
.B1(n_195),
.B2(n_196),
.Y(n_234)
);

OAI21x1_ASAP7_75t_L g235 ( 
.A1(n_188),
.A2(n_79),
.B(n_147),
.Y(n_235)
);

AND2x2_ASAP7_75t_SL g236 ( 
.A(n_182),
.B(n_24),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

OAI22x1_ASAP7_75t_SL g238 ( 
.A1(n_179),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g239 ( 
.A(n_156),
.Y(n_239)
);

AND2x4_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_4),
.Y(n_240)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_171),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_203),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_171),
.Y(n_246)
);

BUFx6f_ASAP7_75t_SL g247 ( 
.A(n_236),
.Y(n_247)
);

AOI21x1_ASAP7_75t_L g248 ( 
.A1(n_233),
.A2(n_204),
.B(n_180),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_209),
.B(n_193),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_209),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_208),
.B(n_216),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_208),
.B(n_157),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_215),
.Y(n_258)
);

OR2x6_ASAP7_75t_L g259 ( 
.A(n_214),
.B(n_210),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_217),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_213),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_212),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_220),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_213),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_220),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_217),
.B(n_159),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_228),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_215),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_228),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_236),
.B(n_162),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_227),
.A2(n_206),
.B1(n_201),
.B2(n_164),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_246),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_210),
.B(n_168),
.Y(n_275)
);

NOR2x1p5_ASAP7_75t_L g276 ( 
.A(n_207),
.B(n_170),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_231),
.B(n_224),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_232),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_233),
.B(n_244),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_243),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_244),
.B(n_172),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_243),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_237),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_243),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_224),
.B(n_173),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_237),
.Y(n_287)
);

INVx8_ASAP7_75t_L g288 ( 
.A(n_221),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_236),
.B(n_177),
.Y(n_289)
);

NAND2xp33_ASAP7_75t_SL g290 ( 
.A(n_230),
.B(n_184),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_245),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_230),
.Y(n_292)
);

NOR2x1p5_ASAP7_75t_L g293 ( 
.A(n_207),
.B(n_181),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

NOR3xp33_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_226),
.C(n_240),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_254),
.B(n_239),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_286),
.B(n_239),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_252),
.B(n_230),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_252),
.B(n_230),
.Y(n_299)
);

AOI221xp5_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_238),
.B1(n_277),
.B2(n_260),
.C(n_227),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_263),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_252),
.B(n_240),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_240),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_240),
.Y(n_305)
);

NOR3xp33_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_227),
.C(n_225),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_245),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_263),
.B(n_242),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_287),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_265),
.B(n_242),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_254),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_288),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_247),
.A2(n_197),
.B1(n_211),
.B2(n_225),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_267),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_267),
.B(n_273),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_287),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_275),
.B(n_229),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_273),
.B(n_242),
.Y(n_319)
);

AOI221xp5_ASAP7_75t_L g320 ( 
.A1(n_290),
.A2(n_219),
.B1(n_229),
.B2(n_223),
.C(n_185),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_274),
.B(n_219),
.Y(n_321)
);

A2O1A1Ixp33_ASAP7_75t_L g322 ( 
.A1(n_279),
.A2(n_235),
.B(n_223),
.C(n_190),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g323 ( 
.A(n_266),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_274),
.B(n_215),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_250),
.B(n_223),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_257),
.B(n_215),
.Y(n_326)
);

O2A1O1Ixp33_ASAP7_75t_L g327 ( 
.A1(n_255),
.A2(n_211),
.B(n_6),
.C(n_8),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_279),
.B(n_215),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_281),
.B(n_215),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_272),
.B(n_280),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_259),
.B(n_211),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_280),
.B(n_180),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_291),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_282),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_282),
.B(n_218),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_291),
.B(n_218),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_261),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_261),
.B(n_180),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_264),
.B(n_218),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_264),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_259),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_247),
.A2(n_211),
.B1(n_234),
.B2(n_235),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_268),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_268),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_259),
.B(n_221),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_L g346 ( 
.A1(n_259),
.A2(n_234),
.B1(n_180),
.B2(n_204),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_270),
.B(n_218),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_270),
.B(n_218),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_278),
.B(n_204),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_278),
.B(n_218),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_293),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_283),
.B(n_241),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_283),
.B(n_241),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_284),
.B(n_241),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_284),
.B(n_241),
.Y(n_355)
);

NAND2xp33_ASAP7_75t_L g356 ( 
.A(n_288),
.B(n_221),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_288),
.B(n_204),
.Y(n_357)
);

OAI21xp33_ASAP7_75t_L g358 ( 
.A1(n_304),
.A2(n_247),
.B(n_248),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_305),
.A2(n_253),
.B(n_251),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_298),
.A2(n_302),
.B(n_299),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_323),
.B(n_293),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_328),
.A2(n_251),
.B(n_249),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_316),
.A2(n_253),
.B(n_249),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_344),
.B(n_276),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_329),
.A2(n_307),
.B(n_324),
.Y(n_365)
);

BUFx4f_ASAP7_75t_SL g366 ( 
.A(n_318),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_301),
.A2(n_315),
.B(n_314),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_321),
.Y(n_368)
);

NOR3xp33_ASAP7_75t_L g369 ( 
.A(n_300),
.B(n_256),
.C(n_262),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_294),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_309),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_308),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_296),
.B(n_5),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_344),
.B(n_256),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_320),
.B(n_241),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_311),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_317),
.Y(n_377)
);

OAI21xp33_ASAP7_75t_L g378 ( 
.A1(n_295),
.A2(n_248),
.B(n_262),
.Y(n_378)
);

BUFx4f_ASAP7_75t_L g379 ( 
.A(n_345),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_335),
.A2(n_258),
.B(n_269),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_306),
.B(n_258),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_306),
.B(n_221),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_356),
.A2(n_269),
.B(n_241),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_345),
.B(n_269),
.Y(n_384)
);

O2A1O1Ixp33_ASAP7_75t_L g385 ( 
.A1(n_295),
.A2(n_6),
.B(n_10),
.C(n_11),
.Y(n_385)
);

OAI21xp33_ASAP7_75t_L g386 ( 
.A1(n_343),
.A2(n_12),
.B(n_13),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_333),
.B(n_221),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_322),
.A2(n_222),
.B(n_221),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_341),
.B(n_221),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_303),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_331),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_330),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_334),
.A2(n_222),
.B(n_269),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_333),
.A2(n_269),
.B(n_222),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_310),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_347),
.A2(n_222),
.B(n_86),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_327),
.A2(n_222),
.B(n_85),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_319),
.Y(n_398)
);

AOI21xp33_ASAP7_75t_L g399 ( 
.A1(n_313),
.A2(n_12),
.B(n_13),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_346),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_337),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_340),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_303),
.B(n_14),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_348),
.A2(n_222),
.B(n_89),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_325),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_332),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_350),
.A2(n_222),
.B(n_88),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_297),
.B(n_14),
.Y(n_408)
);

NOR2x1_ASAP7_75t_L g409 ( 
.A(n_346),
.B(n_28),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_351),
.B(n_15),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_342),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_326),
.B(n_15),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_303),
.B(n_16),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_338),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_303),
.B(n_16),
.Y(n_415)
);

OAI21x1_ASAP7_75t_L g416 ( 
.A1(n_352),
.A2(n_91),
.B(n_146),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_353),
.A2(n_90),
.B(n_145),
.Y(n_417)
);

AOI21xp33_ASAP7_75t_L g418 ( 
.A1(n_339),
.A2(n_17),
.B(n_18),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_312),
.B(n_17),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_355),
.A2(n_92),
.B(n_142),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_357),
.A2(n_18),
.B(n_19),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_349),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_336),
.A2(n_19),
.B(n_20),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_354),
.A2(n_20),
.B(n_29),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_379),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_411),
.A2(n_354),
.B1(n_339),
.B2(n_312),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_402),
.Y(n_427)
);

OAI21xp33_ASAP7_75t_L g428 ( 
.A1(n_373),
.A2(n_312),
.B(n_32),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_360),
.A2(n_312),
.B(n_33),
.Y(n_429)
);

OAI21x1_ASAP7_75t_L g430 ( 
.A1(n_365),
.A2(n_31),
.B(n_34),
.Y(n_430)
);

OAI21x1_ASAP7_75t_L g431 ( 
.A1(n_393),
.A2(n_35),
.B(n_37),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_360),
.A2(n_38),
.B(n_39),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_387),
.A2(n_374),
.B(n_367),
.Y(n_433)
);

OAI21x1_ASAP7_75t_L g434 ( 
.A1(n_362),
.A2(n_40),
.B(n_41),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_392),
.Y(n_435)
);

BUFx4f_ASAP7_75t_L g436 ( 
.A(n_389),
.Y(n_436)
);

NAND2x1_ASAP7_75t_L g437 ( 
.A(n_390),
.B(n_45),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_390),
.A2(n_46),
.B(n_47),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_359),
.A2(n_48),
.B(n_50),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_359),
.A2(n_51),
.B(n_52),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_400),
.B(n_54),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_391),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_370),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_379),
.B(n_55),
.Y(n_444)
);

CKINVDCx14_ASAP7_75t_R g445 ( 
.A(n_408),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_399),
.A2(n_409),
.B1(n_368),
.B2(n_401),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_372),
.A2(n_59),
.B(n_60),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_395),
.B(n_64),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_371),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_405),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_398),
.B(n_65),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_376),
.Y(n_452)
);

NAND2x1p5_ASAP7_75t_L g453 ( 
.A(n_384),
.B(n_66),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_413),
.A2(n_67),
.B(n_72),
.Y(n_454)
);

OAI21x1_ASAP7_75t_L g455 ( 
.A1(n_362),
.A2(n_388),
.B(n_363),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_L g456 ( 
.A(n_390),
.B(n_73),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_397),
.A2(n_74),
.B(n_75),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_369),
.B(n_76),
.Y(n_458)
);

AO221x1_ASAP7_75t_L g459 ( 
.A1(n_377),
.A2(n_77),
.B1(n_80),
.B2(n_81),
.C(n_82),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_364),
.B(n_361),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_410),
.B(n_93),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_366),
.Y(n_462)
);

AOI21x1_ASAP7_75t_L g463 ( 
.A1(n_394),
.A2(n_382),
.B(n_363),
.Y(n_463)
);

AOI221xp5_ASAP7_75t_SL g464 ( 
.A1(n_385),
.A2(n_94),
.B1(n_95),
.B2(n_99),
.C(n_101),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_419),
.A2(n_102),
.B(n_103),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_389),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_377),
.B(n_104),
.Y(n_467)
);

OAI21x1_ASAP7_75t_L g468 ( 
.A1(n_380),
.A2(n_105),
.B(n_106),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_386),
.A2(n_412),
.B1(n_403),
.B2(n_415),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_406),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_381),
.A2(n_107),
.B(n_108),
.Y(n_471)
);

OAI21x1_ASAP7_75t_SL g472 ( 
.A1(n_424),
.A2(n_111),
.B(n_113),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_414),
.B(n_115),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_422),
.Y(n_474)
);

OA21x2_ASAP7_75t_L g475 ( 
.A1(n_358),
.A2(n_118),
.B(n_119),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_375),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_378),
.B(n_124),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_383),
.A2(n_125),
.B(n_126),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_416),
.Y(n_479)
);

OAI21x1_ASAP7_75t_L g480 ( 
.A1(n_396),
.A2(n_127),
.B(n_128),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_427),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_425),
.Y(n_482)
);

NAND2x1p5_ASAP7_75t_L g483 ( 
.A(n_436),
.B(n_421),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_424),
.Y(n_484)
);

BUFx8_ASAP7_75t_L g485 ( 
.A(n_452),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_474),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_425),
.B(n_421),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_443),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_463),
.A2(n_407),
.B(n_404),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_470),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_455),
.A2(n_420),
.B(n_417),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_425),
.B(n_423),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_SL g493 ( 
.A1(n_445),
.A2(n_441),
.B1(n_457),
.B2(n_459),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_466),
.B(n_423),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_442),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_449),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_462),
.Y(n_497)
);

BUFx5_ASAP7_75t_L g498 ( 
.A(n_479),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_462),
.Y(n_499)
);

BUFx2_ASAP7_75t_SL g500 ( 
.A(n_444),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_433),
.A2(n_418),
.B(n_130),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_435),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_436),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_450),
.B(n_148),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_457),
.A2(n_134),
.B(n_135),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_460),
.B(n_136),
.Y(n_506)
);

O2A1O1Ixp33_ASAP7_75t_L g507 ( 
.A1(n_469),
.A2(n_138),
.B(n_140),
.C(n_141),
.Y(n_507)
);

OAI21x1_ASAP7_75t_SL g508 ( 
.A1(n_472),
.A2(n_458),
.B(n_448),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_448),
.Y(n_509)
);

BUFx4f_ASAP7_75t_L g510 ( 
.A(n_453),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_429),
.A2(n_428),
.B(n_469),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_451),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_451),
.Y(n_513)
);

AO21x2_ASAP7_75t_L g514 ( 
.A1(n_477),
.A2(n_467),
.B(n_461),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_430),
.A2(n_431),
.B(n_434),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_446),
.B(n_473),
.Y(n_516)
);

AO21x2_ASAP7_75t_L g517 ( 
.A1(n_477),
.A2(n_467),
.B(n_432),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_468),
.A2(n_480),
.B(n_440),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_439),
.A2(n_471),
.B(n_465),
.Y(n_519)
);

OA21x2_ASAP7_75t_L g520 ( 
.A1(n_464),
.A2(n_454),
.B(n_447),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_426),
.B(n_453),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_456),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_464),
.A2(n_476),
.B1(n_437),
.B2(n_475),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_478),
.A2(n_475),
.B(n_438),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_488),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_481),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_494),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_486),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_494),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_506),
.B(n_490),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_484),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_493),
.A2(n_506),
.B1(n_512),
.B2(n_495),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_515),
.A2(n_524),
.B(n_518),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_484),
.Y(n_534)
);

INVxp33_ASAP7_75t_L g535 ( 
.A(n_497),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_498),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_513),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_498),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_487),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_483),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_495),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_509),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_498),
.Y(n_543)
);

BUFx2_ASAP7_75t_SL g544 ( 
.A(n_482),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_498),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_521),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_493),
.A2(n_516),
.B1(n_496),
.B2(n_505),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_521),
.Y(n_548)
);

BUFx8_ASAP7_75t_SL g549 ( 
.A(n_502),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_498),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_485),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_492),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_492),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_501),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_487),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_483),
.Y(n_556)
);

BUFx2_ASAP7_75t_R g557 ( 
.A(n_500),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_485),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_482),
.B(n_522),
.Y(n_559)
);

AOI21x1_ASAP7_75t_L g560 ( 
.A1(n_511),
.A2(n_508),
.B(n_491),
.Y(n_560)
);

CKINVDCx11_ASAP7_75t_R g561 ( 
.A(n_499),
.Y(n_561)
);

INVx8_ASAP7_75t_L g562 ( 
.A(n_504),
.Y(n_562)
);

AO21x1_ASAP7_75t_SL g563 ( 
.A1(n_505),
.A2(n_523),
.B(n_507),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_489),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_542),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_539),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_546),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_546),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_542),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_548),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_548),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_527),
.B(n_511),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_527),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_539),
.B(n_552),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_529),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_529),
.Y(n_576)
);

BUFx2_ASAP7_75t_SL g577 ( 
.A(n_559),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_549),
.B(n_510),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_539),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_541),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_535),
.B(n_510),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_552),
.B(n_514),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_553),
.B(n_514),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_532),
.A2(n_517),
.B1(n_520),
.B2(n_503),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_530),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_553),
.B(n_507),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_555),
.B(n_528),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_530),
.B(n_520),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_526),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_526),
.B(n_517),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_531),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_528),
.B(n_519),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_537),
.B(n_531),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_534),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_534),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_554),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_537),
.B(n_556),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_556),
.B(n_532),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_564),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_554),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_525),
.B(n_540),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_525),
.B(n_540),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_547),
.B(n_540),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_562),
.B(n_559),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_536),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_540),
.B(n_563),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_564),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_562),
.A2(n_557),
.B1(n_559),
.B2(n_558),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_566),
.Y(n_609)
);

NAND3xp33_ASAP7_75t_SL g610 ( 
.A(n_578),
.B(n_551),
.C(n_561),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_596),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_565),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_566),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_597),
.B(n_545),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_596),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_565),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_597),
.B(n_545),
.Y(n_617)
);

AND2x4_ASAP7_75t_SL g618 ( 
.A(n_566),
.B(n_559),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_580),
.B(n_585),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_600),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_593),
.B(n_562),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_600),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_569),
.B(n_545),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_579),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_606),
.B(n_543),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_569),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_SL g627 ( 
.A1(n_598),
.A2(n_562),
.B1(n_563),
.B2(n_558),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_574),
.B(n_543),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_575),
.B(n_562),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_606),
.B(n_543),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_574),
.B(n_536),
.Y(n_631)
);

NAND2x1p5_ASAP7_75t_SL g632 ( 
.A(n_586),
.B(n_538),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_570),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_570),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_590),
.B(n_538),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_SL g636 ( 
.A1(n_598),
.A2(n_544),
.B1(n_550),
.B2(n_533),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_566),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_567),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_590),
.B(n_550),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_579),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_567),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_568),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_573),
.B(n_560),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_592),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_573),
.B(n_560),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_619),
.B(n_571),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_614),
.B(n_577),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_644),
.B(n_588),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_644),
.B(n_573),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_612),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_614),
.B(n_571),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_617),
.B(n_568),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_617),
.B(n_592),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_635),
.B(n_602),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_628),
.B(n_586),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_627),
.A2(n_603),
.B1(n_584),
.B2(n_608),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_609),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_635),
.B(n_601),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_639),
.B(n_601),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_640),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_638),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_638),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_621),
.B(n_581),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_639),
.B(n_602),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_624),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_628),
.B(n_582),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_631),
.B(n_582),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_631),
.B(n_625),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_610),
.A2(n_603),
.B1(n_595),
.B2(n_594),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_625),
.B(n_630),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_625),
.B(n_566),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_641),
.B(n_595),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_668),
.B(n_640),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_670),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_655),
.B(n_632),
.Y(n_675)
);

NOR2x1_ASAP7_75t_L g676 ( 
.A(n_663),
.B(n_609),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_661),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_660),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_662),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_663),
.B(n_609),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_669),
.B(n_636),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_655),
.B(n_632),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_665),
.B(n_641),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_670),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_651),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_668),
.B(n_625),
.Y(n_686)
);

NOR2xp67_ASAP7_75t_L g687 ( 
.A(n_674),
.B(n_670),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_677),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_681),
.A2(n_669),
.B1(n_656),
.B2(n_630),
.Y(n_689)
);

AOI32xp33_ASAP7_75t_L g690 ( 
.A1(n_681),
.A2(n_656),
.A3(n_646),
.B1(n_647),
.B2(n_653),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_675),
.B(n_652),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_682),
.B(n_653),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_678),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_679),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_680),
.B(n_666),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_683),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_694),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_688),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_L g699 ( 
.A1(n_689),
.A2(n_676),
.B1(n_674),
.B2(n_684),
.Y(n_699)
);

AO22x1_ASAP7_75t_L g700 ( 
.A1(n_696),
.A2(n_674),
.B1(n_684),
.B2(n_685),
.Y(n_700)
);

XNOR2x1_ASAP7_75t_L g701 ( 
.A(n_690),
.B(n_686),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_698),
.Y(n_702)
);

NAND4xp25_ASAP7_75t_SL g703 ( 
.A(n_701),
.B(n_695),
.C(n_692),
.D(n_691),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_697),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_700),
.B(n_693),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_699),
.Y(n_706)
);

OAI221xp5_ASAP7_75t_L g707 ( 
.A1(n_701),
.A2(n_687),
.B1(n_672),
.B2(n_649),
.C(n_648),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_702),
.Y(n_708)
);

NOR4xp25_ASAP7_75t_L g709 ( 
.A(n_703),
.B(n_673),
.C(n_629),
.D(n_642),
.Y(n_709)
);

AOI31xp33_ASAP7_75t_L g710 ( 
.A1(n_705),
.A2(n_673),
.A3(n_686),
.B(n_604),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_704),
.B(n_642),
.Y(n_711)
);

AOI211xp5_ASAP7_75t_L g712 ( 
.A1(n_709),
.A2(n_706),
.B(n_707),
.C(n_620),
.Y(n_712)
);

NOR2x1_ASAP7_75t_L g713 ( 
.A(n_708),
.B(n_544),
.Y(n_713)
);

NOR3xp33_ASAP7_75t_L g714 ( 
.A(n_710),
.B(n_657),
.C(n_611),
.Y(n_714)
);

NOR3x1_ASAP7_75t_L g715 ( 
.A(n_712),
.B(n_711),
.C(n_620),
.Y(n_715)
);

NAND4xp75_ASAP7_75t_L g716 ( 
.A(n_713),
.B(n_667),
.C(n_666),
.D(n_589),
.Y(n_716)
);

OAI221xp5_ASAP7_75t_L g717 ( 
.A1(n_714),
.A2(n_591),
.B1(n_594),
.B2(n_575),
.C(n_576),
.Y(n_717)
);

NOR3xp33_ASAP7_75t_L g718 ( 
.A(n_712),
.B(n_591),
.C(n_576),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_718),
.A2(n_671),
.B1(n_637),
.B2(n_613),
.Y(n_719)
);

NOR3x2_ASAP7_75t_L g720 ( 
.A(n_716),
.B(n_572),
.C(n_657),
.Y(n_720)
);

NAND4xp75_ASAP7_75t_L g721 ( 
.A(n_715),
.B(n_667),
.C(n_589),
.D(n_615),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_717),
.A2(n_671),
.B1(n_637),
.B2(n_613),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_716),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_718),
.A2(n_622),
.B(n_615),
.Y(n_724)
);

NOR2x1_ASAP7_75t_L g725 ( 
.A(n_716),
.B(n_657),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_723),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_724),
.B(n_622),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_721),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_719),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_720),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_722),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_725),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_726),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_730),
.B(n_630),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_732),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_728),
.A2(n_671),
.B1(n_630),
.B2(n_577),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_728),
.A2(n_611),
.B1(n_645),
.B2(n_643),
.Y(n_737)
);

AO22x2_ASAP7_75t_L g738 ( 
.A1(n_729),
.A2(n_634),
.B1(n_664),
.B2(n_659),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_727),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_739),
.Y(n_740)
);

OAI31xp33_ASAP7_75t_L g741 ( 
.A1(n_733),
.A2(n_731),
.A3(n_572),
.B(n_618),
.Y(n_741)
);

AOI21xp33_ASAP7_75t_L g742 ( 
.A1(n_735),
.A2(n_634),
.B(n_605),
.Y(n_742)
);

OA22x2_ASAP7_75t_L g743 ( 
.A1(n_734),
.A2(n_618),
.B1(n_645),
.B2(n_643),
.Y(n_743)
);

AOI22x1_ASAP7_75t_L g744 ( 
.A1(n_738),
.A2(n_737),
.B1(n_736),
.B2(n_623),
.Y(n_744)
);

OAI21xp5_ASAP7_75t_SL g745 ( 
.A1(n_740),
.A2(n_623),
.B(n_587),
.Y(n_745)
);

OAI21xp33_ASAP7_75t_L g746 ( 
.A1(n_743),
.A2(n_742),
.B(n_744),
.Y(n_746)
);

OAI22x1_ASAP7_75t_L g747 ( 
.A1(n_741),
.A2(n_658),
.B1(n_654),
.B2(n_650),
.Y(n_747)
);

OAI22xp33_ASAP7_75t_SL g748 ( 
.A1(n_740),
.A2(n_605),
.B1(n_650),
.B2(n_626),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_746),
.B(n_626),
.Y(n_749)
);

OAI21xp5_ASAP7_75t_L g750 ( 
.A1(n_745),
.A2(n_533),
.B(n_583),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_748),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_749),
.A2(n_747),
.B1(n_587),
.B2(n_583),
.Y(n_752)
);

OAI21xp5_ASAP7_75t_SL g753 ( 
.A1(n_751),
.A2(n_633),
.B(n_612),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_753),
.A2(n_750),
.B(n_599),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_754),
.B(n_752),
.C(n_616),
.Y(n_755)
);

AOI211xp5_ASAP7_75t_L g756 ( 
.A1(n_755),
.A2(n_616),
.B(n_633),
.C(n_607),
.Y(n_756)
);


endmodule