module fake_jpeg_31193_n_366 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_366);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_366;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_1),
.B(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_6),
.B(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_62),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_7),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_19),
.A2(n_7),
.B(n_13),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_63),
.B(n_13),
.Y(n_118)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_68),
.Y(n_80)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_69),
.Y(n_119)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_71),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_27),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_73),
.Y(n_82)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_76),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_75),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_33),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_37),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_84),
.B(n_87),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_37),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_35),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_38),
.B1(n_39),
.B2(n_27),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_88),
.A2(n_89),
.B1(n_94),
.B2(n_97),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_39),
.B1(n_38),
.B2(n_18),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_35),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_93),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_54),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_92),
.B(n_107),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_18),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_73),
.A2(n_38),
.B1(n_39),
.B2(n_27),
.Y(n_94)
);

AO21x1_ASAP7_75t_L g144 ( 
.A1(n_96),
.A2(n_118),
.B(n_124),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_66),
.A2(n_28),
.B1(n_39),
.B2(n_41),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_46),
.B(n_29),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_28),
.B1(n_25),
.B2(n_41),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_105),
.A2(n_106),
.B1(n_32),
.B2(n_43),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_58),
.A2(n_27),
.B1(n_25),
.B2(n_41),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_45),
.B(n_34),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_34),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_110),
.B(n_6),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_47),
.B(n_29),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_120),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_50),
.A2(n_28),
.B1(n_25),
.B2(n_20),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_117),
.A2(n_43),
.B1(n_26),
.B2(n_32),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_52),
.B(n_29),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_72),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_125),
.Y(n_172)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_126),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_61),
.B1(n_60),
.B2(n_56),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_129),
.Y(n_201)
);

O2A1O1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_101),
.A2(n_55),
.B(n_49),
.C(n_43),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_131),
.A2(n_145),
.B(n_162),
.Y(n_188)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_132),
.Y(n_181)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_86),
.A2(n_76),
.B1(n_26),
.B2(n_42),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_137),
.A2(n_158),
.B1(n_95),
.B2(n_83),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_42),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_147),
.Y(n_168)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_140),
.Y(n_192)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_141),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_155),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_112),
.A2(n_42),
.B1(n_36),
.B2(n_20),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_143),
.A2(n_149),
.B(n_153),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_120),
.A2(n_36),
.B(n_43),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_146),
.B(n_150),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_79),
.B(n_36),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_79),
.B(n_43),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_161),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_43),
.B1(n_33),
.B2(n_26),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_98),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_151),
.B(n_164),
.Y(n_200)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_157),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_159),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_82),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_163),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_0),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_96),
.A2(n_32),
.B(n_7),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_99),
.A2(n_111),
.B1(n_90),
.B2(n_113),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_124),
.B1(n_92),
.B2(n_83),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_166),
.B(n_14),
.Y(n_189)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_80),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_167),
.B(n_81),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_169),
.B(n_170),
.Y(n_208)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_127),
.A2(n_134),
.A3(n_161),
.B1(n_138),
.B2(n_147),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_174),
.A2(n_196),
.B1(n_130),
.B2(n_131),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_127),
.B(n_134),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_177),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_81),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_176),
.B(n_178),
.C(n_184),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_119),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_118),
.C(n_119),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_119),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_182),
.B(n_183),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_145),
.B(n_108),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_164),
.B(n_108),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_187),
.B(n_199),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_194),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_159),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_131),
.A2(n_109),
.B1(n_90),
.B2(n_89),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_153),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_144),
.B(n_152),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_153),
.B(n_109),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_202),
.B(n_205),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_78),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_206),
.A2(n_226),
.B1(n_232),
.B2(n_205),
.Y(n_253)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_203),
.Y(n_207)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_209),
.Y(n_245)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_210),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_128),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_212),
.B(n_216),
.Y(n_259)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_215),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_217),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_218),
.A2(n_201),
.B1(n_174),
.B2(n_204),
.Y(n_241)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_219),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_146),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_220),
.A2(n_229),
.B(n_171),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_136),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_222),
.Y(n_246)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_169),
.B(n_140),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_230),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_188),
.A2(n_141),
.B(n_133),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_225),
.A2(n_198),
.B(n_194),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_196),
.A2(n_139),
.B1(n_125),
.B2(n_132),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_231),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_182),
.B(n_156),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_154),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_168),
.B(n_14),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_188),
.A2(n_116),
.B1(n_102),
.B2(n_85),
.Y(n_232)
);

OAI31xp33_ASAP7_75t_L g233 ( 
.A1(n_199),
.A2(n_155),
.A3(n_113),
.B(n_111),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_233),
.A2(n_187),
.B(n_202),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_176),
.B(n_142),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_237),
.Y(n_262)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_180),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_236),
.Y(n_265)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_191),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_191),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_195),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_178),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_241),
.A2(n_266),
.B1(n_242),
.B2(n_269),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_218),
.A2(n_201),
.B1(n_204),
.B2(n_184),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_242),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_175),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_243),
.B(n_249),
.C(n_251),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_211),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_247),
.B(n_250),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_183),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_214),
.C(n_208),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_253),
.A2(n_229),
.B1(n_210),
.B2(n_213),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_214),
.B(n_168),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_258),
.B(n_219),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_233),
.Y(n_260)
);

NOR2xp67_ASAP7_75t_R g278 ( 
.A(n_260),
.B(n_261),
.Y(n_278)
);

AO22x1_ASAP7_75t_L g261 ( 
.A1(n_218),
.A2(n_197),
.B1(n_170),
.B2(n_171),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_263),
.A2(n_269),
.B(n_225),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_267),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_78),
.B1(n_116),
.B2(n_102),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_189),
.Y(n_267)
);

OAI32xp33_ASAP7_75t_L g270 ( 
.A1(n_227),
.A2(n_173),
.A3(n_181),
.B1(n_172),
.B2(n_98),
.Y(n_270)
);

OAI321xp33_ASAP7_75t_L g277 ( 
.A1(n_270),
.A2(n_229),
.A3(n_220),
.B1(n_173),
.B2(n_222),
.C(n_217),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_239),
.Y(n_273)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_273),
.Y(n_303)
);

AOI321xp33_ASAP7_75t_L g275 ( 
.A1(n_261),
.A2(n_227),
.A3(n_238),
.B1(n_220),
.B2(n_231),
.C(n_206),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_247),
.A2(n_226),
.B1(n_216),
.B2(n_232),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_276),
.A2(n_281),
.B1(n_294),
.B2(n_256),
.Y(n_310)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_277),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_215),
.Y(n_279)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_279),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_280),
.B(n_287),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_292),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_243),
.B(n_209),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_288),
.C(n_251),
.Y(n_295)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_286),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_237),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_249),
.B(n_207),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_265),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_290),
.Y(n_299)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_246),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_291),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_236),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_235),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_252),
.C(n_256),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_241),
.A2(n_228),
.B1(n_78),
.B2(n_85),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_295),
.B(n_311),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_258),
.C(n_263),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_298),
.B(n_300),
.C(n_301),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_250),
.C(n_253),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_259),
.C(n_268),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_244),
.C(n_245),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_312),
.C(n_313),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_282),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_310),
.A2(n_290),
.B1(n_294),
.B2(n_254),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_266),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_271),
.B(n_245),
.C(n_244),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_271),
.B(n_254),
.C(n_255),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_289),
.Y(n_314)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_314),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_304),
.A2(n_278),
.B1(n_300),
.B2(n_296),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_315),
.A2(n_328),
.B1(n_309),
.B2(n_295),
.Y(n_331)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_307),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_317),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_306),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_296),
.A2(n_278),
.B(n_277),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_318),
.B(n_320),
.Y(n_333)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_297),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_319),
.B(n_321),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_286),
.Y(n_321)
);

NAND3xp33_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_274),
.C(n_273),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_327),
.Y(n_334)
);

AOI21x1_ASAP7_75t_SL g324 ( 
.A1(n_311),
.A2(n_272),
.B(n_275),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_324),
.A2(n_314),
.B(n_321),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_280),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_14),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_302),
.B(n_255),
.Y(n_327)
);

AOI21x1_ASAP7_75t_L g343 ( 
.A1(n_330),
.A2(n_324),
.B(n_319),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_338),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_329),
.B(n_181),
.C(n_172),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_332),
.B(n_335),
.C(n_339),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_6),
.C(n_12),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_12),
.C(n_10),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_322),
.B(n_8),
.C(n_10),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_337),
.B(n_318),
.Y(n_342)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_342),
.Y(n_350)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_343),
.Y(n_355)
);

NAND4xp25_ASAP7_75t_SL g344 ( 
.A(n_336),
.B(n_0),
.C(n_1),
.D(n_2),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_338),
.B(n_326),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_334),
.A2(n_326),
.B(n_1),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_347),
.A2(n_2),
.B(n_3),
.Y(n_356)
);

NOR2xp67_ASAP7_75t_L g349 ( 
.A(n_333),
.B(n_330),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_349),
.A2(n_339),
.B1(n_341),
.B2(n_335),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_342),
.A2(n_340),
.B(n_332),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_351),
.A2(n_354),
.B(n_353),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_352),
.B(n_356),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_345),
.B(n_1),
.C(n_2),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_346),
.B(n_348),
.C(n_344),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_350),
.A2(n_348),
.B1(n_346),
.B2(n_5),
.Y(n_357)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_357),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_359),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_351),
.A2(n_334),
.B(n_355),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_362),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_363),
.B(n_364),
.Y(n_365)
);

NAND2x1_ASAP7_75t_SL g364 ( 
.A(n_361),
.B(n_360),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_365),
.B(n_358),
.Y(n_366)
);


endmodule