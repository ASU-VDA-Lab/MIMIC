module fake_jpeg_3742_n_271 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_271);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_271;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_33),
.B1(n_32),
.B2(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_16),
.B(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_20),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_14),
.B(n_0),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_14),
.C(n_30),
.Y(n_80)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_52),
.B(n_54),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_58),
.Y(n_103)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_57),
.Y(n_122)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

CKINVDCx6p67_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_35),
.Y(n_64)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_33),
.B1(n_16),
.B2(n_17),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_67),
.A2(n_95),
.B1(n_21),
.B2(n_8),
.Y(n_121)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_46),
.B(n_31),
.Y(n_72)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_48),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_80),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_15),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_75),
.A2(n_28),
.B(n_21),
.C(n_18),
.Y(n_104)
);

INVx5_ASAP7_75t_SL g76 ( 
.A(n_38),
.Y(n_76)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_45),
.B(n_31),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_83),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_22),
.B1(n_20),
.B2(n_19),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_79),
.A2(n_84),
.B1(n_13),
.B2(n_12),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_40),
.A2(n_25),
.B1(n_22),
.B2(n_19),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_47),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_86),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx5_ASAP7_75t_SL g87 ( 
.A(n_36),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_88),
.Y(n_117)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_89),
.A2(n_93),
.B1(n_94),
.B2(n_99),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_91),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_46),
.A2(n_25),
.B1(n_29),
.B2(n_32),
.Y(n_95)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_104),
.B(n_87),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_84),
.A2(n_29),
.B1(n_24),
.B2(n_23),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_111),
.A2(n_125),
.B1(n_13),
.B2(n_12),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_L g115 ( 
.A1(n_76),
.A2(n_21),
.B1(n_18),
.B2(n_24),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_123),
.B1(n_97),
.B2(n_93),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_53),
.A2(n_23),
.B1(n_15),
.B2(n_18),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_116),
.A2(n_98),
.B1(n_51),
.B2(n_65),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_110),
.B1(n_112),
.B2(n_103),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_64),
.A2(n_60),
.B1(n_92),
.B2(n_96),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_121),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_134),
.C(n_122),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_75),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_128),
.B(n_133),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_129),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_130),
.A2(n_132),
.B1(n_155),
.B2(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_56),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_60),
.C(n_57),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_105),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_135),
.B(n_147),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_92),
.B1(n_98),
.B2(n_51),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_136),
.A2(n_139),
.B1(n_145),
.B2(n_154),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_65),
.B1(n_62),
.B2(n_81),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_137),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_61),
.Y(n_138)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_81),
.Y(n_142)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_144),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_63),
.Y(n_146)
);

NOR2x1_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_7),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_21),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_112),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_151),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_77),
.Y(n_149)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_21),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_SL g161 ( 
.A1(n_150),
.A2(n_152),
.B(n_126),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_107),
.B(n_63),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_0),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_114),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_5),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_123),
.A2(n_77),
.B1(n_82),
.B2(n_59),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_100),
.A2(n_59),
.B1(n_86),
.B2(n_83),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_113),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_118),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

HAxp5_ASAP7_75t_SL g159 ( 
.A(n_146),
.B(n_120),
.CON(n_159),
.SN(n_159)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_161),
.A2(n_184),
.B1(n_170),
.B2(n_163),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_136),
.Y(n_205)
);

AO22x1_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_91),
.B1(n_113),
.B2(n_2),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_163),
.A2(n_170),
.B1(n_178),
.B2(n_129),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_114),
.C(n_126),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_127),
.C(n_134),
.Y(n_196)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_11),
.Y(n_168)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_153),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_174),
.Y(n_191)
);

AO22x1_ASAP7_75t_SL g170 ( 
.A1(n_135),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_155),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_154),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_130),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_144),
.Y(n_197)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_188),
.Y(n_195)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_132),
.B1(n_148),
.B2(n_131),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_204),
.B1(n_187),
.B2(n_175),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_206),
.B1(n_179),
.B2(n_159),
.Y(n_220)
);

A2O1A1Ixp33_ASAP7_75t_SL g226 ( 
.A1(n_194),
.A2(n_208),
.B(n_160),
.C(n_185),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_165),
.C(n_173),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_182),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_147),
.Y(n_198)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_198),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_183),
.A2(n_147),
.B(n_150),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_201),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_150),
.Y(n_200)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_183),
.A2(n_152),
.B(n_137),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_141),
.Y(n_203)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_172),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_163),
.B(n_162),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_152),
.Y(n_207)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

XNOR2x2_ASAP7_75t_SL g208 ( 
.A(n_181),
.B(n_145),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_156),
.Y(n_209)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_177),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_211),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_213),
.C(n_218),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_164),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

NAND4xp25_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_207),
.C(n_194),
.D(n_201),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_216),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_173),
.C(n_169),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_220),
.A2(n_223),
.B1(n_190),
.B2(n_208),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_208),
.A2(n_166),
.B1(n_171),
.B2(n_172),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_205),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_200),
.C(n_199),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_225),
.A2(n_226),
.B(n_198),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_232),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_227),
.B(n_195),
.Y(n_229)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_233),
.A2(n_235),
.B(n_236),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_223),
.A2(n_191),
.B1(n_204),
.B2(n_192),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_237),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_226),
.A2(n_195),
.B(n_202),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_189),
.B(n_197),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_221),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_244),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_189),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_213),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_228),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_235),
.A2(n_210),
.B1(n_217),
.B2(n_222),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_248),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_238),
.B(n_234),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_250),
.C(n_255),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_231),
.C(n_218),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_231),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_224),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_219),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_212),
.C(n_237),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_246),
.A2(n_238),
.B1(n_215),
.B2(n_230),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_256),
.A2(n_226),
.B1(n_247),
.B2(n_233),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_249),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_248),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_260),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_262),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_230),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_254),
.A2(n_243),
.B1(n_246),
.B2(n_226),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_259),
.B(n_243),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_265),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_263),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_268),
.A2(n_266),
.B(n_264),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_270),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_261),
.Y(n_270)
);


endmodule