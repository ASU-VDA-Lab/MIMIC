module real_jpeg_31684_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_0),
.Y(n_138)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_0),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_0),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_1),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_1),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_1),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_1),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_1),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_1),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_1),
.B(n_333),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_1),
.Y(n_356)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_2),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_2),
.B(n_113),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_2),
.B(n_349),
.Y(n_348)
);

NAND2xp33_ASAP7_75t_SL g379 ( 
.A(n_2),
.B(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_3),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_4),
.A2(n_19),
.B(n_452),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_4),
.B(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_5),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_5),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_5),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_5),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_5),
.B(n_297),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_6),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_6),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_8),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_9),
.B(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_9),
.B(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_9),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_9),
.B(n_170),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_9),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_10),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_10),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_10),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_10),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_10),
.B(n_79),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_10),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_10),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_10),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_11),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_11),
.B(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_11),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_11),
.B(n_258),
.Y(n_257)
);

AND2x2_ASAP7_75t_SL g347 ( 
.A(n_11),
.B(n_94),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_11),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_11),
.B(n_391),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_12),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_12),
.Y(n_172)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_12),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_13),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_14),
.B(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_14),
.A2(n_137),
.B1(n_139),
.B2(n_141),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_14),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_14),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_14),
.B(n_308),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_14),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_14),
.B(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_14),
.B(n_396),
.Y(n_395)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_15),
.Y(n_95)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_15),
.Y(n_150)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_16),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_16),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_17),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_44),
.Y(n_43)
);

NAND2x1_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_17),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_17),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_17),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_17),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_17),
.B(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_223),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_222),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp67_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_177),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_24),
.B(n_177),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_99),
.C(n_155),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_26),
.B(n_155),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_68),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_47),
.Y(n_27)
);

MAJx2_ASAP7_75t_L g178 ( 
.A(n_28),
.B(n_47),
.C(n_68),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_37),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_29),
.B(n_43),
.C(n_46),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.C(n_35),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_30),
.B(n_35),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_30),
.B(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_30),
.B(n_251),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_31),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_31),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_32),
.B(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_34),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_34),
.Y(n_283)
);

XNOR2x1_ASAP7_75t_L g157 ( 
.A(n_35),
.B(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_35),
.B(n_126),
.C(n_158),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_35),
.B(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_35),
.B(n_329),
.Y(n_363)
);

INVx8_ASAP7_75t_L g405 ( 
.A(n_36),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B1(n_43),
.B2(n_46),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_42),
.A2(n_43),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_45),
.Y(n_134)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_45),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_45),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_61),
.C(n_66),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_48),
.B(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_54),
.C(n_57),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_50),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_50),
.Y(n_245)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_52),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_54),
.B(n_166),
.Y(n_294)
);

OA21x2_ASAP7_75t_L g335 ( 
.A1(n_54),
.A2(n_204),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_54),
.B(n_204),
.Y(n_336)
);

OAI21xp33_ASAP7_75t_L g367 ( 
.A1(n_54),
.A2(n_204),
.B(n_336),
.Y(n_367)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_56),
.Y(n_393)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_59),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_61),
.A2(n_62),
.B1(n_66),
.B2(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_66),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.C(n_86),
.Y(n_68)
);

XNOR2x1_ASAP7_75t_L g234 ( 
.A(n_69),
.B(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_71),
.A2(n_72),
.B1(n_86),
.B2(n_87),
.Y(n_235)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_77),
.C(n_81),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_73),
.A2(n_78),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_78),
.A2(n_106),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_85),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_85),
.Y(n_331)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_85),
.Y(n_362)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_88),
.Y(n_162)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_93),
.Y(n_163)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_95),
.Y(n_208)
);

INVxp33_ASAP7_75t_SL g164 ( 
.A(n_96),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_100),
.B(n_228),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_130),
.C(n_151),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_102),
.B(n_233),
.Y(n_232)
);

MAJx2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.C(n_117),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_103),
.B(n_108),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.C(n_115),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_112),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_114),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_115),
.B(n_248),
.Y(n_247)
);

XOR2x2_ASAP7_75t_L g437 ( 
.A(n_117),
.B(n_438),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_123),
.C(n_126),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_118),
.B(n_126),
.Y(n_317)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2x2_ASAP7_75t_L g316 ( 
.A(n_123),
.B(n_317),
.Y(n_316)
);

NOR2x1_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_124),
.B(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_124),
.B(n_331),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_124),
.B(n_408),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_126),
.B(n_157),
.Y(n_156)
);

OR2x2_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_130),
.B(n_152),
.Y(n_233)
);

MAJx2_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_136),
.C(n_145),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_132),
.B(n_146),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_134),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_135),
.B(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_136),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_136),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx5_ASAP7_75t_L g357 ( 
.A(n_138),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_139),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_148),
.Y(n_384)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx6_ASAP7_75t_L g334 ( 
.A(n_149),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_150),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_156),
.B(n_161),
.C(n_165),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.C(n_164),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_183),
.C(n_184),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_166),
.A2(n_199),
.B1(n_203),
.B2(n_204),
.Y(n_198)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.Y(n_168)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_172),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_173),
.Y(n_185)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_175),
.Y(n_304)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2x1_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

XNOR2x1_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_209),
.Y(n_179)
);

XOR2x2_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_196),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_186),
.B1(n_194),
.B2(n_195),
.Y(n_181)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

XOR2x2_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_188),
.Y(n_190)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_205),
.B2(n_206),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_199),
.Y(n_203)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_205),
.A2(n_206),
.B1(n_257),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_206),
.B(n_257),
.C(n_260),
.Y(n_256)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_221),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_266),
.B(n_450),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_227),
.B(n_230),
.Y(n_451)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.C(n_236),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_232),
.B(n_234),
.Y(n_440)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_237),
.B(n_440),
.Y(n_439)
);

MAJx2_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_242),
.C(n_246),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_238),
.B(n_242),
.Y(n_435)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OA21x2_ASAP7_75t_SL g306 ( 
.A1(n_241),
.A2(n_307),
.B(n_312),
.Y(n_306)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_246),
.B(n_435),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.C(n_255),
.Y(n_246)
);

XOR2x2_ASAP7_75t_L g289 ( 
.A(n_247),
.B(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_250),
.B(n_256),
.Y(n_290)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_259),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_263),
.Y(n_345)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_265),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_431),
.B(n_446),
.Y(n_266)
);

AO21x2_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_337),
.B(n_430),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_318),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_269),
.B(n_318),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_291),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_289),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_271),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_276),
.C(n_277),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_273),
.B(n_321),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_276),
.Y(n_322)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_284),
.C(n_286),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_279),
.A2(n_280),
.B1(n_284),
.B2(n_285),
.Y(n_371)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_286),
.B(n_371),
.Y(n_370)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

MAJx2_ASAP7_75t_L g442 ( 
.A(n_289),
.B(n_291),
.C(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_305),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_292),
.B(n_306),
.C(n_316),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.C(n_300),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_293),
.A2(n_294),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_295),
.A2(n_296),
.B1(n_300),
.B2(n_301),
.Y(n_325)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_316),
.Y(n_305)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_315),
.Y(n_312)
);

BUFx4f_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_323),
.C(n_326),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_319),
.A2(n_320),
.B1(n_428),
.B2(n_429),
.Y(n_427)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_320),
.B(n_424),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_323),
.B(n_326),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_323),
.B(n_326),
.Y(n_429)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_332),
.C(n_335),
.Y(n_326)
);

XNOR2x1_ASAP7_75t_L g365 ( 
.A(n_327),
.B(n_366),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_332),
.A2(n_335),
.B1(n_367),
.B2(n_368),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_332),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_338),
.A2(n_422),
.B(n_426),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_373),
.B(n_421),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_364),
.Y(n_339)
);

NOR2x1_ASAP7_75t_L g421 ( 
.A(n_340),
.B(n_364),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_353),
.C(n_363),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_342),
.B(n_418),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_346),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_343),
.B(n_347),
.C(n_352),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_344),
.B(n_403),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_351),
.B2(n_352),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_347),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_348),
.Y(n_352)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

AO22x1_ASAP7_75t_L g418 ( 
.A1(n_353),
.A2(n_354),
.B1(n_363),
.B2(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_358),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_355),
.A2(n_358),
.B1(n_359),
.B2(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_355),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_363),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_369),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_365),
.B(n_370),
.C(n_372),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_372),
.Y(n_369)
);

OAI21x1_ASAP7_75t_L g373 ( 
.A1(n_374),
.A2(n_415),
.B(n_420),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_399),
.B(n_414),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_376),
.B(n_388),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_376),
.B(n_388),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_378),
.B1(n_385),
.B2(n_386),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_379),
.B(n_382),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_379),
.B(n_382),
.C(n_385),
.Y(n_416)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_394),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_389),
.A2(n_390),
.B1(n_394),
.B2(n_395),
.Y(n_412)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx3_ASAP7_75t_SL g391 ( 
.A(n_392),
.Y(n_391)
);

INVx8_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

OAI21x1_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_406),
.B(n_413),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx5_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_412),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_407),
.B(n_412),
.Y(n_413)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_417),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_416),
.B(n_417),
.Y(n_420)
);

NOR2x1p5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_425),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_425),
.B(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_441),
.Y(n_431)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_432),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_439),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_433),
.B(n_439),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_436),
.C(n_437),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_434),
.B(n_445),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_436),
.B(n_437),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_444),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g447 ( 
.A(n_442),
.B(n_444),
.Y(n_447)
);

OAI21x1_ASAP7_75t_L g446 ( 
.A1(n_447),
.A2(n_448),
.B(n_449),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);


endmodule