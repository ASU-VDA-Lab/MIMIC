module real_jpeg_7063_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g195 ( 
.A(n_0),
.Y(n_195)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_0),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_0),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g283 ( 
.A(n_0),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_0),
.Y(n_414)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_1),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_1),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g326 ( 
.A(n_1),
.Y(n_326)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_1),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_1),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_2),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_2),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_2),
.A2(n_280),
.B1(n_362),
.B2(n_364),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_2),
.A2(n_280),
.B1(n_285),
.B2(n_388),
.Y(n_387)
);

OAI22xp33_ASAP7_75t_L g452 ( 
.A1(n_2),
.A2(n_46),
.B1(n_280),
.B2(n_453),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_3),
.A2(n_209),
.B1(n_213),
.B2(n_214),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_3),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_3),
.A2(n_201),
.B1(n_213),
.B2(n_235),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_3),
.A2(n_85),
.B1(n_213),
.B2(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_3),
.A2(n_213),
.B1(n_325),
.B2(n_425),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_4),
.A2(n_91),
.B1(n_92),
.B2(n_95),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_4),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_4),
.A2(n_95),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_4),
.A2(n_54),
.B1(n_95),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_4),
.A2(n_95),
.B1(n_378),
.B2(n_379),
.Y(n_377)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_6),
.A2(n_127),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_6),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_6),
.A2(n_169),
.B1(n_201),
.B2(n_204),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_6),
.A2(n_169),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_6),
.A2(n_146),
.B1(n_169),
.B2(n_352),
.Y(n_351)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_7),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_8),
.Y(n_534)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_9),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_9),
.Y(n_108)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_9),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_9),
.Y(n_176)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_11),
.A2(n_160),
.B1(n_162),
.B2(n_165),
.Y(n_159)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_11),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_11),
.B(n_176),
.C(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_11),
.B(n_72),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_11),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_11),
.B(n_125),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_11),
.B(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_12),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_12),
.Y(n_119)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_12),
.Y(n_182)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_14),
.A2(n_82),
.B1(n_85),
.B2(n_88),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_14),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_14),
.A2(n_88),
.B1(n_135),
.B2(n_140),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_14),
.A2(n_88),
.B1(n_178),
.B2(n_374),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_14),
.A2(n_88),
.B1(n_403),
.B2(n_407),
.Y(n_402)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_15),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_15),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_15),
.A2(n_127),
.B1(n_188),
.B2(n_210),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_15),
.A2(n_188),
.B1(n_285),
.B2(n_358),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_15),
.A2(n_49),
.B1(n_56),
.B2(n_188),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_16),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_16),
.A2(n_50),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_16),
.A2(n_50),
.B1(n_209),
.B2(n_364),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_16),
.A2(n_50),
.B1(n_392),
.B2(n_394),
.Y(n_391)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_18),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_18),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_18),
.A2(n_57),
.B1(n_338),
.B2(n_340),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_18),
.A2(n_57),
.B1(n_129),
.B2(n_384),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_18),
.A2(n_57),
.B1(n_388),
.B2(n_438),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_529),
.B(n_532),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_149),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_147),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_144),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_23),
.B(n_144),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_133),
.C(n_141),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_24),
.A2(n_25),
.B1(n_525),
.B2(n_526),
.Y(n_524)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_58),
.C(n_96),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g516 ( 
.A(n_26),
.B(n_517),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_45),
.B1(n_51),
.B2(n_53),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_27),
.A2(n_51),
.B1(n_53),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_27),
.A2(n_51),
.B1(n_134),
.B2(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_27),
.A2(n_350),
.B(n_398),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_27),
.A2(n_51),
.B1(n_398),
.B2(n_424),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_27),
.A2(n_45),
.B1(n_51),
.B2(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_28),
.A2(n_347),
.B(n_349),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_28),
.B(n_351),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_34),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_29)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_30),
.Y(n_328)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx8_ASAP7_75t_L g348 ( 
.A(n_31),
.Y(n_348)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B1(n_41),
.B2(n_43),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_37),
.Y(n_330)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_40),
.Y(n_269)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_51),
.B(n_165),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_51),
.A2(n_424),
.B(n_456),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_52),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_52),
.B(n_452),
.Y(n_451)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_54),
.Y(n_140)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_58),
.A2(n_96),
.B1(n_97),
.B2(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_58),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_81),
.B1(n_89),
.B2(n_90),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_59),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_59),
.A2(n_89),
.B1(n_303),
.B2(n_357),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_59),
.A2(n_89),
.B1(n_387),
.B2(n_391),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_59),
.A2(n_81),
.B1(n_89),
.B2(n_506),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_72),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_63),
.B1(n_67),
.B2(n_70),
.Y(n_60)
);

INVx6_ASAP7_75t_L g292 ( 
.A(n_61),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_63),
.Y(n_272)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_66),
.Y(n_264)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_66),
.Y(n_324)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_66),
.Y(n_440)
);

AO22x2_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_73),
.B1(n_77),
.B2(n_79),
.Y(n_72)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_69),
.Y(n_290)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_71),
.Y(n_396)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_72),
.A2(n_142),
.B(n_143),
.Y(n_141)
);

AOI22x1_ASAP7_75t_L g427 ( 
.A1(n_72),
.A2(n_142),
.B1(n_306),
.B2(n_428),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_72),
.A2(n_142),
.B1(n_436),
.B2(n_437),
.Y(n_435)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_76),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g406 ( 
.A(n_76),
.Y(n_406)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_82),
.B(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_84),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_84),
.Y(n_393)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_86),
.Y(n_273)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_89),
.B(n_271),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_89),
.A2(n_303),
.B(n_305),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_91),
.Y(n_285)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_96),
.A2(n_97),
.B1(n_504),
.B2(n_505),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_96),
.B(n_501),
.C(n_504),
.Y(n_512)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_124),
.B(n_126),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_98),
.A2(n_159),
.B(n_166),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_98),
.A2(n_124),
.B1(n_208),
.B2(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_98),
.A2(n_166),
.B(n_260),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_98),
.A2(n_124),
.B1(n_361),
.B2(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_99),
.B(n_167),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_99),
.A2(n_125),
.B1(n_382),
.B2(n_383),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_99),
.A2(n_125),
.B1(n_383),
.B2(n_402),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_99),
.A2(n_125),
.B1(n_402),
.B2(n_443),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_111),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B1(n_106),
.B2(n_109),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g364 ( 
.A(n_101),
.Y(n_364)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_102),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_110),
.Y(n_288)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_111),
.A2(n_208),
.B(n_217),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_114),
.B1(n_118),
.B2(n_120),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_117),
.Y(n_197)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_117),
.Y(n_282)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_117),
.Y(n_311)
);

BUFx8_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_119),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_119),
.Y(n_237)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_124),
.A2(n_217),
.B(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_125),
.B(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_126),
.Y(n_443)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp33_ASAP7_75t_SL g291 ( 
.A(n_130),
.B(n_292),
.Y(n_291)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_132),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_132),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_132),
.Y(n_363)
);

INVx6_ASAP7_75t_L g410 ( 
.A(n_132),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_133),
.B(n_141),
.Y(n_526)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_136),
.B(n_165),
.Y(n_331)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_139),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_142),
.A2(n_263),
.B(n_270),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_142),
.B(n_306),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_142),
.A2(n_270),
.B(n_469),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_523),
.B(n_528),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_495),
.B(n_520),
.Y(n_150)
);

OAI311xp33_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_367),
.A3(n_471),
.B1(n_489),
.C1(n_490),
.Y(n_151)
);

AOI21x1_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_317),
.B(n_366),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_294),
.B(n_316),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_254),
.B(n_293),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_220),
.B(n_253),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_183),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_157),
.B(n_183),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_170),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_158),
.A2(n_170),
.B1(n_171),
.B2(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_158),
.Y(n_251)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_165),
.A2(n_192),
.B(n_198),
.Y(n_231)
);

OAI21xp33_ASAP7_75t_SL g263 ( 
.A1(n_165),
.A2(n_264),
.B(n_265),
.Y(n_263)
);

OAI21xp33_ASAP7_75t_SL g347 ( 
.A1(n_165),
.A2(n_331),
.B(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_180),
.Y(n_339)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_205),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_184),
.B(n_206),
.C(n_219),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_192),
.B(n_198),
.Y(n_184)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_185),
.Y(n_246)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_189),
.Y(n_312)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_191),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_192),
.A2(n_334),
.B1(n_335),
.B2(n_336),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_192),
.A2(n_248),
.B1(n_373),
.B2(n_377),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_192),
.A2(n_377),
.B(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_200),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_193),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_193),
.A2(n_277),
.B1(n_310),
.B2(n_313),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_193),
.A2(n_313),
.B1(n_337),
.B2(n_421),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_194),
.Y(n_239)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_195),
.Y(n_249)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_195),
.Y(n_314)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_203),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_218),
.B2(n_219),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx11_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_243),
.B(n_252),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_232),
.B(n_242),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_231),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_228),
.Y(n_279)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_228),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_241),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_241),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_238),
.B(n_240),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_240),
.A2(n_276),
.B(n_283),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_250),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_250),
.Y(n_252)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_256),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_274),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_259),
.B(n_261),
.C(n_274),
.Y(n_295)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI32xp33_ASAP7_75t_L g284 ( 
.A1(n_266),
.A2(n_285),
.A3(n_286),
.B1(n_289),
.B2(n_291),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_268),
.Y(n_267)
);

INVx6_ASAP7_75t_SL g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_271),
.Y(n_306)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_273),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_284),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_284),
.Y(n_300)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx5_ASAP7_75t_SL g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_295),
.B(n_296),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_301),
.B2(n_315),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_300),
.C(n_315),
.Y(n_318)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_307),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_302),
.B(n_308),
.C(n_309),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_310),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_313),
.Y(n_335)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_318),
.B(n_319),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_344),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_341),
.B1(n_342),
.B2(n_343),
.Y(n_320)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_321),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_332),
.B2(n_333),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_323),
.B(n_332),
.Y(n_467)
);

OAI32xp33_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_325),
.A3(n_327),
.B1(n_329),
.B2(n_331),
.Y(n_323)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_338),
.Y(n_378)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_341),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_341),
.B(n_342),
.C(n_344),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_346),
.B1(n_355),
.B2(n_365),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_345),
.B(n_356),
.C(n_360),
.Y(n_480)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_355),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_360),
.Y(n_355)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_357),
.Y(n_469)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx5_ASAP7_75t_L g390 ( 
.A(n_359),
.Y(n_390)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

NAND2xp33_ASAP7_75t_SL g367 ( 
.A(n_368),
.B(n_457),
.Y(n_367)
);

A2O1A1Ixp33_ASAP7_75t_SL g490 ( 
.A1(n_368),
.A2(n_457),
.B(n_491),
.C(n_494),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_429),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_369),
.B(n_429),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_399),
.C(n_416),
.Y(n_369)
);

FAx1_ASAP7_75t_L g470 ( 
.A(n_370),
.B(n_399),
.CI(n_416),
.CON(n_470),
.SN(n_470)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_385),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_371),
.B(n_386),
.C(n_397),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_381),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_372),
.B(n_381),
.Y(n_463)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_373),
.Y(n_421)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_382),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_397),
.Y(n_385)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_387),
.Y(n_428)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx4_ASAP7_75t_SL g389 ( 
.A(n_390),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_391),
.Y(n_436)
);

INVx6_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_400),
.A2(n_401),
.B1(n_411),
.B2(n_415),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_401),
.B(n_411),
.Y(n_447)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx5_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx8_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_411),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_411),
.A2(n_415),
.B1(n_449),
.B2(n_450),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_411),
.A2(n_447),
.B(n_450),
.Y(n_498)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_422),
.C(n_427),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_417),
.B(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_418),
.B(n_420),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_418),
.B(n_420),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_422),
.A2(n_423),
.B1(n_427),
.B2(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx6_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_427),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_430),
.B(n_433),
.C(n_445),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_433),
.B1(n_445),
.B2(n_446),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_434),
.A2(n_441),
.B(n_444),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_435),
.B(n_442),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_437),
.Y(n_506)
);

INVx5_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

FAx1_ASAP7_75t_SL g497 ( 
.A(n_444),
.B(n_498),
.CI(n_499),
.CON(n_497),
.SN(n_497)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_444),
.B(n_498),
.C(n_499),
.Y(n_519)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_456),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_452),
.Y(n_502)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_470),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_458),
.B(n_470),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_463),
.C(n_464),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_459),
.A2(n_460),
.B1(n_463),
.B2(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_463),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_482),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_467),
.C(n_468),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_465),
.A2(n_466),
.B1(n_468),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_467),
.B(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_468),
.Y(n_477)
);

BUFx24_ASAP7_75t_SL g537 ( 
.A(n_470),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_484),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_473),
.A2(n_492),
.B(n_493),
.Y(n_491)
);

NOR2x1_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_481),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_474),
.B(n_481),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_478),
.C(n_480),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_487),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_478),
.A2(n_479),
.B1(n_480),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_480),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_486),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_485),
.B(n_486),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_509),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_497),
.B(n_508),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_497),
.B(n_508),
.Y(n_521)
);

BUFx24_ASAP7_75t_SL g536 ( 
.A(n_497),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_501),
.B1(n_503),
.B2(n_507),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_500),
.A2(n_501),
.B1(n_515),
.B2(n_516),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_500),
.B(n_511),
.C(n_515),
.Y(n_527)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_503),
.Y(n_507)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_509),
.A2(n_521),
.B(n_522),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_510),
.B(n_519),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_510),
.B(n_519),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_511),
.A2(n_512),
.B1(n_513),
.B2(n_514),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_527),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_524),
.B(n_527),
.Y(n_528)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx13_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx6_ASAP7_75t_L g533 ( 
.A(n_531),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_534),
.Y(n_532)
);


endmodule