module real_aes_15407_n_234 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_234);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_234;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_239;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_238;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_246;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_247;
wire n_264;
wire n_237;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_245;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_248;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_1404;
wire n_733;
wire n_402;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_265;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1403;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_249;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_243;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_241;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_236;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_244;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1352;
wire n_1323;
wire n_1369;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_240;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g440 ( .A(n_0), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g1226 ( .A1(n_0), .A2(n_191), .B1(n_1170), .B2(n_1174), .Y(n_1226) );
INVx1_ASAP7_75t_L g369 ( .A(n_1), .Y(n_369) );
AOI221x1_ASAP7_75t_SL g405 ( .A1(n_1), .A2(n_3), .B1(n_406), .B2(n_409), .C(n_411), .Y(n_405) );
INVx1_ASAP7_75t_L g767 ( .A(n_2), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_3), .A2(n_18), .B1(n_375), .B2(n_377), .Y(n_387) );
OAI211xp5_ASAP7_75t_L g833 ( .A1(n_4), .A2(n_738), .B(n_830), .C(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g851 ( .A(n_4), .Y(n_851) );
AOI221x1_ASAP7_75t_SL g454 ( .A1(n_5), .A2(n_226), .B1(n_455), .B2(n_459), .C(n_461), .Y(n_454) );
AOI21xp33_ASAP7_75t_L g545 ( .A1(n_5), .A2(n_424), .B(n_546), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g1194 ( .A1(n_6), .A2(n_50), .B1(n_1170), .B2(n_1174), .Y(n_1194) );
XNOR2xp5_ASAP7_75t_L g1372 ( .A(n_6), .B(n_1373), .Y(n_1372) );
AOI22xp33_ASAP7_75t_L g1417 ( .A1(n_6), .A2(n_1418), .B1(n_1421), .B2(n_1424), .Y(n_1417) );
INVx1_ASAP7_75t_L g1142 ( .A(n_7), .Y(n_1142) );
INVx1_ASAP7_75t_L g895 ( .A(n_8), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_8), .A2(n_98), .B1(n_549), .B2(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g1055 ( .A(n_9), .Y(n_1055) );
OAI22xp33_ASAP7_75t_L g1099 ( .A1(n_9), .A2(n_112), .B1(n_1100), .B2(n_1101), .Y(n_1099) );
AOI21xp33_ASAP7_75t_L g383 ( .A1(n_10), .A2(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_L g428 ( .A(n_10), .Y(n_428) );
INVx1_ASAP7_75t_L g247 ( .A(n_11), .Y(n_247) );
AND2x2_ASAP7_75t_L g278 ( .A(n_11), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g366 ( .A(n_11), .B(n_206), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_11), .B(n_257), .Y(n_475) );
OAI221xp5_ASAP7_75t_L g1060 ( .A1(n_12), .A2(n_227), .B1(n_1061), .B2(n_1062), .C(n_1066), .Y(n_1060) );
INVx1_ASAP7_75t_L g1096 ( .A(n_12), .Y(n_1096) );
OAI211xp5_ASAP7_75t_L g1113 ( .A1(n_13), .A2(n_368), .B(n_1114), .C(n_1118), .Y(n_1113) );
INVx1_ASAP7_75t_L g1123 ( .A(n_13), .Y(n_1123) );
OAI22xp33_ASAP7_75t_L g609 ( .A1(n_14), .A2(n_190), .B1(n_610), .B2(n_613), .Y(n_609) );
OAI22xp33_ASAP7_75t_L g648 ( .A1(n_14), .A2(n_190), .B1(n_649), .B2(n_652), .Y(n_648) );
INVx1_ASAP7_75t_L g1381 ( .A(n_15), .Y(n_1381) );
INVx2_ASAP7_75t_L g1173 ( .A(n_16), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_16), .B(n_92), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_16), .B(n_1179), .Y(n_1181) );
INVx1_ASAP7_75t_L g1405 ( .A(n_17), .Y(n_1405) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_18), .A2(n_161), .B1(n_409), .B2(n_422), .C(n_425), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_19), .A2(n_144), .B1(n_649), .B2(n_1108), .Y(n_1107) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_19), .A2(n_144), .B1(n_613), .B2(n_1125), .Y(n_1124) );
AOI22xp5_ASAP7_75t_L g1203 ( .A1(n_20), .A2(n_33), .B1(n_1177), .B2(n_1180), .Y(n_1203) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_21), .A2(n_129), .B1(n_495), .B2(n_498), .Y(n_494) );
OAI221xp5_ASAP7_75t_L g506 ( .A1(n_21), .A2(n_209), .B1(n_507), .B2(n_509), .C(n_511), .Y(n_506) );
OAI22xp33_ASAP7_75t_L g959 ( .A1(n_22), .A2(n_223), .B1(n_744), .B2(n_960), .Y(n_959) );
OAI22xp33_ASAP7_75t_L g972 ( .A1(n_22), .A2(n_223), .B1(n_853), .B2(n_973), .Y(n_972) );
INVx1_ASAP7_75t_L g680 ( .A(n_23), .Y(n_680) );
OAI22xp33_ASAP7_75t_L g743 ( .A1(n_24), .A2(n_51), .B1(n_744), .B2(n_745), .Y(n_743) );
OAI22xp33_ASAP7_75t_L g753 ( .A1(n_24), .A2(n_51), .B1(n_754), .B2(n_755), .Y(n_753) );
OAI22xp33_ASAP7_75t_L g1112 ( .A1(n_25), .A2(n_38), .B1(n_249), .B2(n_645), .Y(n_1112) );
OAI22xp33_ASAP7_75t_L g1120 ( .A1(n_25), .A2(n_38), .B1(n_632), .B2(n_716), .Y(n_1120) );
AOI22xp5_ASAP7_75t_L g1225 ( .A1(n_26), .A2(n_110), .B1(n_1177), .B2(n_1180), .Y(n_1225) );
INVx1_ASAP7_75t_L g928 ( .A(n_27), .Y(n_928) );
OAI211xp5_ASAP7_75t_L g1403 ( .A1(n_28), .A2(n_619), .B(n_823), .C(n_1404), .Y(n_1403) );
INVx1_ASAP7_75t_L g1412 ( .A(n_28), .Y(n_1412) );
INVx1_ASAP7_75t_L g560 ( .A(n_29), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g951 ( .A1(n_30), .A2(n_116), .B1(n_952), .B2(n_954), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_30), .A2(n_116), .B1(n_645), .B2(n_965), .Y(n_964) );
OAI22xp33_ASAP7_75t_L g832 ( .A1(n_31), .A2(n_166), .B1(n_634), .B2(n_735), .Y(n_832) );
OAI22xp33_ASAP7_75t_L g842 ( .A1(n_31), .A2(n_166), .B1(n_249), .B2(n_758), .Y(n_842) );
INVx1_ASAP7_75t_L g861 ( .A(n_32), .Y(n_861) );
INVx1_ASAP7_75t_L g1034 ( .A(n_34), .Y(n_1034) );
INVx1_ASAP7_75t_L g1141 ( .A(n_35), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1263 ( .A1(n_36), .A2(n_88), .B1(n_1170), .B2(n_1264), .Y(n_1263) );
INVx1_ASAP7_75t_L g813 ( .A(n_37), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g1200 ( .A1(n_39), .A2(n_84), .B1(n_1170), .B2(n_1191), .Y(n_1200) );
CKINVDCx5p33_ASAP7_75t_R g1003 ( .A(n_40), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_41), .A2(n_67), .B1(n_526), .B2(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g1025 ( .A(n_41), .Y(n_1025) );
AOI221xp5_ASAP7_75t_L g1048 ( .A1(n_42), .A2(n_124), .B1(n_1049), .B2(n_1050), .C(n_1051), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_42), .A2(n_71), .B1(n_995), .B2(n_1088), .Y(n_1094) );
INVx1_ASAP7_75t_L g741 ( .A(n_43), .Y(n_741) );
OAI22xp5_ASAP7_75t_SL g339 ( .A1(n_44), .A2(n_162), .B1(n_340), .B2(n_344), .Y(n_339) );
INVx1_ASAP7_75t_L g351 ( .A(n_44), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_45), .A2(n_152), .B1(n_391), .B2(n_485), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_45), .A2(n_91), .B1(n_406), .B2(n_993), .Y(n_1093) );
INVx1_ASAP7_75t_L g1138 ( .A(n_46), .Y(n_1138) );
INVx1_ASAP7_75t_L g289 ( .A(n_47), .Y(n_289) );
INVx1_ASAP7_75t_L g337 ( .A(n_47), .Y(n_337) );
INVx1_ASAP7_75t_L g805 ( .A(n_48), .Y(n_805) );
OAI22xp5_ASAP7_75t_L g858 ( .A1(n_49), .A2(n_859), .B1(n_919), .B2(n_920), .Y(n_858) );
INVxp67_ASAP7_75t_L g920 ( .A(n_49), .Y(n_920) );
AOI22xp5_ASAP7_75t_L g1190 ( .A1(n_49), .A2(n_119), .B1(n_1170), .B2(n_1191), .Y(n_1190) );
INVx1_ASAP7_75t_L g1406 ( .A(n_52), .Y(n_1406) );
OAI211xp5_ASAP7_75t_L g1410 ( .A1(n_52), .A2(n_658), .B(n_749), .C(n_1411), .Y(n_1410) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_53), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g873 ( .A(n_54), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_55), .A2(n_204), .B1(n_1177), .B2(n_1180), .Y(n_1265) );
OAI22xp33_ASAP7_75t_L g714 ( .A1(n_56), .A2(n_185), .B1(n_715), .B2(n_716), .Y(n_714) );
OAI22xp33_ASAP7_75t_L g719 ( .A1(n_56), .A2(n_185), .B1(n_249), .B2(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g240 ( .A(n_57), .Y(n_240) );
INVx2_ASAP7_75t_L g295 ( .A(n_58), .Y(n_295) );
INVx1_ASAP7_75t_L g568 ( .A(n_59), .Y(n_568) );
XOR2x2_ASAP7_75t_L g729 ( .A(n_60), .B(n_730), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_61), .A2(n_230), .B1(n_375), .B2(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g906 ( .A(n_61), .Y(n_906) );
INVx1_ASAP7_75t_L g685 ( .A(n_62), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g1080 ( .A1(n_63), .A2(n_200), .B1(n_311), .B2(n_1081), .Y(n_1080) );
INVx1_ASAP7_75t_L g1148 ( .A(n_64), .Y(n_1148) );
INVx1_ASAP7_75t_L g1079 ( .A(n_65), .Y(n_1079) );
XOR2xp5_ASAP7_75t_L g1422 ( .A(n_66), .B(n_1423), .Y(n_1422) );
AOI221xp5_ASAP7_75t_L g1005 ( .A1(n_67), .A2(n_114), .B1(n_898), .B2(n_1006), .C(n_1008), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_68), .A2(n_98), .B1(n_377), .B2(n_883), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_68), .A2(n_179), .B1(n_526), .B2(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g1117 ( .A(n_69), .Y(n_1117) );
OAI211xp5_ASAP7_75t_L g1121 ( .A1(n_69), .A2(n_619), .B(n_830), .C(n_1122), .Y(n_1121) );
INVx1_ASAP7_75t_L g780 ( .A(n_70), .Y(n_780) );
INVxp67_ASAP7_75t_SL g1069 ( .A(n_71), .Y(n_1069) );
XOR2x2_ASAP7_75t_L g1103 ( .A(n_72), .B(n_1104), .Y(n_1103) );
INVx1_ASAP7_75t_L g837 ( .A(n_73), .Y(n_837) );
OAI211xp5_ASAP7_75t_L g843 ( .A1(n_73), .A2(n_355), .B(n_844), .C(n_848), .Y(n_843) );
AOI22xp5_ASAP7_75t_L g1176 ( .A1(n_74), .A2(n_115), .B1(n_1177), .B2(n_1180), .Y(n_1176) );
AOI22xp33_ASAP7_75t_L g1211 ( .A1(n_75), .A2(n_96), .B1(n_1170), .B2(n_1174), .Y(n_1211) );
INVx1_ASAP7_75t_L g580 ( .A(n_76), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g1002 ( .A(n_77), .Y(n_1002) );
OAI221xp5_ASAP7_75t_SL g867 ( .A1(n_78), .A2(n_83), .B1(n_868), .B2(n_870), .C(n_872), .Y(n_867) );
INVx1_ASAP7_75t_L g890 ( .A(n_78), .Y(n_890) );
INVx1_ASAP7_75t_L g381 ( .A(n_79), .Y(n_381) );
INVx1_ASAP7_75t_L g818 ( .A(n_80), .Y(n_818) );
INVx1_ASAP7_75t_L g626 ( .A(n_81), .Y(n_626) );
INVx1_ASAP7_75t_L g817 ( .A(n_82), .Y(n_817) );
INVx1_ASAP7_75t_L g900 ( .A(n_83), .Y(n_900) );
OA222x2_ASAP7_75t_L g442 ( .A1(n_85), .A2(n_192), .B1(n_209), .B2(n_443), .C1(n_447), .C2(n_451), .Y(n_442) );
INVx1_ASAP7_75t_L g524 ( .A(n_85), .Y(n_524) );
INVx1_ASAP7_75t_L g935 ( .A(n_86), .Y(n_935) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_87), .Y(n_242) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_87), .B(n_240), .Y(n_1171) );
INVx1_ASAP7_75t_L g931 ( .A(n_89), .Y(n_931) );
CKINVDCx5p33_ASAP7_75t_R g998 ( .A(n_90), .Y(n_998) );
AOI221xp5_ASAP7_75t_L g1070 ( .A1(n_91), .A2(n_141), .B1(n_457), .B2(n_1071), .C(n_1073), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_92), .B(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1179 ( .A(n_92), .Y(n_1179) );
AOI22xp5_ASAP7_75t_L g1189 ( .A1(n_93), .A2(n_151), .B1(n_1177), .B2(n_1180), .Y(n_1189) );
OAI211xp5_ASAP7_75t_SL g615 ( .A1(n_94), .A2(n_616), .B(n_619), .C(n_621), .Y(n_615) );
INVx1_ASAP7_75t_L g670 ( .A(n_94), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_95), .A2(n_100), .B1(n_409), .B2(n_828), .Y(n_989) );
INVx1_ASAP7_75t_L g1027 ( .A(n_95), .Y(n_1027) );
INVx1_ASAP7_75t_L g984 ( .A(n_97), .Y(n_984) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_97), .A2(n_212), .B1(n_464), .B2(n_468), .Y(n_1018) );
INVx1_ASAP7_75t_L g776 ( .A(n_99), .Y(n_776) );
INVx1_ASAP7_75t_L g1010 ( .A(n_100), .Y(n_1010) );
INVx1_ASAP7_75t_L g932 ( .A(n_101), .Y(n_932) );
INVx1_ASAP7_75t_L g865 ( .A(n_102), .Y(n_865) );
INVx1_ASAP7_75t_L g929 ( .A(n_103), .Y(n_929) );
OAI211xp5_ASAP7_75t_L g955 ( .A1(n_104), .A2(n_429), .B(n_738), .C(n_956), .Y(n_955) );
INVx1_ASAP7_75t_L g971 ( .A(n_104), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_105), .B(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g318 ( .A(n_105), .Y(n_318) );
INVx1_ASAP7_75t_L g420 ( .A(n_105), .Y(n_420) );
OAI22xp33_ASAP7_75t_L g838 ( .A1(n_106), .A2(n_214), .B1(n_744), .B2(n_839), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_106), .A2(n_214), .B1(n_853), .B2(n_854), .Y(n_852) );
INVx1_ASAP7_75t_L g682 ( .A(n_107), .Y(n_682) );
OAI22xp33_ASAP7_75t_L g732 ( .A1(n_108), .A2(n_228), .B1(n_733), .B2(n_735), .Y(n_732) );
OAI22xp33_ASAP7_75t_L g757 ( .A1(n_108), .A2(n_228), .B1(n_249), .B2(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g1382 ( .A(n_109), .Y(n_1382) );
INVx1_ASAP7_75t_L g958 ( .A(n_111), .Y(n_958) );
OAI211xp5_ASAP7_75t_L g968 ( .A1(n_111), .A2(n_844), .B(n_969), .C(n_970), .Y(n_968) );
INVx1_ASAP7_75t_L g1057 ( .A(n_112), .Y(n_1057) );
OAI211xp5_ASAP7_75t_L g704 ( .A1(n_113), .A2(n_619), .B(n_705), .C(n_708), .Y(n_704) );
INVx1_ASAP7_75t_L g724 ( .A(n_113), .Y(n_724) );
AOI22xp33_ASAP7_75t_SL g994 ( .A1(n_114), .A2(n_145), .B1(n_988), .B2(n_995), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_117), .A2(n_225), .B1(n_391), .B2(n_485), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_117), .A2(n_211), .B1(n_410), .B2(n_549), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g1212 ( .A1(n_118), .A2(n_216), .B1(n_1177), .B2(n_1180), .Y(n_1212) );
AOI22xp5_ASAP7_75t_L g1169 ( .A1(n_120), .A2(n_121), .B1(n_1170), .B2(n_1174), .Y(n_1169) );
INVx1_ASAP7_75t_L g1377 ( .A(n_122), .Y(n_1377) );
INVx1_ASAP7_75t_L g574 ( .A(n_123), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_124), .A2(n_159), .B1(n_1086), .B2(n_1089), .Y(n_1085) );
INVx1_ASAP7_75t_L g683 ( .A(n_125), .Y(n_683) );
INVx1_ASAP7_75t_L g266 ( .A(n_126), .Y(n_266) );
INVx1_ASAP7_75t_L g692 ( .A(n_127), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g1193 ( .A1(n_128), .A2(n_136), .B1(n_1177), .B2(n_1180), .Y(n_1193) );
INVx1_ASAP7_75t_L g525 ( .A(n_129), .Y(n_525) );
INVx1_ASAP7_75t_L g1391 ( .A(n_130), .Y(n_1391) );
OAI22xp33_ASAP7_75t_L g1407 ( .A1(n_131), .A2(n_146), .B1(n_610), .B2(n_839), .Y(n_1407) );
OAI22xp5_ASAP7_75t_L g1413 ( .A1(n_131), .A2(n_146), .B1(n_755), .B2(n_853), .Y(n_1413) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_132), .Y(n_483) );
INVx1_ASAP7_75t_L g808 ( .A(n_133), .Y(n_808) );
INVx1_ASAP7_75t_L g810 ( .A(n_134), .Y(n_810) );
INVx1_ASAP7_75t_L g1147 ( .A(n_135), .Y(n_1147) );
INVx1_ASAP7_75t_L g934 ( .A(n_137), .Y(n_934) );
BUFx3_ASAP7_75t_L g287 ( .A(n_138), .Y(n_287) );
INVx1_ASAP7_75t_L g709 ( .A(n_139), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g1201 ( .A1(n_140), .A2(n_142), .B1(n_1177), .B2(n_1180), .Y(n_1201) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_141), .A2(n_152), .B1(n_828), .B2(n_1091), .Y(n_1090) );
AOI22xp5_ASAP7_75t_L g1204 ( .A1(n_143), .A2(n_207), .B1(n_1170), .B2(n_1174), .Y(n_1204) );
AOI211xp5_ASAP7_75t_SL g1022 ( .A1(n_145), .A2(n_1023), .B(n_1024), .C(n_1026), .Y(n_1022) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_147), .Y(n_254) );
INVx1_ASAP7_75t_L g864 ( .A(n_148), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_149), .A2(n_181), .B1(n_991), .B2(n_993), .Y(n_990) );
INVx1_ASAP7_75t_L g1009 ( .A(n_149), .Y(n_1009) );
INVx1_ASAP7_75t_L g679 ( .A(n_150), .Y(n_679) );
INVx1_ASAP7_75t_L g939 ( .A(n_153), .Y(n_939) );
INVx1_ASAP7_75t_L g710 ( .A(n_154), .Y(n_710) );
OAI211xp5_ASAP7_75t_L g722 ( .A1(n_154), .A2(n_658), .B(n_661), .C(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g1392 ( .A(n_155), .Y(n_1392) );
INVx1_ASAP7_75t_L g1386 ( .A(n_156), .Y(n_1386) );
XNOR2xp5_ASAP7_75t_L g553 ( .A(n_157), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g742 ( .A(n_158), .Y(n_742) );
OAI211xp5_ASAP7_75t_L g748 ( .A1(n_158), .A2(n_660), .B(n_749), .C(n_750), .Y(n_748) );
INVxp67_ASAP7_75t_SL g1067 ( .A(n_159), .Y(n_1067) );
INVx1_ASAP7_75t_L g1131 ( .A(n_160), .Y(n_1131) );
AOI21xp33_ASAP7_75t_L g370 ( .A1(n_161), .A2(n_371), .B(n_372), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_162), .Y(n_362) );
OAI22xp33_ASAP7_75t_L g631 ( .A1(n_163), .A2(n_221), .B1(n_632), .B2(n_635), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_163), .A2(n_221), .B1(n_644), .B2(n_645), .Y(n_643) );
XNOR2xp5_ASAP7_75t_L g674 ( .A(n_164), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g689 ( .A(n_165), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g980 ( .A(n_167), .Y(n_980) );
XOR2x2_ASAP7_75t_L g1040 ( .A(n_168), .B(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_L g1115 ( .A(n_169), .Y(n_1115) );
INVx1_ASAP7_75t_L g802 ( .A(n_170), .Y(n_802) );
OAI222xp33_ASAP7_75t_L g268 ( .A1(n_171), .A2(n_208), .B1(n_218), .B2(n_269), .C1(n_296), .C2(n_311), .Y(n_268) );
INVx1_ASAP7_75t_L g564 ( .A(n_172), .Y(n_564) );
INVx1_ASAP7_75t_L g765 ( .A(n_173), .Y(n_765) );
INVx1_ASAP7_75t_L g773 ( .A(n_174), .Y(n_773) );
INVx1_ASAP7_75t_L g576 ( .A(n_175), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_176), .A2(n_231), .B1(n_375), .B2(n_377), .Y(n_374) );
INVxp67_ASAP7_75t_SL g426 ( .A(n_176), .Y(n_426) );
XOR2x2_ASAP7_75t_L g795 ( .A(n_177), .B(n_796), .Y(n_795) );
OAI211xp5_ASAP7_75t_L g736 ( .A1(n_178), .A2(n_737), .B(n_738), .C(n_739), .Y(n_736) );
INVx1_ASAP7_75t_L g752 ( .A(n_178), .Y(n_752) );
AOI21xp33_ASAP7_75t_L g896 ( .A1(n_179), .A2(n_384), .B(n_385), .Y(n_896) );
INVx1_ASAP7_75t_L g836 ( .A(n_180), .Y(n_836) );
INVx1_ASAP7_75t_L g1029 ( .A(n_181), .Y(n_1029) );
INVx1_ASAP7_75t_L g687 ( .A(n_182), .Y(n_687) );
INVx1_ASAP7_75t_L g630 ( .A(n_183), .Y(n_630) );
OAI211xp5_ASAP7_75t_L g657 ( .A1(n_183), .A2(n_658), .B(n_661), .C(n_664), .Y(n_657) );
INVx1_ASAP7_75t_L g1134 ( .A(n_184), .Y(n_1134) );
INVx1_ASAP7_75t_L g1387 ( .A(n_186), .Y(n_1387) );
INVx1_ASAP7_75t_L g770 ( .A(n_187), .Y(n_770) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_188), .Y(n_253) );
OAI22xp33_ASAP7_75t_L g1402 ( .A1(n_189), .A2(n_201), .B1(n_735), .B2(n_952), .Y(n_1402) );
OAI22xp33_ASAP7_75t_L g1409 ( .A1(n_189), .A2(n_201), .B1(n_249), .B2(n_720), .Y(n_1409) );
INVx1_ASAP7_75t_L g512 ( .A(n_192), .Y(n_512) );
INVx1_ASAP7_75t_L g579 ( .A(n_193), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_194), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g879 ( .A1(n_195), .A2(n_203), .B1(n_372), .B2(n_460), .C(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g905 ( .A(n_195), .Y(n_905) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_196), .Y(n_330) );
INVx1_ASAP7_75t_L g1379 ( .A(n_197), .Y(n_1379) );
INVx1_ASAP7_75t_L g777 ( .A(n_198), .Y(n_777) );
INVx1_ASAP7_75t_L g812 ( .A(n_199), .Y(n_812) );
OAI211xp5_ASAP7_75t_L g1043 ( .A1(n_200), .A2(n_1044), .B(n_1047), .C(n_1054), .Y(n_1043) );
OAI22xp33_ASAP7_75t_L g711 ( .A1(n_202), .A2(n_233), .B1(n_613), .B2(n_712), .Y(n_711) );
OAI22xp33_ASAP7_75t_L g721 ( .A1(n_202), .A2(n_233), .B1(n_649), .B2(n_652), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_203), .A2(n_230), .B1(n_914), .B2(n_915), .Y(n_913) );
CKINVDCx5p33_ASAP7_75t_R g875 ( .A(n_205), .Y(n_875) );
BUFx3_ASAP7_75t_L g257 ( .A(n_206), .Y(n_257) );
INVx1_ASAP7_75t_L g279 ( .A(n_206), .Y(n_279) );
XOR2x2_ASAP7_75t_L g923 ( .A(n_207), .B(n_924), .Y(n_923) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_210), .Y(n_478) );
INVx1_ASAP7_75t_L g462 ( .A(n_211), .Y(n_462) );
INVx1_ASAP7_75t_L g1032 ( .A(n_212), .Y(n_1032) );
INVx1_ASAP7_75t_L g1139 ( .A(n_213), .Y(n_1139) );
INVx1_ASAP7_75t_L g957 ( .A(n_215), .Y(n_957) );
INVx1_ASAP7_75t_L g276 ( .A(n_217), .Y(n_276) );
INVx1_ASAP7_75t_L g329 ( .A(n_217), .Y(n_329) );
INVx2_ASAP7_75t_L g403 ( .A(n_217), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_218), .A2(n_224), .B1(n_389), .B2(n_393), .Y(n_388) );
INVx1_ASAP7_75t_L g781 ( .A(n_219), .Y(n_781) );
INVx1_ASAP7_75t_L g937 ( .A(n_220), .Y(n_937) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_222), .Y(n_504) );
INVx1_ASAP7_75t_L g338 ( .A(n_224), .Y(n_338) );
INVx1_ASAP7_75t_L g543 ( .A(n_225), .Y(n_543) );
INVx1_ASAP7_75t_L g540 ( .A(n_226), .Y(n_540) );
INVx1_ASAP7_75t_L g1098 ( .A(n_227), .Y(n_1098) );
CKINVDCx5p33_ASAP7_75t_R g985 ( .A(n_229), .Y(n_985) );
INVx1_ASAP7_75t_L g412 ( .A(n_231), .Y(n_412) );
INVx1_ASAP7_75t_L g570 ( .A(n_232), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_258), .B(n_1163), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_243), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g1416 ( .A(n_237), .B(n_246), .Y(n_1416) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_239), .B(n_241), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g1420 ( .A(n_239), .B(n_242), .Y(n_1420) );
INVx1_ASAP7_75t_L g1425 ( .A(n_239), .Y(n_1425) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g1427 ( .A(n_242), .B(n_1425), .Y(n_1427) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_248), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x4_ASAP7_75t_L g672 ( .A(n_246), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x4_ASAP7_75t_L g373 ( .A(n_247), .B(n_256), .Y(n_373) );
AND2x4_ASAP7_75t_L g386 ( .A(n_247), .B(n_257), .Y(n_386) );
INVxp67_ASAP7_75t_SL g644 ( .A(n_248), .Y(n_644) );
AND2x4_ASAP7_75t_SL g1415 ( .A(n_248), .B(n_1416), .Y(n_1415) );
INVx3_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OR2x6_ASAP7_75t_L g249 ( .A(n_250), .B(n_255), .Y(n_249) );
INVx1_ASAP7_75t_L g605 ( .A(n_250), .Y(n_605) );
OR2x6_ASAP7_75t_L g651 ( .A(n_250), .B(n_647), .Y(n_651) );
BUFx4f_ASAP7_75t_L g779 ( .A(n_250), .Y(n_779) );
INVxp67_ASAP7_75t_L g804 ( .A(n_250), .Y(n_804) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx3_ASAP7_75t_L g464 ( .A(n_251), .Y(n_464) );
BUFx4f_ASAP7_75t_L g587 ( .A(n_251), .Y(n_587) );
INVx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
INVx2_ASAP7_75t_L g281 ( .A(n_253), .Y(n_281) );
AND2x2_ASAP7_75t_L g309 ( .A(n_253), .B(n_310), .Y(n_309) );
NAND2x1_ASAP7_75t_L g358 ( .A(n_253), .B(n_254), .Y(n_358) );
INVx2_ASAP7_75t_L g379 ( .A(n_253), .Y(n_379) );
AND2x2_ASAP7_75t_L g398 ( .A(n_253), .B(n_254), .Y(n_398) );
INVx1_ASAP7_75t_L g501 ( .A(n_253), .Y(n_501) );
INVx1_ASAP7_75t_L g282 ( .A(n_254), .Y(n_282) );
INVx2_ASAP7_75t_L g310 ( .A(n_254), .Y(n_310) );
BUFx2_ASAP7_75t_L g361 ( .A(n_254), .Y(n_361) );
AND2x2_ASAP7_75t_L g378 ( .A(n_254), .B(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_254), .B(n_379), .Y(n_469) );
OR2x2_ASAP7_75t_L g481 ( .A(n_254), .B(n_281), .Y(n_481) );
OR2x6_ASAP7_75t_L g967 ( .A(n_255), .B(n_464), .Y(n_967) );
INVxp67_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g663 ( .A(n_256), .Y(n_663) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
BUFx2_ASAP7_75t_L g656 ( .A(n_257), .Y(n_656) );
AND2x4_ASAP7_75t_L g669 ( .A(n_257), .B(n_500), .Y(n_669) );
XNOR2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_725), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
XNOR2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_552), .Y(n_261) );
OAI22xp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_264), .B1(n_437), .B2(n_438), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVxp67_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
XNOR2x1_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
NOR2x1_ASAP7_75t_L g267 ( .A(n_268), .B(n_320), .Y(n_267) );
INVxp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_270), .A2(n_297), .B1(n_864), .B2(n_865), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_283), .Y(n_270) );
INVx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_272), .A2(n_306), .B1(n_503), .B2(n_504), .Y(n_502) );
AND2x4_ASAP7_75t_L g272 ( .A(n_273), .B(n_277), .Y(n_272) );
AND2x4_ASAP7_75t_L g306 ( .A(n_273), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVxp67_ASAP7_75t_L g319 ( .A(n_274), .Y(n_319) );
OR2x2_ASAP7_75t_L g498 ( .A(n_274), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g673 ( .A(n_274), .Y(n_673) );
BUFx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g293 ( .A(n_275), .Y(n_293) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
BUFx6f_ASAP7_75t_L g1056 ( .A(n_277), .Y(n_1056) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
AND2x2_ASAP7_75t_L g307 ( .A(n_278), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g390 ( .A(n_278), .B(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_SL g396 ( .A(n_278), .B(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_278), .B(n_329), .Y(n_450) );
BUFx2_ASAP7_75t_L g1014 ( .A(n_278), .Y(n_1014) );
AND2x4_ASAP7_75t_L g1045 ( .A(n_278), .B(n_1046), .Y(n_1045) );
AND2x4_ASAP7_75t_L g1059 ( .A(n_278), .B(n_308), .Y(n_1059) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_279), .Y(n_647) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_280), .Y(n_353) );
INVx3_ASAP7_75t_L g376 ( .A(n_280), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_280), .B(n_366), .Y(n_446) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_281), .Y(n_364) );
OR2x6_ASAP7_75t_L g283 ( .A(n_284), .B(n_290), .Y(n_283) );
OR2x2_ASAP7_75t_L g1100 ( .A(n_284), .B(n_290), .Y(n_1100) );
INVx2_ASAP7_75t_SL g1161 ( .A(n_284), .Y(n_1161) );
INVx2_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
INVx3_ASAP7_75t_L g414 ( .A(n_285), .Y(n_414) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx4f_ASAP7_75t_L g427 ( .A(n_286), .Y(n_427) );
BUFx3_ASAP7_75t_L g533 ( .A(n_286), .Y(n_533) );
BUFx3_ASAP7_75t_L g563 ( .A(n_286), .Y(n_563) );
OR2x4_ASAP7_75t_L g611 ( .A(n_286), .B(n_612), .Y(n_611) );
OR2x4_ASAP7_75t_L g634 ( .A(n_286), .B(n_316), .Y(n_634) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx2_ASAP7_75t_L g304 ( .A(n_287), .Y(n_304) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_287), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_287), .B(n_337), .Y(n_343) );
AND2x4_ASAP7_75t_L g436 ( .A(n_287), .B(n_336), .Y(n_436) );
INVx1_ASAP7_75t_L g314 ( .A(n_288), .Y(n_314) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVxp67_ASAP7_75t_L g303 ( .A(n_289), .Y(n_303) );
INVxp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g299 ( .A(n_291), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g340 ( .A(n_292), .B(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g344 ( .A(n_292), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g983 ( .A(n_292), .Y(n_983) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g489 ( .A(n_293), .Y(n_489) );
OR2x2_ASAP7_75t_L g558 ( .A(n_293), .B(n_547), .Y(n_558) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_293), .Y(n_641) );
INVx1_ASAP7_75t_L g529 ( .A(n_294), .Y(n_529) );
INVx3_ASAP7_75t_L g316 ( .A(n_295), .Y(n_316) );
BUFx3_ASAP7_75t_L g433 ( .A(n_295), .Y(n_433) );
NAND2xp33_ASAP7_75t_SL g547 ( .A(n_295), .B(n_318), .Y(n_547) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2x1_ASAP7_75t_L g297 ( .A(n_298), .B(n_305), .Y(n_297) );
INVx2_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g825 ( .A(n_300), .Y(n_825) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g914 ( .A(n_301), .Y(n_914) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_302), .Y(n_408) );
BUFx8_ASAP7_75t_L g424 ( .A(n_302), .Y(n_424) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_302), .Y(n_539) );
AND2x4_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
AND2x4_ASAP7_75t_L g313 ( .A(n_304), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_308), .Y(n_384) );
INVx1_ASAP7_75t_L g881 ( .A(n_308), .Y(n_881) );
INVx2_ASAP7_75t_L g1017 ( .A(n_308), .Y(n_1017) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx3_ASAP7_75t_L g371 ( .A(n_309), .Y(n_371) );
INVx2_ASAP7_75t_L g458 ( .A(n_309), .Y(n_458) );
AND2x4_ASAP7_75t_L g646 ( .A(n_309), .B(n_647), .Y(n_646) );
INVx3_ASAP7_75t_L g862 ( .A(n_311), .Y(n_862) );
INVx5_ASAP7_75t_L g1033 ( .A(n_311), .Y(n_1033) );
OR2x6_ASAP7_75t_L g311 ( .A(n_312), .B(n_319), .Y(n_311) );
NAND2x1p5_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
INVx8_ASAP7_75t_L g514 ( .A(n_313), .Y(n_514) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_313), .Y(n_520) );
BUFx3_ASAP7_75t_L g910 ( .A(n_313), .Y(n_910) );
BUFx3_ASAP7_75t_L g1088 ( .A(n_313), .Y(n_1088) );
AND2x4_ASAP7_75t_L g327 ( .A(n_315), .B(n_328), .Y(n_327) );
AND2x6_ASAP7_75t_L g508 ( .A(n_315), .B(n_324), .Y(n_508) );
AND2x2_ASAP7_75t_L g510 ( .A(n_315), .B(n_334), .Y(n_510) );
INVx1_ASAP7_75t_L g517 ( .A(n_315), .Y(n_517) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NAND3x1_ASAP7_75t_L g418 ( .A(n_316), .B(n_419), .C(n_420), .Y(n_418) );
NAND2x1p5_ASAP7_75t_L g535 ( .A(n_316), .B(n_420), .Y(n_535) );
INVx1_ASAP7_75t_L g612 ( .A(n_316), .Y(n_612) );
OR2x6_ASAP7_75t_L g614 ( .A(n_316), .B(n_572), .Y(n_614) );
AND2x4_ASAP7_75t_L g620 ( .A(n_316), .B(n_436), .Y(n_620) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND3x4_ASAP7_75t_L g432 ( .A(n_318), .B(n_402), .C(n_433), .Y(n_432) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_318), .Y(n_639) );
NAND3xp33_ASAP7_75t_SL g320 ( .A(n_321), .B(n_348), .C(n_404), .Y(n_320) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_330), .B1(n_331), .B2(n_338), .C(n_339), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2x1_ASAP7_75t_L g323 ( .A(n_324), .B(n_327), .Y(n_323) );
AND2x4_ASAP7_75t_SL g869 ( .A(n_324), .B(n_327), .Y(n_869) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_324), .B(n_327), .Y(n_1097) );
INVx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2x1p5_ASAP7_75t_L g346 ( .A(n_326), .B(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g410 ( .A(n_326), .B(n_335), .Y(n_410) );
BUFx2_ASAP7_75t_L g625 ( .A(n_326), .Y(n_625) );
AND2x4_ASAP7_75t_L g331 ( .A(n_327), .B(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g434 ( .A(n_327), .B(n_435), .Y(n_434) );
AND2x4_ASAP7_75t_SL g871 ( .A(n_327), .B(n_332), .Y(n_871) );
OR2x2_ASAP7_75t_L g445 ( .A(n_328), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g419 ( .A(n_329), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_330), .A2(n_360), .B1(n_362), .B2(n_363), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_331), .A2(n_1096), .B1(n_1097), .B2(n_1098), .Y(n_1095) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g347 ( .A(n_337), .Y(n_347) );
INVx1_ASAP7_75t_L g874 ( .A(n_340), .Y(n_874) );
AND2x4_ASAP7_75t_L g1078 ( .A(n_340), .B(n_445), .Y(n_1078) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_342), .Y(n_542) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx2_ASAP7_75t_L g572 ( .A(n_343), .Y(n_572) );
INVx2_ASAP7_75t_L g876 ( .A(n_344), .Y(n_876) );
AND2x4_ASAP7_75t_L g1081 ( .A(n_344), .B(n_498), .Y(n_1081) );
INVx4_ASAP7_75t_L g416 ( .A(n_345), .Y(n_416) );
INVx3_ASAP7_75t_L g430 ( .A(n_345), .Y(n_430) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g566 ( .A(n_346), .Y(n_566) );
BUFx2_ASAP7_75t_L g618 ( .A(n_346), .Y(n_618) );
BUFx2_ASAP7_75t_L g629 ( .A(n_347), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_388), .B(n_399), .Y(n_348) );
NAND3xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_367), .C(n_380), .Y(n_349) );
A2O1A1Ixp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_352), .B(n_354), .C(n_365), .Y(n_350) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx3_ASAP7_75t_L g1007 ( .A(n_353), .Y(n_1007) );
A2O1A1Ixp33_ASAP7_75t_L g1019 ( .A1(n_353), .A2(n_365), .B(n_985), .C(n_1020), .Y(n_1019) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_355), .B(n_359), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g368 ( .A(n_356), .Y(n_368) );
INVx2_ASAP7_75t_L g382 ( .A(n_356), .Y(n_382) );
INVx4_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx4f_ASAP7_75t_L g482 ( .A(n_357), .Y(n_482) );
OR2x6_ASAP7_75t_L g490 ( .A(n_357), .B(n_491), .Y(n_490) );
BUFx4f_ASAP7_75t_L g660 ( .A(n_357), .Y(n_660) );
BUFx4f_ASAP7_75t_L g696 ( .A(n_357), .Y(n_696) );
BUFx4f_ASAP7_75t_L g969 ( .A(n_357), .Y(n_969) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx3_ASAP7_75t_L g452 ( .A(n_358), .Y(n_452) );
BUFx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g497 ( .A(n_361), .Y(n_497) );
AND2x4_ASAP7_75t_L g666 ( .A(n_361), .B(n_656), .Y(n_666) );
AND2x2_ASAP7_75t_L g751 ( .A(n_361), .B(n_656), .Y(n_751) );
INVx1_ASAP7_75t_L g889 ( .A(n_361), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_361), .A2(n_363), .B1(n_980), .B2(n_1002), .Y(n_1021) );
AOI221xp5_ASAP7_75t_L g887 ( .A1(n_363), .A2(n_875), .B1(n_888), .B2(n_890), .C(n_891), .Y(n_887) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g893 ( .A(n_365), .Y(n_893) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_366), .B(n_403), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_366), .B(n_500), .Y(n_499) );
AND2x6_ASAP7_75t_L g1053 ( .A(n_366), .B(n_397), .Y(n_1053) );
INVx1_ASAP7_75t_L g1065 ( .A(n_366), .Y(n_1065) );
OAI211xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_369), .B(n_370), .C(n_374), .Y(n_367) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI221xp5_ASAP7_75t_L g1008 ( .A1(n_373), .A2(n_382), .B1(n_1009), .B2(n_1010), .C(n_1011), .Y(n_1008) );
INVx3_ASAP7_75t_L g1073 ( .A(n_373), .Y(n_1073) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g485 ( .A(n_376), .Y(n_485) );
INVx2_ASAP7_75t_L g883 ( .A(n_376), .Y(n_883) );
INVx2_ASAP7_75t_SL g886 ( .A(n_376), .Y(n_886) );
BUFx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g392 ( .A(n_378), .Y(n_392) );
BUFx3_ASAP7_75t_L g898 ( .A(n_378), .Y(n_898) );
BUFx6f_ASAP7_75t_L g1046 ( .A(n_378), .Y(n_1046) );
OAI211xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B(n_383), .C(n_387), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_381), .A2(n_412), .B1(n_413), .B2(n_415), .Y(n_411) );
INVx4_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g487 ( .A(n_386), .B(n_488), .Y(n_487) );
OAI21xp33_ASAP7_75t_L g1024 ( .A1(n_386), .A2(n_599), .B(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_SL g1051 ( .A(n_386), .Y(n_1051) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_386), .B(n_488), .Y(n_1145) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_390), .A2(n_861), .B1(n_900), .B2(n_901), .Y(n_899) );
AND2x4_ASAP7_75t_L g448 ( .A(n_391), .B(n_449), .Y(n_448) );
INVx3_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g1061 ( .A(n_394), .Y(n_1061) );
INVx4_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx3_ASAP7_75t_L g901 ( .A(n_396), .Y(n_901) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_397), .Y(n_460) );
AND2x2_ASAP7_75t_L g662 ( .A(n_397), .B(n_663), .Y(n_662) );
BUFx3_ASAP7_75t_L g1023 ( .A(n_397), .Y(n_1023) );
BUFx3_ASAP7_75t_L g1049 ( .A(n_397), .Y(n_1049) );
INVx1_ASAP7_75t_L g1072 ( .A(n_397), .Y(n_1072) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g847 ( .A(n_398), .Y(n_847) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g1075 ( .A(n_400), .Y(n_1075) );
BUFx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OAI31xp33_ASAP7_75t_L g1004 ( .A1(n_401), .A2(n_1005), .A3(n_1012), .B(n_1022), .Y(n_1004) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx2_ASAP7_75t_L g474 ( .A(n_403), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_417), .B1(n_421), .B2(n_431), .C(n_434), .Y(n_404) );
INVx2_ASAP7_75t_L g569 ( .A(n_406), .Y(n_569) );
INVx1_ASAP7_75t_L g1378 ( .A(n_406), .Y(n_1378) );
INVx8_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g790 ( .A1(n_407), .A2(n_773), .B1(n_781), .B2(n_787), .Y(n_790) );
BUFx3_ASAP7_75t_L g1390 ( .A(n_407), .Y(n_1390) );
INVx5_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx3_ASAP7_75t_L g522 ( .A(n_408), .Y(n_522) );
INVx2_ASAP7_75t_SL g992 ( .A(n_408), .Y(n_992) );
HB1xp67_ASAP7_75t_L g1158 ( .A(n_408), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_409), .A2(n_524), .B1(n_525), .B2(n_526), .Y(n_523) );
BUFx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx12f_ASAP7_75t_L g915 ( .A(n_410), .Y(n_915) );
BUFx3_ASAP7_75t_L g993 ( .A(n_410), .Y(n_993) );
INVx5_ASAP7_75t_L g1092 ( .A(n_410), .Y(n_1092) );
BUFx4f_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
OAI22xp33_ASAP7_75t_L g941 ( .A1(n_414), .A2(n_928), .B1(n_934), .B2(n_942), .Y(n_941) );
OAI22xp33_ASAP7_75t_L g946 ( .A1(n_414), .A2(n_929), .B1(n_935), .B2(n_947), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g1380 ( .A1(n_414), .A2(n_690), .B1(n_1381), .B2(n_1382), .Y(n_1380) );
OAI22xp33_ASAP7_75t_L g794 ( .A1(n_415), .A2(n_561), .B1(n_767), .B2(n_777), .Y(n_794) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g532 ( .A(n_416), .Y(n_532) );
INVx1_ASAP7_75t_L g785 ( .A(n_416), .Y(n_785) );
INVx1_ASAP7_75t_L g830 ( .A(n_416), .Y(n_830) );
INVx1_ASAP7_75t_L g942 ( .A(n_416), .Y(n_942) );
INVx2_ASAP7_75t_L g581 ( .A(n_417), .Y(n_581) );
NAND3xp33_ASAP7_75t_L g912 ( .A(n_417), .B(n_913), .C(n_916), .Y(n_912) );
CKINVDCx5p33_ASAP7_75t_R g1388 ( .A(n_417), .Y(n_1388) );
INVx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx3_ASAP7_75t_L g793 ( .A(n_418), .Y(n_793) );
OAI33xp33_ASAP7_75t_L g819 ( .A1(n_418), .A2(n_783), .A3(n_820), .B1(n_824), .B2(n_826), .B3(n_829), .Y(n_819) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx3_ASAP7_75t_L g686 ( .A(n_424), .Y(n_686) );
AND2x4_ASAP7_75t_L g999 ( .A(n_424), .B(n_983), .Y(n_999) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B1(n_428), .B2(n_429), .Y(n_425) );
INVx1_ASAP7_75t_L g1152 ( .A(n_427), .Y(n_1152) );
OAI211xp5_ASAP7_75t_L g544 ( .A1(n_429), .A2(n_478), .B(n_545), .C(n_548), .Y(n_544) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_429), .Y(n_737) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx3_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AOI33xp33_ASAP7_75t_L g986 ( .A1(n_432), .A2(n_987), .A3(n_989), .B1(n_990), .B2(n_994), .B3(n_996), .Y(n_986) );
AOI33xp33_ASAP7_75t_L g1084 ( .A1(n_432), .A2(n_996), .A3(n_1085), .B1(n_1090), .B2(n_1093), .B3(n_1094), .Y(n_1084) );
INVx3_ASAP7_75t_L g624 ( .A(n_433), .Y(n_624) );
INVx3_ASAP7_75t_L g911 ( .A(n_434), .Y(n_911) );
AOI221xp5_ASAP7_75t_L g1001 ( .A1(n_434), .A2(n_869), .B1(n_871), .B2(n_1002), .C(n_1003), .Y(n_1001) );
BUFx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx3_ASAP7_75t_L g515 ( .A(n_436), .Y(n_515) );
BUFx2_ASAP7_75t_L g526 ( .A(n_436), .Y(n_526) );
INVx2_ASAP7_75t_L g918 ( .A(n_436), .Y(n_918) );
BUFx2_ASAP7_75t_L g1089 ( .A(n_436), .Y(n_1089) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
XNOR2x1_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
NAND4xp75_ASAP7_75t_L g441 ( .A(n_442), .B(n_453), .C(n_502), .D(n_505), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g451 ( .A(n_450), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_SL g596 ( .A(n_452), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_452), .B(n_1021), .Y(n_1020) );
BUFx2_ASAP7_75t_SL g1399 ( .A(n_452), .Y(n_1399) );
AOI211x1_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_471), .B(n_476), .C(n_494), .Y(n_453) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g1050 ( .A(n_456), .Y(n_1050) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AOI221xp5_ASAP7_75t_L g1015 ( .A1(n_460), .A2(n_998), .B1(n_1003), .B2(n_1016), .C(n_1018), .Y(n_1015) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B1(n_465), .B2(n_470), .Y(n_461) );
INVx1_ASAP7_75t_L g1133 ( .A(n_463), .Y(n_1133) );
BUFx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx3_ASAP7_75t_L g766 ( .A(n_464), .Y(n_766) );
INVx2_ASAP7_75t_SL g816 ( .A(n_464), .Y(n_816) );
OAI22xp33_ASAP7_75t_L g927 ( .A1(n_465), .A2(n_779), .B1(n_928), .B2(n_929), .Y(n_927) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_467), .Y(n_589) );
INVx1_ASAP7_75t_L g607 ( .A(n_467), .Y(n_607) );
INVx2_ASAP7_75t_L g768 ( .A(n_467), .Y(n_768) );
INVx2_ASAP7_75t_SL g806 ( .A(n_467), .Y(n_806) );
INVx4_ASAP7_75t_L g1030 ( .A(n_467), .Y(n_1030) );
INVx1_ASAP7_75t_L g1395 ( .A(n_467), .Y(n_1395) );
INVx8_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OR2x2_ASAP7_75t_L g655 ( .A(n_468), .B(n_656), .Y(n_655) );
BUFx2_ASAP7_75t_L g1068 ( .A(n_468), .Y(n_1068) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OAI221xp5_ASAP7_75t_L g531 ( .A1(n_470), .A2(n_483), .B1(n_532), .B2(n_533), .C(n_534), .Y(n_531) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OAI33xp33_ASAP7_75t_L g1393 ( .A1(n_472), .A2(n_600), .A3(n_1394), .B1(n_1396), .B2(n_1397), .B3(n_1400), .Y(n_1393) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g583 ( .A(n_473), .Y(n_583) );
INVx4_ASAP7_75t_L g763 ( .A(n_473), .Y(n_763) );
INVx2_ASAP7_75t_L g800 ( .A(n_473), .Y(n_800) );
INVx2_ASAP7_75t_L g1129 ( .A(n_473), .Y(n_1129) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g551 ( .A(n_474), .Y(n_551) );
OR2x6_ASAP7_75t_L g948 ( .A(n_474), .B(n_535), .Y(n_948) );
OAI21xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_486), .B(n_490), .Y(n_476) );
OAI221xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B1(n_482), .B2(n_483), .C(n_484), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_479), .A2(n_595), .B1(n_812), .B2(n_813), .Y(n_811) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g594 ( .A(n_481), .Y(n_594) );
BUFx3_ASAP7_75t_L g599 ( .A(n_481), .Y(n_599) );
BUFx2_ASAP7_75t_L g700 ( .A(n_481), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_482), .A2(n_775), .B1(n_776), .B2(n_777), .Y(n_774) );
OAI33xp33_ASAP7_75t_L g760 ( .A1(n_486), .A2(n_761), .A3(n_764), .B1(n_769), .B2(n_774), .B3(n_778), .Y(n_760) );
OAI33xp33_ASAP7_75t_L g798 ( .A1(n_486), .A2(n_799), .A3(n_801), .B1(n_807), .B2(n_811), .B3(n_814), .Y(n_798) );
OAI33xp33_ASAP7_75t_L g926 ( .A1(n_486), .A2(n_761), .A3(n_927), .B1(n_930), .B2(n_933), .B3(n_936), .Y(n_926) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g600 ( .A(n_487), .Y(n_600) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2x2_ASAP7_75t_L g495 ( .A(n_492), .B(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_503), .A2(n_504), .B1(n_520), .B2(n_521), .Y(n_519) );
OAI31xp67_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_518), .A3(n_530), .B(n_550), .Y(n_505) );
INVx4_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B(n_515), .C(n_516), .Y(n_511) );
CKINVDCx5p33_ASAP7_75t_R g513 ( .A(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g549 ( .A(n_514), .Y(n_549) );
INVx2_ASAP7_75t_L g982 ( .A(n_514), .Y(n_982) );
INVx8_ASAP7_75t_L g988 ( .A(n_514), .Y(n_988) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AOI21xp33_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_523), .B(n_527), .Y(n_518) );
INVx2_ASAP7_75t_L g575 ( .A(n_521), .Y(n_575) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
OAI21xp5_ASAP7_75t_SL g530 ( .A1(n_531), .A2(n_536), .B(n_544), .Y(n_530) );
OAI22xp33_ASAP7_75t_L g1385 ( .A1(n_533), .A2(n_690), .B1(n_1386), .B2(n_1387), .Y(n_1385) );
INVx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_540), .B1(n_541), .B2(n_543), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_537), .A2(n_770), .B1(n_780), .B2(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x4_ASAP7_75t_L g636 ( .A(n_539), .B(n_612), .Y(n_636) );
BUFx6f_ASAP7_75t_L g828 ( .A(n_539), .Y(n_828) );
INVx2_ASAP7_75t_L g904 ( .A(n_539), .Y(n_904) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_541), .A2(n_808), .B1(n_817), .B2(n_825), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_541), .A2(n_904), .B1(n_932), .B2(n_939), .Y(n_949) );
CKINVDCx8_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
INVx3_ASAP7_75t_L g577 ( .A(n_542), .Y(n_577) );
INVx3_ASAP7_75t_L g945 ( .A(n_542), .Y(n_945) );
INVx3_ASAP7_75t_L g1155 ( .A(n_542), .Y(n_1155) );
BUFx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AOI31xp33_ASAP7_75t_L g877 ( .A1(n_550), .A2(n_878), .A3(n_894), .B(n_899), .Y(n_877) );
BUFx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
XOR2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_674), .Y(n_552) );
AND3x1_ASAP7_75t_L g554 ( .A(n_555), .B(n_608), .C(n_642), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_582), .Y(n_555) );
OAI33xp33_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_559), .A3(n_567), .B1(n_573), .B2(n_578), .B3(n_581), .Y(n_556) );
OAI33xp33_ASAP7_75t_L g677 ( .A1(n_557), .A2(n_581), .A3(n_678), .B1(n_681), .B2(n_684), .B3(n_688), .Y(n_677) );
OAI211xp5_ASAP7_75t_SL g902 ( .A1(n_557), .A2(n_903), .B(n_911), .C(n_912), .Y(n_902) );
OAI33xp33_ASAP7_75t_L g1149 ( .A1(n_557), .A2(n_581), .A3(n_1150), .B1(n_1153), .B2(n_1156), .B3(n_1159), .Y(n_1149) );
BUFx4f_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx8_ASAP7_75t_L g783 ( .A(n_558), .Y(n_783) );
BUFx4f_ASAP7_75t_L g1384 ( .A(n_558), .Y(n_1384) );
OAI22xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B1(n_564), .B2(n_565), .Y(n_559) );
OAI22xp33_ASAP7_75t_L g584 ( .A1(n_560), .A2(n_579), .B1(n_585), .B2(n_588), .Y(n_584) );
OAI22xp33_ASAP7_75t_L g578 ( .A1(n_561), .A2(n_565), .B1(n_579), .B2(n_580), .Y(n_578) );
OAI22xp33_ASAP7_75t_L g678 ( .A1(n_561), .A2(n_565), .B1(n_679), .B2(n_680), .Y(n_678) );
OAI22xp33_ASAP7_75t_L g688 ( .A1(n_561), .A2(n_689), .B1(n_690), .B2(n_692), .Y(n_688) );
OAI22xp33_ASAP7_75t_L g784 ( .A1(n_561), .A2(n_765), .B1(n_776), .B2(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g822 ( .A(n_563), .Y(n_822) );
OAI22xp33_ASAP7_75t_L g597 ( .A1(n_564), .A2(n_580), .B1(n_595), .B2(n_598), .Y(n_597) );
OAI22xp33_ASAP7_75t_L g1159 ( .A1(n_565), .A2(n_1134), .B1(n_1142), .B2(n_1160), .Y(n_1159) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g691 ( .A(n_566), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B1(n_570), .B2(n_571), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_568), .A2(n_574), .B1(n_591), .B2(n_595), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_569), .A2(n_571), .B1(n_682), .B2(n_683), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_570), .A2(n_576), .B1(n_602), .B2(n_606), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g1389 ( .A1(n_571), .A2(n_1390), .B1(n_1391), .B2(n_1392), .Y(n_1389) );
BUFx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g789 ( .A(n_572), .Y(n_789) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_575), .B1(n_576), .B2(n_577), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_577), .A2(n_685), .B1(n_686), .B2(n_687), .Y(n_684) );
OAI33xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .A3(n_590), .B1(n_597), .B2(n_600), .B3(n_601), .Y(n_582) );
OAI33xp33_ASAP7_75t_L g693 ( .A1(n_583), .A2(n_600), .A3(n_694), .B1(n_695), .B2(n_697), .B3(n_701), .Y(n_693) );
OAI22xp33_ASAP7_75t_L g694 ( .A1(n_585), .A2(n_588), .B1(n_679), .B2(n_689), .Y(n_694) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx3_ASAP7_75t_L g938 ( .A(n_586), .Y(n_938) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx4_ASAP7_75t_L g1028 ( .A(n_587), .Y(n_1028) );
OAI22xp5_ASAP7_75t_L g1400 ( .A1(n_588), .A2(n_766), .B1(n_1379), .B2(n_1392), .Y(n_1400) );
INVx6_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx5_ASAP7_75t_L g702 ( .A(n_589), .Y(n_702) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g1137 ( .A1(n_593), .A2(n_969), .B1(n_1138), .B2(n_1139), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g1140 ( .A1(n_593), .A2(n_595), .B1(n_1141), .B2(n_1142), .Y(n_1140) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g1011 ( .A(n_594), .Y(n_1011) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_595), .A2(n_680), .B1(n_692), .B2(n_698), .Y(n_697) );
OAI211xp5_ASAP7_75t_L g894 ( .A1(n_595), .A2(n_895), .B(n_896), .C(n_897), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_595), .A2(n_775), .B1(n_931), .B2(n_932), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g1396 ( .A1(n_595), .A2(n_775), .B1(n_1377), .B2(n_1391), .Y(n_1396) );
INVx5_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_599), .A2(n_682), .B1(n_685), .B2(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g772 ( .A(n_599), .Y(n_772) );
OAI22xp33_ASAP7_75t_L g701 ( .A1(n_602), .A2(n_683), .B1(n_687), .B2(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx3_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OAI31xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_615), .A3(n_631), .B(n_637), .Y(n_608) );
BUFx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_SL g713 ( .A(n_611), .Y(n_713) );
BUFx3_ASAP7_75t_L g744 ( .A(n_611), .Y(n_744) );
BUFx2_ASAP7_75t_L g1125 ( .A(n_611), .Y(n_1125) );
BUFx3_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g746 ( .A(n_614), .Y(n_746) );
INVx1_ASAP7_75t_L g840 ( .A(n_614), .Y(n_840) );
INVx2_ASAP7_75t_L g961 ( .A(n_614), .Y(n_961) );
INVxp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g947 ( .A(n_617), .Y(n_947) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g707 ( .A(n_618), .Y(n_707) );
CKINVDCx8_ASAP7_75t_R g619 ( .A(n_620), .Y(n_619) );
CKINVDCx8_ASAP7_75t_R g738 ( .A(n_620), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_626), .B1(n_627), .B2(n_630), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_622), .A2(n_627), .B1(n_709), .B2(n_710), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_622), .A2(n_627), .B1(n_1115), .B2(n_1123), .Y(n_1122) );
BUFx3_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
BUFx3_ASAP7_75t_L g740 ( .A(n_623), .Y(n_740) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
AND2x4_ASAP7_75t_L g628 ( .A(n_624), .B(n_629), .Y(n_628) );
AND2x4_ASAP7_75t_L g835 ( .A(n_624), .B(n_625), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_626), .A2(n_665), .B1(n_667), .B2(n_670), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g1404 ( .A1(n_627), .A2(n_740), .B1(n_1405), .B2(n_1406), .Y(n_1404) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_SL g739 ( .A1(n_628), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_628), .A2(n_835), .B1(n_836), .B2(n_837), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_628), .A2(n_835), .B1(n_957), .B2(n_958), .Y(n_956) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_634), .Y(n_715) );
INVx2_ASAP7_75t_SL g734 ( .A(n_634), .Y(n_734) );
INVx1_ASAP7_75t_L g953 ( .A(n_634), .Y(n_953) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g716 ( .A(n_636), .Y(n_716) );
INVx2_ASAP7_75t_L g735 ( .A(n_636), .Y(n_735) );
INVxp67_ASAP7_75t_L g954 ( .A(n_636), .Y(n_954) );
OAI31xp33_ASAP7_75t_L g831 ( .A1(n_637), .A2(n_832), .A3(n_833), .B(n_838), .Y(n_831) );
OAI31xp33_ASAP7_75t_L g1401 ( .A1(n_637), .A2(n_1402), .A3(n_1403), .B(n_1407), .Y(n_1401) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
AND2x4_ASAP7_75t_L g717 ( .A(n_638), .B(n_640), .Y(n_717) );
AND2x2_ASAP7_75t_L g962 ( .A(n_638), .B(n_640), .Y(n_962) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OAI31xp33_ASAP7_75t_SL g642 ( .A1(n_643), .A2(n_648), .A3(n_657), .B(n_671), .Y(n_642) );
INVx3_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
CKINVDCx16_ASAP7_75t_R g720 ( .A(n_646), .Y(n_720) );
INVx4_ASAP7_75t_L g758 ( .A(n_646), .Y(n_758) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
BUFx2_ASAP7_75t_L g754 ( .A(n_651), .Y(n_754) );
BUFx6f_ASAP7_75t_L g853 ( .A(n_651), .Y(n_853) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx2_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
BUFx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g756 ( .A(n_655), .Y(n_756) );
INVx1_ASAP7_75t_L g1111 ( .A(n_655), .Y(n_1111) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_660), .A2(n_770), .B1(n_771), .B2(n_773), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_660), .A2(n_808), .B1(n_809), .B2(n_810), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g933 ( .A1(n_660), .A2(n_809), .B1(n_934), .B2(n_935), .Y(n_933) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g749 ( .A(n_662), .Y(n_749) );
INVx3_ASAP7_75t_L g1118 ( .A(n_662), .Y(n_1118) );
AND2x2_ASAP7_75t_L g845 ( .A(n_663), .B(n_846), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_665), .A2(n_667), .B1(n_709), .B2(n_724), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_665), .A2(n_1115), .B1(n_1116), .B2(n_1117), .Y(n_1114) );
BUFx3_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_666), .A2(n_669), .B1(n_957), .B2(n_971), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_667), .A2(n_741), .B1(n_751), .B2(n_752), .Y(n_750) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g850 ( .A(n_669), .Y(n_850) );
BUFx3_ASAP7_75t_L g1116 ( .A(n_669), .Y(n_1116) );
OAI31xp33_ASAP7_75t_L g718 ( .A1(n_671), .A2(n_719), .A3(n_721), .B(n_722), .Y(n_718) );
OAI31xp33_ASAP7_75t_L g747 ( .A1(n_671), .A2(n_748), .A3(n_753), .B(n_757), .Y(n_747) );
BUFx2_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
BUFx3_ASAP7_75t_L g855 ( .A(n_672), .Y(n_855) );
BUFx2_ASAP7_75t_L g974 ( .A(n_672), .Y(n_974) );
INVx1_ASAP7_75t_L g1105 ( .A(n_672), .Y(n_1105) );
AND3x1_ASAP7_75t_L g675 ( .A(n_676), .B(n_703), .C(n_718), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_693), .Y(n_676) );
OAI22xp33_ASAP7_75t_L g1150 ( .A1(n_690), .A2(n_1131), .B1(n_1141), .B2(n_1151), .Y(n_1150) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx4_ASAP7_75t_L g775 ( .A(n_699), .Y(n_775) );
INVx2_ASAP7_75t_L g809 ( .A(n_699), .Y(n_809) );
INVx2_ASAP7_75t_L g1398 ( .A(n_699), .Y(n_1398) );
INVx4_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_702), .A2(n_779), .B1(n_780), .B2(n_781), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_702), .A2(n_815), .B1(n_817), .B2(n_818), .Y(n_814) );
OAI31xp33_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_711), .A3(n_714), .B(n_717), .Y(n_703) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVxp67_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g823 ( .A(n_707), .Y(n_823) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
OAI31xp33_ASAP7_75t_L g731 ( .A1(n_717), .A2(n_732), .A3(n_736), .B(n_743), .Y(n_731) );
CKINVDCx14_ASAP7_75t_R g1126 ( .A(n_717), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_1036), .B1(n_1037), .B2(n_1162), .Y(n_725) );
INVx1_ASAP7_75t_L g1162 ( .A(n_726), .Y(n_1162) );
XNOR2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_856), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
XNOR2x1_ASAP7_75t_L g728 ( .A(n_729), .B(n_795), .Y(n_728) );
NAND3xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_747), .C(n_759), .Y(n_730) );
INVx2_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_751), .A2(n_836), .B1(n_849), .B2(n_851), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g1411 ( .A1(n_751), .A2(n_849), .B1(n_1405), .B2(n_1412), .Y(n_1411) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g854 ( .A(n_756), .Y(n_854) );
INVx1_ASAP7_75t_L g973 ( .A(n_756), .Y(n_973) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_782), .Y(n_759) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
OAI22xp33_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B1(n_767), .B2(n_768), .Y(n_764) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_768), .A2(n_937), .B1(n_938), .B2(n_939), .Y(n_936) );
INVx3_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
OAI22xp33_ASAP7_75t_L g1394 ( .A1(n_779), .A2(n_1381), .B1(n_1386), .B2(n_1395), .Y(n_1394) );
OAI33xp33_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_784), .A3(n_786), .B1(n_790), .B2(n_791), .B3(n_794), .Y(n_782) );
OAI33xp33_ASAP7_75t_L g940 ( .A1(n_783), .A2(n_941), .A3(n_943), .B1(n_946), .B2(n_948), .B3(n_949), .Y(n_940) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_787), .A2(n_810), .B1(n_818), .B2(n_827), .Y(n_826) );
OAI221xp5_ASAP7_75t_L g903 ( .A1(n_787), .A2(n_904), .B1(n_905), .B2(n_906), .C(n_907), .Y(n_903) );
OAI22xp33_ASAP7_75t_SL g1376 ( .A1(n_787), .A2(n_1377), .B1(n_1378), .B2(n_1379), .Y(n_1376) );
INVx3_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
BUFx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
BUFx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NAND3xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_831), .C(n_841), .Y(n_796) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_798), .B(n_819), .Y(n_797) );
BUFx6f_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
OAI22xp33_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_803), .B1(n_805), .B2(n_806), .Y(n_801) );
OAI22xp33_ASAP7_75t_L g820 ( .A1(n_802), .A2(n_812), .B1(n_821), .B2(n_823), .Y(n_820) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
OAI22xp33_ASAP7_75t_L g829 ( .A1(n_805), .A2(n_813), .B1(n_821), .B2(n_830), .Y(n_829) );
OAI221xp5_ASAP7_75t_L g1066 ( .A1(n_815), .A2(n_1067), .B1(n_1068), .B2(n_1069), .C(n_1070), .Y(n_1066) );
INVx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g944 ( .A(n_828), .Y(n_944) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
OAI31xp33_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_843), .A3(n_852), .B(n_855), .Y(n_841) );
INVx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
BUFx2_ASAP7_75t_L g892 ( .A(n_847), .Y(n_892) );
INVx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
OAI31xp33_ASAP7_75t_L g1408 ( .A1(n_855), .A2(n_1409), .A3(n_1410), .B(n_1413), .Y(n_1408) );
XNOR2xp5_ASAP7_75t_L g856 ( .A(n_857), .B(n_921), .Y(n_856) );
HB1xp67_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g919 ( .A(n_859), .Y(n_919) );
NAND3xp33_ASAP7_75t_L g859 ( .A(n_860), .B(n_863), .C(n_866), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_861), .B(n_862), .Y(n_860) );
NOR3xp33_ASAP7_75t_SL g866 ( .A(n_867), .B(n_877), .C(n_902), .Y(n_866) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_873), .A2(n_874), .B1(n_875), .B2(n_876), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_873), .B(n_886), .Y(n_885) );
AOI222xp33_ASAP7_75t_L g979 ( .A1(n_874), .A2(n_876), .B1(n_980), .B2(n_981), .C1(n_984), .C2(n_985), .Y(n_979) );
AOI21xp5_ASAP7_75t_L g878 ( .A1(n_879), .A2(n_882), .B(n_884), .Y(n_878) );
INVx2_ASAP7_75t_SL g880 ( .A(n_881), .Y(n_880) );
AOI21xp5_ASAP7_75t_L g884 ( .A1(n_885), .A2(n_887), .B(n_893), .Y(n_884) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
NOR2x1_ASAP7_75t_L g1064 ( .A(n_889), .B(n_1065), .Y(n_1064) );
INVx2_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx2_ASAP7_75t_SL g1102 ( .A(n_911), .Y(n_1102) );
INVx1_ASAP7_75t_L g1154 ( .A(n_914), .Y(n_1154) );
INVx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g995 ( .A(n_918), .Y(n_995) );
AOI22xp5_ASAP7_75t_L g921 ( .A1(n_922), .A2(n_923), .B1(n_975), .B2(n_1035), .Y(n_921) );
INVx2_ASAP7_75t_SL g922 ( .A(n_923), .Y(n_922) );
NAND3xp33_ASAP7_75t_L g924 ( .A(n_925), .B(n_950), .C(n_963), .Y(n_924) );
NOR2xp33_ASAP7_75t_L g925 ( .A(n_926), .B(n_940), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_931), .A2(n_937), .B1(n_944), .B2(n_945), .Y(n_943) );
OAI22xp5_ASAP7_75t_L g1156 ( .A1(n_945), .A2(n_1139), .B1(n_1148), .B2(n_1157), .Y(n_1156) );
INVx1_ASAP7_75t_L g996 ( .A(n_948), .Y(n_996) );
OAI31xp33_ASAP7_75t_L g950 ( .A1(n_951), .A2(n_955), .A3(n_959), .B(n_962), .Y(n_950) );
INVx1_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
INVx2_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
OAI31xp33_ASAP7_75t_SL g963 ( .A1(n_964), .A2(n_968), .A3(n_972), .B(n_974), .Y(n_963) );
INVx1_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
HB1xp67_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
INVx1_ASAP7_75t_L g1035 ( .A(n_976), .Y(n_1035) );
XNOR2x1_ASAP7_75t_L g976 ( .A(n_977), .B(n_1034), .Y(n_976) );
OR2x2_ASAP7_75t_L g977 ( .A(n_978), .B(n_1000), .Y(n_977) );
NAND3xp33_ASAP7_75t_L g978 ( .A(n_979), .B(n_986), .C(n_997), .Y(n_978) );
AND2x4_ASAP7_75t_L g981 ( .A(n_982), .B(n_983), .Y(n_981) );
INVx2_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_998), .B(n_999), .Y(n_997) );
INVx2_ASAP7_75t_L g1101 ( .A(n_999), .Y(n_1101) );
NAND3xp33_ASAP7_75t_SL g1000 ( .A(n_1001), .B(n_1004), .C(n_1031), .Y(n_1000) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
OAI21xp33_ASAP7_75t_L g1012 ( .A1(n_1013), .A2(n_1015), .B(n_1019), .Y(n_1012) );
INVxp67_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
INVx2_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_1027), .A2(n_1028), .B1(n_1029), .B2(n_1030), .Y(n_1026) );
INVx2_ASAP7_75t_L g1136 ( .A(n_1030), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1033), .Y(n_1031) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
XNOR2xp5_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1103), .Y(n_1039) );
NAND3xp33_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1076), .C(n_1082), .Y(n_1041) );
OAI21xp33_ASAP7_75t_L g1042 ( .A1(n_1043), .A2(n_1060), .B(n_1074), .Y(n_1042) );
INVx2_ASAP7_75t_SL g1044 ( .A(n_1045), .Y(n_1044) );
AOI21xp5_ASAP7_75t_SL g1047 ( .A1(n_1048), .A2(n_1052), .B(n_1053), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_1055), .A2(n_1056), .B1(n_1057), .B2(n_1058), .Y(n_1054) );
HB1xp67_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
BUFx2_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
INVx2_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
AOI21xp33_ASAP7_75t_SL g1076 ( .A1(n_1077), .A2(n_1079), .B(n_1080), .Y(n_1076) );
INVx8_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
NOR3xp33_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1099), .C(n_1102), .Y(n_1082) );
NAND2xp5_ASAP7_75t_SL g1083 ( .A(n_1084), .B(n_1095), .Y(n_1083) );
INVx2_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
INVx2_ASAP7_75t_SL g1087 ( .A(n_1088), .Y(n_1087) );
INVx2_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
OAI221xp5_ASAP7_75t_L g1104 ( .A1(n_1105), .A2(n_1106), .B1(n_1119), .B2(n_1126), .C(n_1127), .Y(n_1104) );
NOR3xp33_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1112), .C(n_1113), .Y(n_1106) );
INVx2_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
INVx2_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
INVx2_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
NOR3xp33_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1121), .C(n_1124), .Y(n_1119) );
NOR2xp33_ASAP7_75t_L g1127 ( .A(n_1128), .B(n_1149), .Y(n_1127) );
OAI33xp33_ASAP7_75t_L g1128 ( .A1(n_1129), .A2(n_1130), .A3(n_1137), .B1(n_1140), .B2(n_1143), .B3(n_1146), .Y(n_1128) );
OAI22xp5_ASAP7_75t_L g1130 ( .A1(n_1131), .A2(n_1132), .B1(n_1134), .B2(n_1135), .Y(n_1130) );
OAI22xp5_ASAP7_75t_L g1146 ( .A1(n_1132), .A2(n_1135), .B1(n_1147), .B2(n_1148), .Y(n_1146) );
INVx2_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
INVx2_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
OAI22xp5_ASAP7_75t_L g1153 ( .A1(n_1138), .A2(n_1147), .B1(n_1154), .B2(n_1155), .Y(n_1153) );
INVx2_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
INVx2_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
OAI221xp5_ASAP7_75t_L g1163 ( .A1(n_1164), .A2(n_1367), .B1(n_1369), .B2(n_1414), .C(n_1417), .Y(n_1163) );
NOR2xp67_ASAP7_75t_SL g1164 ( .A(n_1165), .B(n_1305), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1266), .Y(n_1165) );
A2O1A1Ixp33_ASAP7_75t_SL g1166 ( .A1(n_1167), .A2(n_1182), .B(n_1215), .C(n_1261), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1167), .B(n_1232), .Y(n_1231) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1167), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1303 ( .A(n_1167), .B(n_1304), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1328 ( .A(n_1167), .B(n_1253), .Y(n_1328) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1167), .Y(n_1359) );
AND2x2_ASAP7_75t_L g1364 ( .A(n_1167), .B(n_1199), .Y(n_1364) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1168), .Y(n_1218) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1168), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1168), .B(n_1213), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1168), .B(n_1260), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_1168), .B(n_1199), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1176), .Y(n_1168) );
AND2x6_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1172), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1171), .B(n_1175), .Y(n_1174) );
AND2x4_ASAP7_75t_L g1177 ( .A(n_1171), .B(n_1178), .Y(n_1177) );
AND2x6_ASAP7_75t_L g1180 ( .A(n_1171), .B(n_1181), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1171), .B(n_1175), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1171), .B(n_1175), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1173), .B(n_1179), .Y(n_1178) );
OAI21xp5_ASAP7_75t_L g1424 ( .A1(n_1175), .A2(n_1425), .B(n_1426), .Y(n_1424) );
OAI22xp5_ASAP7_75t_L g1182 ( .A1(n_1183), .A2(n_1198), .B1(n_1205), .B2(n_1214), .Y(n_1182) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
NOR2xp33_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1195), .Y(n_1184) );
NAND2xp5_ASAP7_75t_L g1315 ( .A(n_1185), .B(n_1202), .Y(n_1315) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1227 ( .A(n_1186), .B(n_1224), .Y(n_1227) );
OR2x2_ASAP7_75t_L g1279 ( .A(n_1186), .B(n_1230), .Y(n_1279) );
OR2x2_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1192), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1187), .B(n_1224), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1187), .B(n_1247), .Y(n_1246) );
A2O1A1Ixp33_ASAP7_75t_L g1308 ( .A1(n_1187), .A2(n_1290), .B(n_1309), .C(n_1311), .Y(n_1308) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
OR2x2_ASAP7_75t_L g1196 ( .A(n_1188), .B(n_1197), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1188), .B(n_1192), .Y(n_1239) );
OR2x2_ASAP7_75t_L g1334 ( .A(n_1188), .B(n_1224), .Y(n_1334) );
NOR2xp33_ASAP7_75t_L g1339 ( .A(n_1188), .B(n_1340), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1190), .Y(n_1188) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1192), .Y(n_1197) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1192), .Y(n_1214) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1192), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_1192), .B(n_1230), .Y(n_1299) );
NAND2x1_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1194), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1195), .B(n_1230), .Y(n_1331) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
OR2x2_ASAP7_75t_L g1229 ( .A(n_1196), .B(n_1230), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1198 ( .A(n_1199), .B(n_1202), .Y(n_1198) );
CKINVDCx5p33_ASAP7_75t_R g1213 ( .A(n_1199), .Y(n_1213) );
OR2x2_ASAP7_75t_L g1233 ( .A(n_1199), .B(n_1210), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1199), .B(n_1250), .Y(n_1249) );
OAI22xp5_ASAP7_75t_L g1329 ( .A1(n_1199), .A2(n_1293), .B1(n_1312), .B2(n_1330), .Y(n_1329) );
AND2x4_ASAP7_75t_L g1199 ( .A(n_1200), .B(n_1201), .Y(n_1199) );
INVx3_ASAP7_75t_L g1207 ( .A(n_1202), .Y(n_1207) );
CKINVDCx5p33_ASAP7_75t_R g1222 ( .A(n_1202), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1202), .B(n_1224), .Y(n_1248) );
NAND2xp5_ASAP7_75t_L g1272 ( .A(n_1202), .B(n_1246), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1202), .B(n_1276), .Y(n_1300) );
AND2x4_ASAP7_75t_SL g1202 ( .A(n_1203), .B(n_1204), .Y(n_1202) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
NOR2xp33_ASAP7_75t_L g1206 ( .A(n_1207), .B(n_1208), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1207), .B(n_1230), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1207), .B(n_1209), .Y(n_1260) );
NOR2xp33_ASAP7_75t_L g1318 ( .A(n_1207), .B(n_1319), .Y(n_1318) );
NAND2xp5_ASAP7_75t_L g1326 ( .A(n_1207), .B(n_1239), .Y(n_1326) );
CKINVDCx14_ASAP7_75t_R g1345 ( .A(n_1207), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1207), .B(n_1228), .Y(n_1348) );
AOI211xp5_ASAP7_75t_L g1274 ( .A1(n_1208), .A2(n_1275), .B(n_1277), .C(n_1280), .Y(n_1274) );
OR2x2_ASAP7_75t_L g1208 ( .A(n_1209), .B(n_1213), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1209), .B(n_1270), .Y(n_1269) );
INVx2_ASAP7_75t_L g1319 ( .A(n_1209), .Y(n_1319) );
NOR2xp33_ASAP7_75t_L g1342 ( .A(n_1209), .B(n_1271), .Y(n_1342) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_1209), .B(n_1344), .Y(n_1343) );
INVx2_ASAP7_75t_SL g1209 ( .A(n_1210), .Y(n_1209) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_1210), .B(n_1213), .Y(n_1243) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1210), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1211), .B(n_1212), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1217 ( .A(n_1213), .B(n_1218), .Y(n_1217) );
NAND3xp33_ASAP7_75t_L g1317 ( .A(n_1213), .B(n_1239), .C(n_1318), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1214), .B(n_1230), .Y(n_1322) );
NAND4xp25_ASAP7_75t_SL g1215 ( .A(n_1216), .B(n_1234), .C(n_1251), .D(n_1257), .Y(n_1215) );
AOI22xp5_ASAP7_75t_L g1216 ( .A1(n_1217), .A2(n_1219), .B1(n_1228), .B2(n_1231), .Y(n_1216) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1218), .Y(n_1273) );
OAI211xp5_ASAP7_75t_L g1337 ( .A1(n_1218), .A2(n_1338), .B(n_1341), .C(n_1343), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1220), .B(n_1227), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
OAI21xp5_ASAP7_75t_L g1285 ( .A1(n_1221), .A2(n_1232), .B(n_1286), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1222), .B(n_1223), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1222), .B(n_1242), .Y(n_1241) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1222), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1222), .B(n_1292), .Y(n_1294) );
OR2x2_ASAP7_75t_L g1310 ( .A(n_1222), .B(n_1249), .Y(n_1310) );
NOR2xp33_ASAP7_75t_L g1311 ( .A(n_1222), .B(n_1312), .Y(n_1311) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1224), .Y(n_1230) );
OR2x2_ASAP7_75t_L g1271 ( .A(n_1224), .B(n_1272), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1224), .B(n_1247), .Y(n_1292) );
AOI22xp33_ASAP7_75t_L g1332 ( .A1(n_1224), .A2(n_1333), .B1(n_1335), .B2(n_1336), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1225), .B(n_1226), .Y(n_1224) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1227), .Y(n_1235) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
NOR2xp33_ASAP7_75t_L g1258 ( .A(n_1229), .B(n_1259), .Y(n_1258) );
OR2x2_ASAP7_75t_L g1237 ( .A(n_1230), .B(n_1238), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1302 ( .A(n_1230), .B(n_1246), .Y(n_1302) );
OR2x2_ASAP7_75t_L g1362 ( .A(n_1230), .B(n_1326), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1232), .B(n_1289), .Y(n_1288) );
INVx2_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
O2A1O1Ixp33_ASAP7_75t_L g1234 ( .A1(n_1235), .A2(n_1236), .B(n_1240), .C(n_1244), .Y(n_1234) );
AOI22xp5_ASAP7_75t_L g1338 ( .A1(n_1235), .A2(n_1243), .B1(n_1319), .B2(n_1339), .Y(n_1338) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
AOI21xp5_ASAP7_75t_L g1244 ( .A1(n_1237), .A2(n_1245), .B(n_1249), .Y(n_1244) );
OR2x2_ASAP7_75t_L g1255 ( .A(n_1238), .B(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1239), .B(n_1248), .Y(n_1270) );
OAI211xp5_ASAP7_75t_L g1297 ( .A1(n_1239), .A2(n_1242), .B(n_1298), .C(n_1300), .Y(n_1297) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1242), .Y(n_1312) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
OR2x2_ASAP7_75t_L g1358 ( .A(n_1243), .B(n_1359), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1246), .B(n_1248), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_1246), .B(n_1351), .Y(n_1350) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1248), .Y(n_1340) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1249), .Y(n_1284) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1249), .Y(n_1304) );
INVx2_ASAP7_75t_L g1253 ( .A(n_1250), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1252), .B(n_1254), .Y(n_1251) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
OR2x2_ASAP7_75t_L g1275 ( .A(n_1253), .B(n_1276), .Y(n_1275) );
AOI21xp5_ASAP7_75t_L g1349 ( .A1(n_1253), .A2(n_1350), .B(n_1352), .Y(n_1349) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
A2O1A1Ixp33_ASAP7_75t_L g1281 ( .A1(n_1255), .A2(n_1282), .B(n_1283), .C(n_1285), .Y(n_1281) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1256), .Y(n_1351) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
CKINVDCx14_ASAP7_75t_R g1280 ( .A(n_1261), .Y(n_1280) );
A2O1A1Ixp33_ASAP7_75t_L g1346 ( .A1(n_1261), .A2(n_1347), .B(n_1349), .C(n_1354), .Y(n_1346) );
INVx3_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
OAI221xp5_ASAP7_75t_L g1320 ( .A1(n_1262), .A2(n_1291), .B1(n_1295), .B2(n_1321), .C(n_1323), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1263), .B(n_1265), .Y(n_1262) );
HB1xp67_ASAP7_75t_L g1368 ( .A(n_1264), .Y(n_1368) );
NOR5xp2_ASAP7_75t_L g1266 ( .A(n_1267), .B(n_1274), .C(n_1281), .D(n_1287), .E(n_1301), .Y(n_1266) );
AOI21xp33_ASAP7_75t_L g1267 ( .A1(n_1268), .A2(n_1271), .B(n_1273), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
INVxp67_ASAP7_75t_L g1282 ( .A(n_1270), .Y(n_1282) );
OR2x2_ASAP7_75t_L g1277 ( .A(n_1278), .B(n_1279), .Y(n_1277) );
INVx2_ASAP7_75t_L g1286 ( .A(n_1279), .Y(n_1286) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
AOI211xp5_ASAP7_75t_L g1313 ( .A1(n_1284), .A2(n_1314), .B(n_1316), .C(n_1320), .Y(n_1313) );
NAND2xp5_ASAP7_75t_L g1353 ( .A(n_1286), .B(n_1345), .Y(n_1353) );
OAI221xp5_ASAP7_75t_SL g1287 ( .A1(n_1288), .A2(n_1291), .B1(n_1293), .B2(n_1295), .C(n_1297), .Y(n_1287) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1288), .Y(n_1336) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
NOR2xp33_ASAP7_75t_L g1301 ( .A(n_1302), .B(n_1303), .Y(n_1301) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1302), .Y(n_1327) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1303), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1306), .B(n_1356), .Y(n_1305) );
OAI21xp5_ASAP7_75t_L g1306 ( .A1(n_1307), .A2(n_1337), .B(n_1346), .Y(n_1306) );
NAND4xp25_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1313), .C(n_1324), .D(n_1332), .Y(n_1307) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
OAI21xp5_ASAP7_75t_SL g1357 ( .A1(n_1321), .A2(n_1358), .B(n_1360), .Y(n_1357) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
O2A1O1Ixp33_ASAP7_75t_L g1324 ( .A1(n_1325), .A2(n_1327), .B(n_1328), .C(n_1329), .Y(n_1324) );
AOI22xp5_ASAP7_75t_L g1356 ( .A1(n_1325), .A2(n_1345), .B1(n_1357), .B2(n_1365), .Y(n_1356) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
INVx2_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1331), .B(n_1345), .Y(n_1344) );
OAI31xp33_ASAP7_75t_L g1360 ( .A1(n_1333), .A2(n_1361), .A3(n_1363), .B(n_1364), .Y(n_1360) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
A2O1A1Ixp33_ASAP7_75t_L g1365 ( .A1(n_1334), .A2(n_1358), .B(n_1362), .C(n_1366), .Y(n_1365) );
INVxp67_ASAP7_75t_SL g1341 ( .A(n_1342), .Y(n_1341) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1358), .Y(n_1363) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1364), .Y(n_1366) );
INVx4_ASAP7_75t_L g1367 ( .A(n_1368), .Y(n_1367) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
HB1xp67_ASAP7_75t_L g1423 ( .A(n_1373), .Y(n_1423) );
NAND3xp33_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1401), .C(n_1408), .Y(n_1373) );
NOR2xp33_ASAP7_75t_L g1374 ( .A(n_1375), .B(n_1393), .Y(n_1374) );
OAI33xp33_ASAP7_75t_L g1375 ( .A1(n_1376), .A2(n_1380), .A3(n_1383), .B1(n_1385), .B2(n_1388), .B3(n_1389), .Y(n_1375) );
OAI22xp5_ASAP7_75t_L g1397 ( .A1(n_1382), .A2(n_1387), .B1(n_1398), .B2(n_1399), .Y(n_1397) );
BUFx3_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
INVx2_ASAP7_75t_L g1414 ( .A(n_1415), .Y(n_1414) );
BUFx3_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
BUFx3_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
INVxp33_ASAP7_75t_L g1421 ( .A(n_1422), .Y(n_1421) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
endmodule