module fake_jpeg_11525_n_435 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_435);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_435;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_14),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_55),
.B(n_97),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_56),
.Y(n_151)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_57),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_58),
.B(n_62),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_22),
.B(n_11),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_61),
.B(n_85),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_22),
.B(n_11),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_65),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_66),
.Y(n_164)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_70),
.Y(n_160)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_71),
.Y(n_168)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_23),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_78),
.Y(n_119)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_75),
.Y(n_115)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_23),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_81),
.Y(n_171)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_83),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_26),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_84),
.B(n_88),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_26),
.B(n_9),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_32),
.B(n_0),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_32),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_93),
.Y(n_140)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_91),
.Y(n_183)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_92),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_41),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_95),
.Y(n_170)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_96),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_41),
.B(n_43),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_98),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_43),
.B(n_0),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_104),
.Y(n_143)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_100),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

BUFx10_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_102),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_34),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_20),
.Y(n_105)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_106),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_51),
.B(n_50),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_112),
.Y(n_154)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_36),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_L g158 ( 
.A1(n_108),
.A2(n_111),
.B(n_2),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_109),
.B(n_110),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

INVx6_ASAP7_75t_SL g112 ( 
.A(n_34),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_35),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_113),
.B(n_35),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_30),
.B1(n_45),
.B2(n_31),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g204 ( 
.A1(n_122),
.A2(n_130),
.B1(n_151),
.B2(n_162),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_110),
.A2(n_45),
.B1(n_51),
.B2(n_31),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_127),
.A2(n_136),
.B1(n_152),
.B2(n_163),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_69),
.A2(n_31),
.B1(n_35),
.B2(n_45),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_130),
.A2(n_153),
.B1(n_159),
.B2(n_162),
.Y(n_188)
);

AO22x1_ASAP7_75t_SL g131 ( 
.A1(n_72),
.A2(n_54),
.B1(n_52),
.B2(n_39),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_131),
.B(n_175),
.Y(n_208)
);

OR2x4_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_20),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_132),
.B(n_122),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_71),
.A2(n_27),
.B1(n_46),
.B2(n_42),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_133),
.A2(n_144),
.B1(n_172),
.B2(n_175),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_73),
.A2(n_27),
.B1(n_46),
.B2(n_42),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_137),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_56),
.A2(n_17),
.B1(n_37),
.B2(n_28),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_76),
.A2(n_54),
.B1(n_52),
.B2(n_39),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_145),
.A2(n_157),
.B(n_115),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_59),
.A2(n_37),
.B1(n_28),
.B2(n_24),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_67),
.A2(n_24),
.B1(n_17),
.B2(n_4),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_64),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_156),
.A2(n_159),
.B(n_131),
.C(n_153),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_77),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_158),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_66),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_66),
.A2(n_91),
.B1(n_108),
.B2(n_106),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_65),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_111),
.A2(n_8),
.B1(n_95),
.B2(n_105),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_165),
.A2(n_174),
.B1(n_115),
.B2(n_114),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_80),
.A2(n_103),
.B1(n_102),
.B2(n_94),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_82),
.A2(n_87),
.B1(n_98),
.B2(n_79),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_92),
.A2(n_113),
.B1(n_79),
.B2(n_101),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_68),
.B(n_70),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_179),
.B(n_132),
.Y(n_201)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_185),
.Y(n_250)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_186),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_128),
.B(n_75),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_187),
.B(n_189),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_119),
.B(n_75),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_190),
.Y(n_249)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_191),
.Y(n_254)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_126),
.Y(n_192)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_192),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_193),
.B(n_208),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_140),
.B(n_161),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_194),
.B(n_202),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_125),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_195),
.B(n_203),
.Y(n_247)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_196),
.Y(n_275)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_197),
.Y(n_256)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_198),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_200),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_201),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_118),
.B(n_139),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_143),
.B(n_154),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_204),
.A2(n_228),
.B1(n_227),
.B2(n_220),
.Y(n_284)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_205),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_148),
.B(n_149),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_206),
.B(n_214),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_137),
.A2(n_156),
.B(n_131),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_207),
.A2(n_184),
.B(n_204),
.Y(n_269)
);

NOR2x1_ASAP7_75t_R g264 ( 
.A(n_209),
.B(n_221),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_150),
.B(n_166),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_210),
.B(n_231),
.Y(n_262)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_211),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_151),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_213),
.A2(n_229),
.B1(n_234),
.B2(n_235),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_177),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_215),
.Y(n_255)
);

O2A1O1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_129),
.A2(n_141),
.B(n_180),
.C(n_160),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_216),
.A2(n_208),
.B(n_221),
.C(n_243),
.Y(n_258)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

INVx13_ASAP7_75t_L g260 ( 
.A(n_217),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

CKINVDCx10_ASAP7_75t_R g253 ( 
.A(n_218),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_171),
.B(n_173),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_219),
.B(n_223),
.Y(n_266)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_147),
.Y(n_220)
);

INVx13_ASAP7_75t_L g267 ( 
.A(n_220),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_129),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_142),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_225),
.B(n_226),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_114),
.B(n_164),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_147),
.Y(n_227)
);

INVx13_ASAP7_75t_L g280 ( 
.A(n_227),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_114),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_228),
.B(n_230),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_116),
.B(n_120),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_121),
.B(n_138),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_120),
.B(n_155),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_232),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_129),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_233),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_123),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_155),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_135),
.B(n_174),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_236),
.B(n_237),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_141),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_141),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_238),
.B(n_241),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_165),
.B(n_124),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_239),
.A2(n_240),
.B1(n_193),
.B2(n_188),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_124),
.A2(n_134),
.B1(n_123),
.B2(n_167),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_135),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_168),
.B(n_134),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_242),
.B(n_243),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_168),
.B(n_167),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_146),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_222),
.C(n_231),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_246),
.B(n_218),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_248),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g252 ( 
.A(n_224),
.B(n_207),
.CI(n_210),
.CON(n_252),
.SN(n_252)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_252),
.B(n_199),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_258),
.B(n_253),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_184),
.A2(n_224),
.B1(n_212),
.B2(n_209),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_268),
.A2(n_286),
.B1(n_185),
.B2(n_186),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_269),
.A2(n_238),
.B(n_211),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_200),
.B(n_192),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_274),
.B(n_279),
.C(n_283),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_190),
.B(n_196),
.C(n_235),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_216),
.B(n_241),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_284),
.A2(n_257),
.B1(n_285),
.B2(n_259),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_198),
.A2(n_213),
.B1(n_234),
.B2(n_205),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_290),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_291),
.B(n_310),
.Y(n_337)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_292),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_293),
.A2(n_317),
.B(n_316),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_273),
.A2(n_217),
.B(n_197),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_295),
.A2(n_302),
.B(n_317),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_296),
.A2(n_298),
.B1(n_312),
.B2(n_314),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_297),
.B(n_306),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_273),
.A2(n_218),
.B1(n_269),
.B2(n_262),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_299),
.A2(n_300),
.B1(n_318),
.B2(n_319),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_262),
.B1(n_288),
.B2(n_273),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_259),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_301),
.B(n_303),
.Y(n_335)
);

NAND3xp33_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_265),
.C(n_266),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_278),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_256),
.Y(n_304)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_304),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_287),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_305),
.B(n_315),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_288),
.B(n_276),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_309),
.Y(n_330)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_308),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_274),
.B(n_251),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_277),
.B(n_247),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_246),
.B(n_289),
.C(n_252),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_311),
.B(n_260),
.C(n_307),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_258),
.A2(n_286),
.B1(n_283),
.B2(n_285),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_263),
.Y(n_313)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_313),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_264),
.A2(n_252),
.B1(n_279),
.B2(n_287),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_272),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_264),
.B(n_255),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_316),
.B(n_323),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_254),
.A2(n_249),
.B1(n_275),
.B2(n_281),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_281),
.A2(n_249),
.B1(n_275),
.B2(n_263),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_282),
.A2(n_256),
.B1(n_261),
.B2(n_250),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_320),
.B(n_324),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_282),
.B(n_250),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_321),
.B(n_322),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_261),
.B(n_253),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_245),
.B(n_267),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_245),
.B(n_267),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_298),
.A2(n_260),
.B1(n_280),
.B2(n_314),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_325),
.A2(n_349),
.B1(n_294),
.B2(n_299),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_280),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_326),
.B(n_331),
.C(n_348),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_318),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_301),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_332),
.C(n_348),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_306),
.C(n_297),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_295),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_313),
.Y(n_368)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_290),
.Y(n_342)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_342),
.Y(n_352)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_292),
.Y(n_345)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_345),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_346),
.B(n_321),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_317),
.B(n_300),
.C(n_305),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_296),
.A2(n_294),
.B1(n_291),
.B2(n_293),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_351),
.A2(n_355),
.B(n_364),
.Y(n_383)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_353),
.Y(n_375)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_327),
.Y(n_357)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_357),
.Y(n_382)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_327),
.Y(n_358)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_358),
.Y(n_384)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_329),
.Y(n_359)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_359),
.Y(n_386)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_329),
.Y(n_360)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_360),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_337),
.B(n_310),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_361),
.B(n_365),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_333),
.A2(n_315),
.B1(n_302),
.B2(n_324),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_362),
.A2(n_344),
.B1(n_346),
.B2(n_343),
.Y(n_374)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_342),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_363),
.B(n_366),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_349),
.A2(n_322),
.B1(n_323),
.B2(n_320),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_337),
.B(n_335),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_325),
.A2(n_304),
.B1(n_319),
.B2(n_308),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_367),
.B(n_371),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_368),
.B(n_369),
.C(n_326),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_339),
.B(n_332),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_347),
.B(n_330),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_370),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_373),
.B(n_380),
.C(n_371),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_350),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_369),
.B(n_330),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_379),
.B(n_381),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_354),
.B(n_344),
.C(n_343),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_354),
.B(n_336),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_362),
.B(n_347),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_387),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_375),
.Y(n_390)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_390),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_391),
.B(n_397),
.Y(n_403)
);

A2O1A1O1Ixp25_ASAP7_75t_L g392 ( 
.A1(n_387),
.A2(n_355),
.B(n_335),
.C(n_340),
.D(n_351),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_392),
.B(n_396),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_368),
.C(n_340),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_393),
.B(n_394),
.C(n_395),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_377),
.B(n_364),
.C(n_333),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_380),
.B(n_356),
.C(n_357),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_372),
.A2(n_366),
.B(n_352),
.Y(n_396)
);

XOR2x1_ASAP7_75t_SL g397 ( 
.A(n_374),
.B(n_350),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_398),
.A2(n_378),
.B(n_383),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_373),
.B(n_352),
.C(n_360),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_399),
.B(n_379),
.C(n_381),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_385),
.B(n_334),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_400),
.B(n_385),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_404),
.B(n_407),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_398),
.A2(n_383),
.B(n_378),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_406),
.A2(n_392),
.B(n_376),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_389),
.A2(n_328),
.B1(n_376),
.B2(n_386),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_408),
.B(n_356),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_409),
.B(n_410),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_391),
.B(n_384),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_410),
.B(n_393),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_412),
.B(n_413),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_402),
.B(n_382),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_409),
.B(n_388),
.C(n_394),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_416),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_405),
.B(n_388),
.C(n_397),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_417),
.A2(n_401),
.B(n_404),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_418),
.A2(n_406),
.B1(n_402),
.B2(n_359),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_419),
.B(n_420),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_411),
.A2(n_401),
.B(n_403),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_415),
.A2(n_405),
.B(n_407),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_421),
.B(n_414),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_422),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_425),
.B(n_428),
.C(n_423),
.Y(n_429)
);

MAJx2_ASAP7_75t_L g428 ( 
.A(n_424),
.B(n_416),
.C(n_403),
.Y(n_428)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_429),
.Y(n_431)
);

AOI322xp5_ASAP7_75t_L g430 ( 
.A1(n_427),
.A2(n_426),
.A3(n_423),
.B1(n_408),
.B2(n_358),
.C1(n_363),
.C2(n_345),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_430),
.B(n_338),
.C(n_341),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_432),
.B(n_338),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_433),
.B(n_431),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_434),
.B(n_334),
.Y(n_435)
);


endmodule