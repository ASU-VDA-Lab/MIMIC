module fake_jpeg_18910_n_154 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_154);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_15),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_0),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_26),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_4),
.Y(n_71)
);

BUFx4f_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_6),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_78),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_77),
.Y(n_86)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_1),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_78),
.A2(n_48),
.B1(n_71),
.B2(n_72),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_84),
.B(n_59),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_54),
.B1(n_55),
.B2(n_62),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_53),
.C(n_54),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_92),
.A2(n_59),
.B1(n_70),
.B2(n_65),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_53),
.C(n_58),
.Y(n_118)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_97),
.Y(n_109)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_67),
.B1(n_66),
.B2(n_63),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_51),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_99),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_56),
.B1(n_49),
.B2(n_61),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_101),
.A2(n_8),
.B(n_9),
.C(n_13),
.Y(n_123)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_103),
.Y(n_115)
);

INVx6_ASAP7_75t_SL g103 ( 
.A(n_83),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_104),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_SL g110 ( 
.A(n_105),
.B(n_46),
.C(n_49),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_69),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_1),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_110),
.B(n_116),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_114),
.B1(n_120),
.B2(n_8),
.Y(n_124)
);

FAx1_ASAP7_75t_SL g113 ( 
.A(n_102),
.B(n_61),
.CI(n_2),
.CON(n_113),
.SN(n_113)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_113),
.B(n_121),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_50),
.B1(n_3),
.B2(n_5),
.Y(n_114)
);

AND2x6_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_56),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_118),
.A2(n_123),
.B1(n_19),
.B2(n_21),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_96),
.B(n_25),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_23),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_101),
.B1(n_5),
.B2(n_7),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_7),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_122),
.A2(n_14),
.B(n_17),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_124),
.A2(n_108),
.B1(n_132),
.B2(n_112),
.Y(n_140)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_132),
.Y(n_141)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_130),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_119),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_131),
.B(n_127),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_133),
.A2(n_134),
.B(n_135),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_28),
.Y(n_135)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_140),
.A2(n_141),
.B1(n_139),
.B2(n_123),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_136),
.C(n_137),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_142),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_138),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_146),
.A2(n_112),
.B1(n_130),
.B2(n_128),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_33),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_35),
.B(n_36),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g151 ( 
.A(n_150),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_37),
.B(n_39),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_42),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_43),
.Y(n_154)
);


endmodule