module fake_jpeg_20047_n_46 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_46);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_46;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_32;
wire n_15;

INVxp67_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_17),
.A2(n_5),
.B(n_29),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_32),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_28),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_37),
.B1(n_31),
.B2(n_36),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_38),
.B(n_14),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_39),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_18),
.C(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_44),
.B(n_43),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_21),
.Y(n_46)
);


endmodule