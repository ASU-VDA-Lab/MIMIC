module fake_aes_8590_n_739 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_739);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_739;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_23), .Y(n_82) );
INVxp33_ASAP7_75t_L g83 ( .A(n_48), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_79), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_73), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_8), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_5), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_28), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_46), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_62), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_71), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_20), .Y(n_92) );
CKINVDCx16_ASAP7_75t_R g93 ( .A(n_4), .Y(n_93) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_30), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_42), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_27), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_66), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_74), .Y(n_98) );
BUFx3_ASAP7_75t_L g99 ( .A(n_14), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_33), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_5), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_59), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_45), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_63), .Y(n_104) );
INVxp33_ASAP7_75t_SL g105 ( .A(n_17), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_67), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_15), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_55), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_80), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_34), .B(n_7), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_19), .Y(n_111) );
INVxp33_ASAP7_75t_L g112 ( .A(n_38), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_72), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_22), .Y(n_114) );
BUFx2_ASAP7_75t_SL g115 ( .A(n_49), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_16), .Y(n_116) );
CKINVDCx14_ASAP7_75t_R g117 ( .A(n_68), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_61), .Y(n_118) );
BUFx3_ASAP7_75t_L g119 ( .A(n_54), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_35), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_57), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_39), .Y(n_122) );
INVxp67_ASAP7_75t_L g123 ( .A(n_3), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_0), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_29), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_16), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_1), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_1), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_51), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_52), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_81), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_94), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_93), .B(n_0), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_85), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_84), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_88), .Y(n_137) );
CKINVDCx11_ASAP7_75t_R g138 ( .A(n_99), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_84), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_123), .B(n_2), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_94), .B(n_2), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_88), .Y(n_142) );
INVx4_ASAP7_75t_L g143 ( .A(n_119), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_89), .Y(n_144) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_105), .A2(n_3), .B1(n_4), .B2(n_6), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_89), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_90), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_94), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_90), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_91), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_91), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_99), .B(n_6), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_95), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_128), .Y(n_154) );
BUFx2_ASAP7_75t_L g155 ( .A(n_86), .Y(n_155) );
INVxp67_ASAP7_75t_L g156 ( .A(n_111), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_95), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_96), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g159 ( .A1(n_87), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_127), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_83), .B(n_9), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_128), .B(n_10), .Y(n_162) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_87), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_96), .Y(n_164) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_101), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_112), .B(n_10), .Y(n_166) );
BUFx8_ASAP7_75t_L g167 ( .A(n_94), .Y(n_167) );
BUFx2_ASAP7_75t_L g168 ( .A(n_117), .Y(n_168) );
OAI22xp33_ASAP7_75t_L g169 ( .A1(n_101), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_97), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_94), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_97), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_98), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_98), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_116), .B(n_11), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_109), .B(n_12), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_100), .Y(n_177) );
INVx4_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_152), .B(n_114), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_168), .B(n_121), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_172), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_160), .Y(n_182) );
BUFx2_ASAP7_75t_L g183 ( .A(n_168), .Y(n_183) );
OR2x6_ASAP7_75t_L g184 ( .A(n_159), .B(n_115), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_155), .B(n_82), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_172), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_132), .Y(n_187) );
INVxp67_ASAP7_75t_L g188 ( .A(n_155), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_132), .Y(n_189) );
AND2x4_ASAP7_75t_L g190 ( .A(n_152), .B(n_114), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_167), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_172), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_132), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_156), .B(n_106), .Y(n_194) );
NAND3xp33_ASAP7_75t_L g195 ( .A(n_163), .B(n_107), .C(n_124), .Y(n_195) );
OAI221xp5_ASAP7_75t_L g196 ( .A1(n_165), .A2(n_107), .B1(n_126), .B2(n_124), .C(n_92), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_162), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_162), .Y(n_198) );
INVx6_ASAP7_75t_L g199 ( .A(n_167), .Y(n_199) );
OA22x2_ASAP7_75t_L g200 ( .A1(n_145), .A2(n_126), .B1(n_131), .B2(n_129), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_132), .Y(n_201) );
INVx4_ASAP7_75t_L g202 ( .A(n_152), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_132), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_134), .B(n_113), .Y(n_204) );
INVx4_ASAP7_75t_L g205 ( .A(n_143), .Y(n_205) );
INVx1_ASAP7_75t_SL g206 ( .A(n_138), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_132), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_148), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_162), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_148), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_172), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_162), .B(n_131), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_134), .B(n_135), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_177), .B(n_130), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_148), .Y(n_215) );
BUFx3_ASAP7_75t_L g216 ( .A(n_167), .Y(n_216) );
INVx4_ASAP7_75t_L g217 ( .A(n_143), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_177), .B(n_130), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_135), .B(n_129), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_148), .Y(n_220) );
INVxp33_ASAP7_75t_L g221 ( .A(n_161), .Y(n_221) );
NAND2x1p5_ASAP7_75t_L g222 ( .A(n_137), .B(n_125), .Y(n_222) );
INVx2_ASAP7_75t_SL g223 ( .A(n_167), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_148), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_137), .B(n_120), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_144), .B(n_125), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_161), .B(n_119), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_144), .B(n_122), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_136), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_142), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_146), .B(n_122), .Y(n_231) );
NOR2xp33_ASAP7_75t_SL g232 ( .A(n_166), .B(n_118), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_142), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_151), .Y(n_234) );
OR2x6_ASAP7_75t_L g235 ( .A(n_133), .B(n_115), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_146), .B(n_108), .Y(n_236) );
INVx2_ASAP7_75t_SL g237 ( .A(n_166), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_147), .B(n_108), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_147), .B(n_103), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_149), .B(n_103), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_151), .Y(n_241) );
NAND2x1p5_ASAP7_75t_L g242 ( .A(n_149), .B(n_102), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_148), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_171), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_171), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_181), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_221), .B(n_150), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_181), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_222), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_186), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_222), .Y(n_251) );
INVx5_ASAP7_75t_L g252 ( .A(n_199), .Y(n_252) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_199), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_222), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_237), .B(n_145), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_242), .Y(n_256) );
INVx3_ASAP7_75t_L g257 ( .A(n_178), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_186), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_227), .B(n_153), .Y(n_259) );
BUFx12f_ASAP7_75t_L g260 ( .A(n_183), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_237), .B(n_140), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_191), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_242), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_227), .B(n_170), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_182), .Y(n_265) );
NOR2x1_ASAP7_75t_R g266 ( .A(n_182), .B(n_104), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_242), .B(n_153), .Y(n_267) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_199), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_192), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_206), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_229), .Y(n_271) );
OAI22xp5_ASAP7_75t_SL g272 ( .A1(n_184), .A2(n_169), .B1(n_175), .B2(n_176), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_191), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_199), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_235), .B(n_174), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_214), .B(n_174), .Y(n_276) );
INVx3_ASAP7_75t_L g277 ( .A(n_178), .Y(n_277) );
INVxp67_ASAP7_75t_SL g278 ( .A(n_216), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_229), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_192), .Y(n_280) );
INVx2_ASAP7_75t_SL g281 ( .A(n_216), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_211), .Y(n_282) );
BUFx12f_ASAP7_75t_L g283 ( .A(n_183), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_235), .B(n_173), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_198), .Y(n_285) );
BUFx2_ASAP7_75t_L g286 ( .A(n_188), .Y(n_286) );
OR2x6_ASAP7_75t_L g287 ( .A(n_235), .B(n_173), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_235), .B(n_158), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_185), .B(n_150), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_200), .A2(n_157), .B1(n_170), .B2(n_164), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_221), .B(n_158), .Y(n_291) );
INVx2_ASAP7_75t_SL g292 ( .A(n_178), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_198), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_214), .B(n_164), .Y(n_294) );
BUFx2_ASAP7_75t_L g295 ( .A(n_202), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_202), .B(n_157), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_198), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_202), .Y(n_298) );
AND2x6_ASAP7_75t_SL g299 ( .A(n_184), .B(n_110), .Y(n_299) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_223), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_223), .Y(n_301) );
OR2x6_ASAP7_75t_L g302 ( .A(n_184), .B(n_141), .Y(n_302) );
BUFx4f_ASAP7_75t_L g303 ( .A(n_179), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_211), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_214), .B(n_143), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_209), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_209), .Y(n_307) );
AO22x1_ASAP7_75t_L g308 ( .A1(n_179), .A2(n_100), .B1(n_102), .B2(n_154), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_209), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_179), .Y(n_310) );
BUFx12f_ASAP7_75t_SL g311 ( .A(n_184), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_218), .B(n_143), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_218), .Y(n_313) );
INVx5_ASAP7_75t_L g314 ( .A(n_205), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_218), .B(n_154), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_219), .Y(n_316) );
INVx4_ASAP7_75t_L g317 ( .A(n_190), .Y(n_317) );
CKINVDCx6p67_ASAP7_75t_R g318 ( .A(n_190), .Y(n_318) );
INVx4_ASAP7_75t_L g319 ( .A(n_318), .Y(n_319) );
HAxp5_ASAP7_75t_L g320 ( .A(n_255), .B(n_200), .CON(n_320), .SN(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_287), .B(n_190), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_247), .B(n_291), .Y(n_322) );
AOI21x1_ASAP7_75t_L g323 ( .A1(n_308), .A2(n_197), .B(n_228), .Y(n_323) );
O2A1O1Ixp33_ASAP7_75t_L g324 ( .A1(n_259), .A2(n_196), .B(n_236), .C(n_240), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_287), .B(n_212), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_247), .B(n_232), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_313), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_246), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_291), .B(n_289), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_285), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_253), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_318), .A2(n_212), .B1(n_226), .B2(n_238), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_286), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g334 ( .A1(n_316), .A2(n_200), .B1(n_212), .B2(n_226), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_287), .B(n_219), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_313), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_313), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_293), .Y(n_338) );
INVx2_ASAP7_75t_SL g339 ( .A(n_303), .Y(n_339) );
AND2x2_ASAP7_75t_SL g340 ( .A(n_249), .B(n_219), .Y(n_340) );
BUFx2_ASAP7_75t_R g341 ( .A(n_270), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_286), .B(n_239), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_246), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_248), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_253), .Y(n_345) );
A2O1A1Ixp33_ASAP7_75t_L g346 ( .A1(n_276), .A2(n_213), .B(n_195), .C(n_238), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_248), .Y(n_347) );
AO21x1_ASAP7_75t_L g348 ( .A1(n_267), .A2(n_226), .B(n_238), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_255), .B(n_180), .Y(n_349) );
AO21x2_ASAP7_75t_L g350 ( .A1(n_267), .A2(n_231), .B(n_225), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_297), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_306), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_255), .A2(n_239), .B1(n_241), .B2(n_233), .Y(n_353) );
INVx2_ASAP7_75t_SL g354 ( .A(n_303), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_307), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_309), .Y(n_356) );
AND3x2_ASAP7_75t_L g357 ( .A(n_270), .B(n_136), .C(n_139), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_296), .A2(n_205), .B(n_217), .Y(n_358) );
AOI222xp33_ASAP7_75t_L g359 ( .A1(n_272), .A2(n_194), .B1(n_154), .B2(n_234), .C1(n_230), .C2(n_204), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_250), .Y(n_360) );
BUFx12f_ASAP7_75t_L g361 ( .A(n_260), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_250), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_258), .Y(n_363) );
BUFx2_ASAP7_75t_L g364 ( .A(n_260), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_258), .Y(n_365) );
CKINVDCx11_ASAP7_75t_R g366 ( .A(n_283), .Y(n_366) );
AND2x2_ASAP7_75t_SL g367 ( .A(n_251), .B(n_205), .Y(n_367) );
INVx1_ASAP7_75t_SL g368 ( .A(n_283), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_254), .A2(n_263), .B1(n_256), .B2(n_303), .Y(n_369) );
INVx2_ASAP7_75t_SL g370 ( .A(n_262), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_269), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_261), .B(n_217), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_313), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_269), .Y(n_374) );
NAND2x1p5_ASAP7_75t_L g375 ( .A(n_317), .B(n_217), .Y(n_375) );
INVxp67_ASAP7_75t_L g376 ( .A(n_333), .Y(n_376) );
INVx3_ASAP7_75t_L g377 ( .A(n_327), .Y(n_377) );
BUFx2_ASAP7_75t_L g378 ( .A(n_335), .Y(n_378) );
AOI22xp33_ASAP7_75t_SL g379 ( .A1(n_340), .A2(n_265), .B1(n_361), .B2(n_364), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_360), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_353), .B(n_290), .Y(n_381) );
BUFx3_ASAP7_75t_L g382 ( .A(n_335), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_349), .A2(n_261), .B1(n_265), .B2(n_264), .C(n_294), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_360), .Y(n_384) );
NAND3xp33_ASAP7_75t_L g385 ( .A(n_359), .B(n_302), .C(n_287), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_340), .A2(n_311), .B1(n_284), .B2(n_288), .Y(n_386) );
AO31x2_ASAP7_75t_L g387 ( .A1(n_348), .A2(n_139), .A3(n_271), .B(n_279), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_340), .A2(n_311), .B1(n_275), .B2(n_288), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_335), .Y(n_389) );
AOI21xp5_ASAP7_75t_SL g390 ( .A1(n_332), .A2(n_275), .B(n_288), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_366), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_321), .B(n_262), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_361), .Y(n_393) );
OAI22xp33_ASAP7_75t_L g394 ( .A1(n_329), .A2(n_317), .B1(n_302), .B2(n_313), .Y(n_394) );
AND2x6_ASAP7_75t_L g395 ( .A(n_325), .B(n_321), .Y(n_395) );
BUFx3_ASAP7_75t_L g396 ( .A(n_325), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_341), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_342), .A2(n_284), .B1(n_275), .B2(n_317), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_364), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_363), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_328), .Y(n_401) );
INVx2_ASAP7_75t_SL g402 ( .A(n_325), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_363), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_328), .Y(n_404) );
INVx3_ASAP7_75t_L g405 ( .A(n_327), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_374), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_367), .A2(n_284), .B1(n_302), .B2(n_310), .Y(n_407) );
AOI211xp5_ASAP7_75t_L g408 ( .A1(n_342), .A2(n_266), .B(n_261), .C(n_315), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_343), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_343), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_374), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g412 ( .A1(n_390), .A2(n_369), .B(n_367), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_380), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_380), .Y(n_414) );
OAI21xp5_ASAP7_75t_SL g415 ( .A1(n_379), .A2(n_357), .B(n_334), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_383), .A2(n_322), .B1(n_324), .B2(n_326), .C(n_346), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_385), .A2(n_302), .B1(n_321), .B2(n_367), .Y(n_417) );
BUFx2_ASAP7_75t_L g418 ( .A(n_395), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_384), .Y(n_419) );
OAI22xp5_ASAP7_75t_SL g420 ( .A1(n_408), .A2(n_368), .B1(n_334), .B2(n_319), .Y(n_420) );
OAI221xp5_ASAP7_75t_L g421 ( .A1(n_408), .A2(n_339), .B1(n_354), .B2(n_372), .C(n_319), .Y(n_421) );
HB1xp67_ASAP7_75t_SL g422 ( .A(n_393), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_385), .A2(n_348), .B1(n_319), .B2(n_354), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_407), .A2(n_339), .B1(n_330), .B2(n_338), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_407), .A2(n_351), .B1(n_330), .B2(n_338), .Y(n_425) );
INVx5_ASAP7_75t_SL g426 ( .A(n_395), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_376), .A2(n_352), .B1(n_351), .B2(n_355), .C(n_356), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_394), .A2(n_355), .B1(n_352), .B2(n_356), .Y(n_428) );
AOI222xp33_ASAP7_75t_L g429 ( .A1(n_381), .A2(n_320), .B1(n_154), .B2(n_344), .C1(n_371), .C2(n_347), .Y(n_429) );
AOI221x1_ASAP7_75t_SL g430 ( .A1(n_381), .A2(n_320), .B1(n_299), .B2(n_15), .C(n_17), .Y(n_430) );
AO21x2_ASAP7_75t_L g431 ( .A1(n_384), .A2(n_323), .B(n_350), .Y(n_431) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_400), .A2(n_323), .B(n_358), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_395), .A2(n_350), .B1(n_373), .B2(n_336), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_400), .B(n_344), .Y(n_434) );
OAI211xp5_ASAP7_75t_L g435 ( .A1(n_390), .A2(n_312), .B(n_305), .C(n_296), .Y(n_435) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_395), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_395), .B(n_347), .Y(n_437) );
OA21x2_ASAP7_75t_L g438 ( .A1(n_403), .A2(n_371), .B(n_365), .Y(n_438) );
AOI22xp33_ASAP7_75t_SL g439 ( .A1(n_395), .A2(n_278), .B1(n_370), .B2(n_362), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_403), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_401), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_420), .A2(n_395), .B1(n_378), .B2(n_389), .Y(n_442) );
OA21x2_ASAP7_75t_L g443 ( .A1(n_432), .A2(n_411), .B(n_406), .Y(n_443) );
NAND3xp33_ASAP7_75t_L g444 ( .A(n_416), .B(n_411), .C(n_406), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_438), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_420), .A2(n_395), .B1(n_378), .B2(n_382), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_438), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_413), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_430), .B(n_398), .Y(n_449) );
AOI221xp5_ASAP7_75t_L g450 ( .A1(n_430), .A2(n_386), .B1(n_388), .B2(n_399), .C(n_397), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_415), .B(n_391), .Y(n_451) );
AOI22xp33_ASAP7_75t_SL g452 ( .A1(n_426), .A2(n_418), .B1(n_412), .B2(n_436), .Y(n_452) );
AOI33xp33_ASAP7_75t_L g453 ( .A1(n_425), .A2(n_402), .A3(n_410), .B1(n_404), .B2(n_409), .B3(n_401), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_413), .B(n_402), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_414), .B(n_387), .Y(n_455) );
OAI21xp5_ASAP7_75t_SL g456 ( .A1(n_415), .A2(n_392), .B(n_375), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_434), .Y(n_457) );
AOI221xp5_ASAP7_75t_L g458 ( .A1(n_427), .A2(n_382), .B1(n_389), .B2(n_396), .C(n_404), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_414), .B(n_382), .Y(n_459) );
OAI221xp5_ASAP7_75t_L g460 ( .A1(n_417), .A2(n_389), .B1(n_396), .B2(n_375), .C(n_370), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_419), .B(n_396), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_419), .Y(n_462) );
INVx2_ASAP7_75t_SL g463 ( .A(n_436), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_440), .B(n_401), .Y(n_464) );
AO31x2_ASAP7_75t_L g465 ( .A1(n_441), .A2(n_410), .A3(n_409), .B(n_404), .Y(n_465) );
OAI322xp33_ASAP7_75t_L g466 ( .A1(n_440), .A2(n_410), .A3(n_409), .B1(n_365), .B2(n_362), .C1(n_171), .C2(n_21), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_426), .A2(n_405), .B1(n_377), .B2(n_375), .Y(n_467) );
AND2x4_ASAP7_75t_SL g468 ( .A(n_436), .B(n_377), .Y(n_468) );
OAI21xp33_ASAP7_75t_L g469 ( .A1(n_428), .A2(n_405), .B(n_377), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_426), .A2(n_405), .B1(n_377), .B2(n_298), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_429), .A2(n_350), .B1(n_336), .B2(n_373), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_429), .A2(n_373), .B1(n_337), .B2(n_336), .Y(n_472) );
OAI221xp5_ASAP7_75t_SL g473 ( .A1(n_424), .A2(n_337), .B1(n_327), .B2(n_405), .C(n_295), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_426), .A2(n_295), .B1(n_298), .B2(n_337), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_418), .A2(n_300), .B1(n_301), .B2(n_331), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_434), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_438), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_438), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_457), .B(n_441), .Y(n_479) );
AND3x1_ASAP7_75t_L g480 ( .A(n_451), .B(n_422), .C(n_423), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_455), .B(n_387), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_455), .B(n_387), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_445), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_473), .A2(n_436), .B1(n_437), .B2(n_439), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_442), .A2(n_436), .B1(n_421), .B2(n_433), .Y(n_485) );
AND2x4_ASAP7_75t_L g486 ( .A(n_445), .B(n_431), .Y(n_486) );
AOI33xp33_ASAP7_75t_L g487 ( .A1(n_450), .A2(n_13), .A3(n_14), .B1(n_18), .B2(n_19), .B3(n_20), .Y(n_487) );
AOI221xp5_ASAP7_75t_SL g488 ( .A1(n_449), .A2(n_171), .B1(n_207), .B2(n_215), .C(n_243), .Y(n_488) );
BUFx2_ASAP7_75t_L g489 ( .A(n_447), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_456), .A2(n_435), .B1(n_431), .B2(n_281), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_447), .Y(n_491) );
OAI31xp33_ASAP7_75t_L g492 ( .A1(n_456), .A2(n_273), .A3(n_281), .B(n_277), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_477), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_448), .B(n_387), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_476), .B(n_387), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_448), .B(n_387), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_477), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_478), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_462), .B(n_431), .Y(n_499) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_478), .Y(n_500) );
BUFx2_ASAP7_75t_SL g501 ( .A(n_463), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_463), .B(n_345), .Y(n_502) );
INVx1_ASAP7_75t_SL g503 ( .A(n_468), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_462), .B(n_18), .Y(n_504) );
INVxp67_ASAP7_75t_L g505 ( .A(n_464), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_468), .B(n_345), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_443), .B(n_21), .Y(n_507) );
OAI321xp33_ASAP7_75t_L g508 ( .A1(n_446), .A2(n_171), .A3(n_331), .B1(n_345), .B2(n_282), .C(n_304), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_465), .Y(n_509) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_444), .A2(n_282), .B(n_304), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_443), .B(n_22), .Y(n_511) );
OAI31xp33_ASAP7_75t_SL g512 ( .A1(n_452), .A2(n_280), .A3(n_25), .B(n_26), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_465), .Y(n_513) );
OAI21xp33_ASAP7_75t_L g514 ( .A1(n_453), .A2(n_171), .B(n_193), .Y(n_514) );
AOI211xp5_ASAP7_75t_L g515 ( .A1(n_466), .A2(n_273), .B(n_280), .C(n_331), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_443), .B(n_24), .Y(n_516) );
OAI33xp33_ASAP7_75t_L g517 ( .A1(n_459), .A2(n_193), .A3(n_245), .B1(n_244), .B2(n_224), .B3(n_220), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_443), .Y(n_518) );
AND4x1_ASAP7_75t_L g519 ( .A(n_471), .B(n_31), .C(n_32), .D(n_36), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_465), .B(n_345), .Y(n_520) );
INVxp67_ASAP7_75t_L g521 ( .A(n_461), .Y(n_521) );
AND2x4_ASAP7_75t_L g522 ( .A(n_465), .B(n_345), .Y(n_522) );
BUFx3_ASAP7_75t_L g523 ( .A(n_465), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_454), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_444), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_469), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_470), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_467), .Y(n_528) );
INVx1_ASAP7_75t_SL g529 ( .A(n_470), .Y(n_529) );
INVx4_ASAP7_75t_L g530 ( .A(n_466), .Y(n_530) );
NAND4xp25_ASAP7_75t_L g531 ( .A(n_458), .B(n_257), .C(n_277), .D(n_201), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_521), .B(n_460), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_505), .B(n_472), .Y(n_533) );
BUFx3_ASAP7_75t_L g534 ( .A(n_489), .Y(n_534) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_489), .Y(n_535) );
AOI211xp5_ASAP7_75t_L g536 ( .A1(n_512), .A2(n_469), .B(n_474), .C(n_245), .Y(n_536) );
NAND3xp33_ASAP7_75t_SL g537 ( .A(n_487), .B(n_475), .C(n_201), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_503), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_481), .B(n_331), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_479), .B(n_331), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_483), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_504), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_524), .B(n_37), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_524), .B(n_40), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_494), .B(n_41), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_497), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_483), .B(n_43), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_499), .B(n_44), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_504), .Y(n_549) );
NOR3xp33_ASAP7_75t_L g550 ( .A(n_531), .B(n_244), .C(n_187), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_480), .A2(n_277), .B1(n_257), .B2(n_300), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_494), .B(n_47), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_496), .B(n_50), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_491), .B(n_53), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_491), .Y(n_555) );
OAI31xp33_ASAP7_75t_SL g556 ( .A1(n_484), .A2(n_56), .A3(n_58), .B(n_60), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_496), .B(n_64), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_499), .B(n_65), .Y(n_558) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_493), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_493), .Y(n_560) );
OAI211xp5_ASAP7_75t_L g561 ( .A1(n_530), .A2(n_314), .B(n_210), .C(n_187), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_481), .B(n_69), .Y(n_562) );
INVx1_ASAP7_75t_SL g563 ( .A(n_501), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_501), .Y(n_564) );
NAND5xp2_ASAP7_75t_L g565 ( .A(n_492), .B(n_70), .C(n_75), .D(n_76), .E(n_77), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_497), .Y(n_566) );
INVx2_ASAP7_75t_SL g567 ( .A(n_500), .Y(n_567) );
NAND3xp33_ASAP7_75t_L g568 ( .A(n_530), .B(n_243), .C(n_215), .Y(n_568) );
AOI221xp5_ASAP7_75t_L g569 ( .A1(n_530), .A2(n_210), .B1(n_189), .B2(n_203), .C(n_224), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_507), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_507), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_527), .B(n_78), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_495), .B(n_314), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_506), .Y(n_574) );
INVx3_ASAP7_75t_L g575 ( .A(n_500), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_529), .B(n_207), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_511), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_482), .B(n_314), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_523), .B(n_207), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_511), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_482), .B(n_189), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_498), .B(n_203), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_498), .B(n_208), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_486), .B(n_208), .Y(n_584) );
O2A1O1Ixp33_ASAP7_75t_L g585 ( .A1(n_525), .A2(n_220), .B(n_257), .C(n_292), .Y(n_585) );
INVxp67_ASAP7_75t_L g586 ( .A(n_520), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_513), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_509), .Y(n_588) );
INVx2_ASAP7_75t_SL g589 ( .A(n_500), .Y(n_589) );
INVx2_ASAP7_75t_SL g590 ( .A(n_500), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_525), .B(n_314), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_486), .B(n_207), .Y(n_592) );
NOR2x1_ASAP7_75t_L g593 ( .A(n_568), .B(n_523), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_541), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_559), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_586), .B(n_509), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_560), .B(n_500), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_570), .B(n_486), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_561), .A2(n_519), .B(n_515), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_542), .B(n_528), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_555), .Y(n_601) );
NAND2x1p5_ASAP7_75t_L g602 ( .A(n_563), .B(n_548), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_571), .B(n_518), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_549), .Y(n_604) );
NOR2xp67_ASAP7_75t_L g605 ( .A(n_564), .B(n_508), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_535), .Y(n_606) );
NAND2xp33_ASAP7_75t_L g607 ( .A(n_564), .B(n_485), .Y(n_607) );
OAI31xp33_ASAP7_75t_L g608 ( .A1(n_565), .A2(n_528), .A3(n_526), .B(n_516), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_538), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_577), .B(n_518), .Y(n_610) );
NOR2x1_ASAP7_75t_R g611 ( .A(n_548), .B(n_516), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_580), .B(n_490), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_532), .B(n_522), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_587), .Y(n_614) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_534), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_532), .B(n_522), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_581), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_588), .B(n_526), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_581), .B(n_510), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_539), .B(n_506), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_588), .B(n_502), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_534), .B(n_506), .Y(n_622) );
BUFx2_ASAP7_75t_L g623 ( .A(n_592), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_546), .B(n_502), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g625 ( .A1(n_562), .A2(n_488), .B(n_514), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_533), .B(n_517), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_566), .Y(n_627) );
NAND3xp33_ASAP7_75t_SL g628 ( .A(n_536), .B(n_314), .C(n_252), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_578), .B(n_207), .Y(n_629) );
NAND3xp33_ASAP7_75t_SL g630 ( .A(n_572), .B(n_252), .C(n_300), .Y(n_630) );
INVx1_ASAP7_75t_SL g631 ( .A(n_574), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_562), .B(n_215), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_566), .B(n_215), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_573), .B(n_215), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_592), .B(n_243), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_540), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_552), .B(n_243), .Y(n_637) );
NAND4xp25_ASAP7_75t_SL g638 ( .A(n_553), .B(n_252), .C(n_301), .D(n_274), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_567), .B(n_301), .Y(n_639) );
INVx2_ASAP7_75t_SL g640 ( .A(n_579), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_591), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_553), .B(n_301), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_556), .B(n_252), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_594), .Y(n_644) );
OAI21xp5_ASAP7_75t_L g645 ( .A1(n_628), .A2(n_537), .B(n_585), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_595), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_614), .B(n_584), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_606), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_604), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_601), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_603), .B(n_584), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_636), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_607), .A2(n_616), .B1(n_613), .B2(n_641), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_615), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_623), .B(n_575), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_618), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_603), .B(n_558), .Y(n_657) );
XNOR2xp5_ASAP7_75t_L g658 ( .A(n_609), .B(n_557), .Y(n_658) );
OAI21xp5_ASAP7_75t_SL g659 ( .A1(n_608), .A2(n_554), .B(n_547), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_631), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_600), .Y(n_661) );
INVx3_ASAP7_75t_L g662 ( .A(n_602), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_617), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_598), .B(n_545), .Y(n_664) );
AND2x4_ASAP7_75t_L g665 ( .A(n_640), .B(n_567), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_598), .B(n_576), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_605), .B(n_579), .Y(n_667) );
OR2x2_ASAP7_75t_L g668 ( .A(n_596), .B(n_590), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_610), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_627), .Y(n_670) );
INVx1_ASAP7_75t_SL g671 ( .A(n_615), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_618), .Y(n_672) );
OAI22xp33_ASAP7_75t_L g673 ( .A1(n_602), .A2(n_544), .B1(n_543), .B2(n_589), .Y(n_673) );
NOR2x1_ASAP7_75t_L g674 ( .A(n_630), .B(n_579), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_612), .Y(n_675) );
INVx2_ASAP7_75t_SL g676 ( .A(n_640), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_624), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_626), .B(n_576), .Y(n_678) );
OR2x2_ASAP7_75t_L g679 ( .A(n_620), .B(n_590), .Y(n_679) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_597), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_624), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_607), .A2(n_611), .B(n_599), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_619), .A2(n_589), .B1(n_575), .B2(n_569), .C(n_583), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_625), .B(n_551), .C(n_575), .Y(n_684) );
OA22x2_ASAP7_75t_L g685 ( .A1(n_643), .A2(n_583), .B1(n_582), .B2(n_550), .Y(n_685) );
XOR2xp5_ASAP7_75t_L g686 ( .A(n_622), .B(n_292), .Y(n_686) );
OAI21xp5_ASAP7_75t_SL g687 ( .A1(n_643), .A2(n_274), .B(n_253), .Y(n_687) );
OAI22xp33_ASAP7_75t_L g688 ( .A1(n_593), .A2(n_252), .B1(n_274), .B2(n_268), .Y(n_688) );
OAI21xp33_ASAP7_75t_SL g689 ( .A1(n_638), .A2(n_253), .B(n_268), .Y(n_689) );
INVxp67_ASAP7_75t_L g690 ( .A(n_621), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_629), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_635), .B(n_633), .Y(n_692) );
XNOR2xp5_ASAP7_75t_L g693 ( .A(n_637), .B(n_642), .Y(n_693) );
OAI21xp5_ASAP7_75t_SL g694 ( .A1(n_632), .A2(n_634), .B(n_639), .Y(n_694) );
XNOR2xp5_ASAP7_75t_L g695 ( .A(n_633), .B(n_639), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_594), .Y(n_696) );
INVx1_ASAP7_75t_SL g697 ( .A(n_609), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_602), .A2(n_564), .B1(n_605), .B2(n_530), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_594), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_594), .Y(n_700) );
OAI22x1_ASAP7_75t_L g701 ( .A1(n_697), .A2(n_667), .B1(n_660), .B2(n_653), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_680), .Y(n_702) );
NOR3xp33_ASAP7_75t_SL g703 ( .A(n_682), .B(n_698), .C(n_659), .Y(n_703) );
INVxp67_ASAP7_75t_SL g704 ( .A(n_654), .Y(n_704) );
AOI32xp33_ASAP7_75t_L g705 ( .A1(n_667), .A2(n_671), .A3(n_674), .B1(n_676), .B2(n_662), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_685), .A2(n_675), .B1(n_687), .B2(n_694), .Y(n_706) );
OAI21xp5_ASAP7_75t_L g707 ( .A1(n_685), .A2(n_687), .B(n_645), .Y(n_707) );
A2O1A1Ixp33_ASAP7_75t_L g708 ( .A1(n_689), .A2(n_694), .B(n_676), .C(n_654), .Y(n_708) );
XNOR2xp5_ASAP7_75t_L g709 ( .A(n_658), .B(n_693), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_695), .A2(n_684), .B(n_678), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_651), .A2(n_690), .B1(n_662), .B2(n_680), .Y(n_711) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_661), .Y(n_712) );
NAND2x1_ASAP7_75t_L g713 ( .A(n_665), .B(n_656), .Y(n_713) );
AOI211xp5_ASAP7_75t_L g714 ( .A1(n_673), .A2(n_683), .B(n_691), .C(n_688), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_656), .Y(n_715) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_712), .Y(n_716) );
NOR3xp33_ASAP7_75t_L g717 ( .A(n_707), .B(n_673), .C(n_646), .Y(n_717) );
AOI32xp33_ASAP7_75t_L g718 ( .A1(n_711), .A2(n_665), .A3(n_655), .B1(n_652), .B2(n_648), .Y(n_718) );
NOR4xp25_ASAP7_75t_L g719 ( .A(n_708), .B(n_644), .C(n_699), .D(n_696), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_701), .A2(n_700), .B1(n_669), .B2(n_649), .C(n_650), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_705), .A2(n_663), .B1(n_672), .B2(n_647), .C(n_677), .Y(n_721) );
OAI211xp5_ASAP7_75t_SL g722 ( .A1(n_703), .A2(n_657), .B(n_666), .C(n_664), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_706), .A2(n_692), .B1(n_665), .B2(n_686), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_709), .B(n_681), .Y(n_724) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_716), .Y(n_725) );
OAI22xp33_ASAP7_75t_SL g726 ( .A1(n_724), .A2(n_706), .B1(n_713), .B2(n_704), .Y(n_726) );
OAI211xp5_ASAP7_75t_SL g727 ( .A1(n_723), .A2(n_714), .B(n_710), .C(n_702), .Y(n_727) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_717), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_722), .B(n_715), .Y(n_729) );
NAND3xp33_ASAP7_75t_L g730 ( .A(n_728), .B(n_720), .C(n_721), .Y(n_730) );
XOR2xp5_ASAP7_75t_L g731 ( .A(n_725), .B(n_679), .Y(n_731) );
OR2x2_ASAP7_75t_L g732 ( .A(n_729), .B(n_719), .Y(n_732) );
INVx4_ASAP7_75t_L g733 ( .A(n_732), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_731), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_734), .A2(n_727), .B1(n_730), .B2(n_726), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_733), .A2(n_718), .B1(n_668), .B2(n_670), .Y(n_736) );
INVxp67_ASAP7_75t_L g737 ( .A(n_735), .Y(n_737) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_737), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_738), .A2(n_733), .B(n_736), .Y(n_739) );
endmodule