module fake_ariane_975_n_184 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_184);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_184;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_30;
wire n_82;
wire n_178;
wire n_42;
wire n_31;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_144;
wire n_130;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_121;
wire n_118;
wire n_93;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_125;
wire n_168;
wire n_43;
wire n_87;
wire n_81;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_21),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVxp67_ASAP7_75t_SL g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_29),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_51),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_0),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_1),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_30),
.B(n_2),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_3),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_34),
.B(n_3),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_4),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_5),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_43),
.B(n_37),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_34),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_57),
.B(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

AND3x1_ASAP7_75t_SL g80 ( 
.A(n_66),
.B(n_48),
.C(n_46),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_36),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

OR2x6_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_43),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_52),
.Y(n_85)
);

AND2x4_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_48),
.Y(n_86)
);

NAND3xp33_ASAP7_75t_SL g87 ( 
.A(n_62),
.B(n_45),
.C(n_44),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_58),
.B(n_32),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_58),
.B(n_31),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_76),
.B(n_69),
.Y(n_91)
);

AO32x2_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_52),
.A3(n_54),
.B1(n_68),
.B2(n_65),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_54),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_55),
.B(n_64),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_69),
.B(n_73),
.Y(n_95)
);

NAND2x1_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_63),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_52),
.Y(n_97)
);

AO32x2_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_68),
.A3(n_65),
.B1(n_70),
.B2(n_53),
.Y(n_98)
);

INVxp67_ASAP7_75t_SL g99 ( 
.A(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

AOI221x1_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_64),
.B1(n_59),
.B2(n_60),
.C(n_63),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_83),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_72),
.B(n_74),
.C(n_83),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_95),
.A2(n_84),
.B1(n_49),
.B2(n_38),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_84),
.B1(n_83),
.B2(n_82),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_101),
.A2(n_84),
.B(n_90),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_84),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_87),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_98),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_89),
.Y(n_116)
);

OA21x2_ASAP7_75t_L g117 ( 
.A1(n_115),
.A2(n_103),
.B(n_107),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_98),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

OA21x2_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_53),
.B(n_71),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_112),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_98),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_98),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_98),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_119),
.Y(n_130)
);

A2O1A1O1Ixp25_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_37),
.B(n_46),
.C(n_72),
.D(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

OAI221xp5_ASAP7_75t_L g133 ( 
.A1(n_123),
.A2(n_70),
.B1(n_116),
.B2(n_78),
.C(n_109),
.Y(n_133)
);

OAI221xp5_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_109),
.B1(n_114),
.B2(n_66),
.C(n_67),
.Y(n_134)
);

AOI32xp33_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_59),
.A3(n_60),
.B1(n_63),
.B2(n_67),
.Y(n_135)
);

AOI21xp33_ASAP7_75t_SL g136 ( 
.A1(n_122),
.A2(n_60),
.B(n_59),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_119),
.B(n_96),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_118),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_108),
.B1(n_114),
.B2(n_77),
.Y(n_140)
);

AOI221xp5_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_61),
.B1(n_71),
.B2(n_129),
.C(n_127),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_117),
.B(n_132),
.Y(n_142)
);

OAI221xp5_ASAP7_75t_L g143 ( 
.A1(n_135),
.A2(n_131),
.B1(n_61),
.B2(n_71),
.C(n_117),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_117),
.B(n_132),
.Y(n_144)
);

OAI221xp5_ASAP7_75t_L g145 ( 
.A1(n_140),
.A2(n_61),
.B1(n_71),
.B2(n_117),
.C(n_129),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_127),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_136),
.A2(n_117),
.B(n_118),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_128),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_117),
.B(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_146),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_148),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_5),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_SL g153 ( 
.A1(n_149),
.A2(n_126),
.B(n_125),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_144),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_117),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_117),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_126),
.B1(n_68),
.B2(n_65),
.Y(n_160)
);

NAND2x1p5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_120),
.Y(n_161)
);

AOI311xp33_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_6),
.A3(n_7),
.B(n_8),
.C(n_9),
.Y(n_162)
);

OAI211xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_152),
.B(n_154),
.C(n_157),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_156),
.B(n_120),
.Y(n_164)
);

NAND4xp75_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_120),
.C(n_75),
.D(n_77),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_120),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_155),
.C(n_96),
.Y(n_167)
);

AOI221xp5_ASAP7_75t_L g168 ( 
.A1(n_159),
.A2(n_81),
.B1(n_86),
.B2(n_8),
.C(n_9),
.Y(n_168)
);

OAI221xp5_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_159),
.B1(n_160),
.B2(n_166),
.C(n_161),
.Y(n_169)
);

OAI221xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_120),
.B1(n_81),
.B2(n_10),
.C(n_11),
.Y(n_170)
);

AOI221xp5_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_81),
.B1(n_86),
.B2(n_10),
.C(n_12),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_6),
.A3(n_7),
.B1(n_13),
.B2(n_14),
.C1(n_16),
.C2(n_92),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_169),
.Y(n_173)
);

OAI211xp5_ASAP7_75t_SL g174 ( 
.A1(n_171),
.A2(n_164),
.B(n_85),
.C(n_161),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_167),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_170),
.A2(n_120),
.B(n_165),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_172),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_23),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_178),
.A2(n_92),
.B1(n_93),
.B2(n_99),
.Y(n_180)
);

NOR3xp33_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_92),
.C(n_27),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_175),
.B(n_174),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_175),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_183),
.A2(n_182),
.B1(n_181),
.B2(n_177),
.Y(n_184)
);


endmodule