module real_jpeg_33940_n_20 (n_17, n_649, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_649;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_578;
wire n_149;
wire n_620;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_611;
wire n_221;
wire n_393;
wire n_489;
wire n_634;
wire n_153;
wire n_104;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_642;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_641;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_0),
.Y(n_78)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_0),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_0),
.Y(n_339)
);

BUFx12f_ASAP7_75t_L g472 ( 
.A(n_0),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_1),
.A2(n_196),
.B1(n_197),
.B2(n_199),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_1),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_1),
.A2(n_196),
.B1(n_209),
.B2(n_212),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_1),
.A2(n_196),
.B1(n_226),
.B2(n_230),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_1),
.A2(n_196),
.B1(n_341),
.B2(n_344),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_2),
.A2(n_93),
.B1(n_96),
.B2(n_101),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_2),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_2),
.A2(n_101),
.B1(n_241),
.B2(n_244),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_2),
.A2(n_101),
.B1(n_142),
.B2(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_2),
.A2(n_101),
.B1(n_331),
.B2(n_333),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_3),
.Y(n_109)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_3),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_4),
.A2(n_50),
.B1(n_56),
.B2(n_60),
.Y(n_49)
);

INVx2_ASAP7_75t_R g60 ( 
.A(n_4),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_4),
.A2(n_60),
.B1(n_153),
.B2(n_156),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_4),
.A2(n_60),
.B1(n_370),
.B2(n_373),
.Y(n_369)
);

AO22x1_ASAP7_75t_L g621 ( 
.A1(n_4),
.A2(n_60),
.B1(n_357),
.B2(n_622),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_5),
.A2(n_301),
.B1(n_304),
.B2(n_308),
.Y(n_300)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_5),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_5),
.A2(n_308),
.B1(n_397),
.B2(n_400),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g464 ( 
.A1(n_5),
.A2(n_308),
.B1(n_465),
.B2(n_467),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_5),
.A2(n_308),
.B1(n_540),
.B2(n_542),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_6),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_7),
.A2(n_270),
.B1(n_271),
.B2(n_274),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_7),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_7),
.A2(n_270),
.B1(n_320),
.B2(n_323),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_7),
.A2(n_270),
.B1(n_458),
.B2(n_461),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_7),
.A2(n_270),
.B1(n_521),
.B2(n_522),
.Y(n_520)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_8),
.A2(n_117),
.B1(n_121),
.B2(n_122),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_8),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_8),
.A2(n_121),
.B1(n_290),
.B2(n_293),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_8),
.A2(n_121),
.B1(n_404),
.B2(n_406),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_8),
.A2(n_121),
.B1(n_333),
.B2(n_534),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_9),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_9),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_9),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_10),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_10),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_11),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_11),
.Y(n_345)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_11),
.Y(n_491)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_12),
.Y(n_507)
);

CKINVDCx11_ASAP7_75t_R g639 ( 
.A(n_13),
.Y(n_639)
);

CKINVDCx11_ASAP7_75t_R g647 ( 
.A(n_13),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_14),
.A2(n_277),
.B(n_279),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_14),
.B(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_14),
.Y(n_347)
);

OAI22xp33_ASAP7_75t_SL g475 ( 
.A1(n_14),
.A2(n_75),
.B1(n_235),
.B2(n_457),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_14),
.B(n_190),
.Y(n_536)
);

OAI32xp33_ASAP7_75t_L g553 ( 
.A1(n_14),
.A2(n_167),
.A3(n_554),
.B1(n_557),
.B2(n_558),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_14),
.A2(n_347),
.B1(n_568),
.B2(n_571),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_15),
.A2(n_251),
.B1(n_255),
.B2(n_256),
.Y(n_250)
);

INVx2_ASAP7_75t_R g255 ( 
.A(n_15),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_15),
.A2(n_255),
.B1(n_310),
.B2(n_315),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_15),
.A2(n_255),
.B1(n_487),
.B2(n_492),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_15),
.A2(n_255),
.B1(n_575),
.B2(n_578),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_16),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_16),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_16),
.A2(n_87),
.B1(n_142),
.B2(n_145),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g627 ( 
.A1(n_16),
.A2(n_87),
.B1(n_153),
.B2(n_179),
.Y(n_627)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_18),
.A2(n_65),
.B1(n_70),
.B2(n_71),
.Y(n_64)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_18),
.A2(n_70),
.B1(n_179),
.B2(n_183),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_18),
.A2(n_70),
.B1(n_85),
.B2(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_19),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_19),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_19),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_19),
.Y(n_188)
);

OAI321xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_260),
.A3(n_261),
.B1(n_610),
.B2(n_641),
.C(n_646),
.Y(n_20)
);

AOI322xp5_ASAP7_75t_L g646 ( 
.A1(n_21),
.A2(n_611),
.A3(n_634),
.B1(n_642),
.B2(n_643),
.C1(n_647),
.C2(n_649),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_215),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_23),
.B(n_215),
.Y(n_645)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_191),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_136),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_25),
.B(n_630),
.C(n_631),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_74),
.B(n_88),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_26),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_74),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_27),
.A2(n_74),
.B1(n_220),
.B2(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_27),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_49),
.B1(n_61),
.B2(n_64),
.Y(n_27)
);

AO21x1_ASAP7_75t_L g139 ( 
.A1(n_28),
.A2(n_140),
.B(n_141),
.Y(n_139)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_28),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_28),
.A2(n_49),
.B1(n_61),
.B2(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_28),
.A2(n_140),
.B1(n_285),
.B2(n_289),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_28),
.A2(n_140),
.B1(n_225),
.B2(n_285),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_28),
.A2(n_140),
.B1(n_538),
.B2(n_539),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_28),
.A2(n_591),
.B(n_592),
.Y(n_590)
);

AO21x2_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_37),
.B(n_41),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_34),
.Y(n_288)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_36),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_36),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_37),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_43),
.Y(n_332)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_43),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_43),
.Y(n_513)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_44),
.Y(n_343)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_53),
.Y(n_521)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_55),
.Y(n_519)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_58),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_59),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_59),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_62),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_62),
.A2(n_204),
.B1(n_574),
.B2(n_581),
.Y(n_573)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_64),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_69),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_69),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_69),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_69),
.Y(n_541)
);

BUFx6f_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_74),
.A2(n_89),
.B1(n_90),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_74),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_79),
.B(n_84),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_75),
.A2(n_84),
.B1(n_232),
.B2(n_235),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_75),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_75),
.A2(n_232),
.B1(n_369),
.B2(n_384),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_75),
.A2(n_457),
.B1(n_464),
.B2(n_471),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_75),
.A2(n_486),
.B1(n_494),
.B2(n_532),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_76),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx4f_ASAP7_75t_L g479 ( 
.A(n_78),
.Y(n_479)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_83),
.Y(n_387)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_115),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_102),
.Y(n_91)
);

AO22x1_ASAP7_75t_L g206 ( 
.A1(n_92),
.A2(n_125),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_99),
.Y(n_211)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_99),
.Y(n_399)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_100),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_103),
.Y(n_207)
);

OAI22x1_ASAP7_75t_SL g248 ( 
.A1(n_103),
.A2(n_249),
.B1(n_250),
.B2(n_259),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_103),
.A2(n_249),
.B1(n_269),
.B2(n_276),
.Y(n_268)
);

NOR2xp67_ASAP7_75t_SL g346 ( 
.A(n_103),
.B(n_347),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_103),
.A2(n_249),
.B1(n_250),
.B2(n_396),
.Y(n_419)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_103),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_108),
.B1(n_110),
.B2(n_112),
.Y(n_104)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_106),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g303 ( 
.A(n_107),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_107),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_107),
.Y(n_314)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_108),
.Y(n_361)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_109),
.Y(n_356)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_110),
.Y(n_316)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_110),
.Y(n_352)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_125),
.Y(n_115)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_116),
.Y(n_259)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_120),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_120),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_120),
.Y(n_624)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_125),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_125),
.A2(n_207),
.B1(n_394),
.B2(n_395),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g630 ( 
.A1(n_136),
.A2(n_137),
.B1(n_206),
.B2(n_615),
.Y(n_630)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_149),
.B2(n_150),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_138),
.B(n_150),
.C(n_615),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_138),
.A2(n_139),
.B1(n_626),
.B2(n_628),
.Y(n_625)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_140),
.B(n_347),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_140),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_141),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_144),
.Y(n_523)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_147),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_148),
.Y(n_560)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_148),
.Y(n_580)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_160),
.B1(n_178),
.B2(n_189),
.Y(n_150)
);

INVxp67_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_152),
.A2(n_190),
.B1(n_195),
.B2(n_201),
.Y(n_194)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_158),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_159),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_160),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_160),
.A2(n_189),
.B1(n_300),
.B2(n_309),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_160),
.A2(n_189),
.B1(n_300),
.B2(n_319),
.Y(n_318)
);

OA22x2_ASAP7_75t_L g402 ( 
.A1(n_160),
.A2(n_189),
.B1(n_309),
.B2(n_403),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_160),
.A2(n_189),
.B1(n_240),
.B2(n_403),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_160),
.A2(n_189),
.B1(n_319),
.B2(n_567),
.Y(n_566)
);

OAI22xp33_ASAP7_75t_SL g626 ( 
.A1(n_160),
.A2(n_178),
.B1(n_189),
.B2(n_627),
.Y(n_626)
);

AO21x2_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_167),
.B(n_171),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_SL g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_165),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_185),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_187),
.Y(n_322)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_187),
.Y(n_405)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_190),
.A2(n_195),
.B1(n_201),
.B2(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_206),
.Y(n_191)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_192),
.Y(n_631)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OA21x2_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_194),
.B(n_202),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_202),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_204),
.A2(n_516),
.B1(n_520),
.B2(n_524),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_206),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_206),
.B(n_618),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_SL g618 ( 
.A1(n_208),
.A2(n_619),
.B1(n_620),
.B2(n_621),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_212),
.Y(n_400)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_214),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_221),
.C(n_222),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_217),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_218),
.B(n_221),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_222),
.B(n_429),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_237),
.C(n_247),
.Y(n_222)
);

XNOR2x1_ASAP7_75t_L g423 ( 
.A(n_223),
.B(n_424),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_231),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_224),
.B(n_231),
.Y(n_441)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVxp33_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_238),
.B(n_248),
.Y(n_424)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_243),
.Y(n_326)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_243),
.Y(n_364)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_249),
.Y(n_619)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx3_ASAP7_75t_SL g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx4f_ASAP7_75t_SL g278 ( 
.A(n_258),
.Y(n_278)
);

BUFx12f_ASAP7_75t_L g358 ( 
.A(n_258),
.Y(n_358)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_449),
.B(n_605),
.Y(n_262)
);

NAND4xp25_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_410),
.C(n_430),
.D(n_443),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_380),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_265),
.B(n_380),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_317),
.C(n_348),
.Y(n_265)
);

XOR2x2_ASAP7_75t_L g601 ( 
.A(n_266),
.B(n_602),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_283),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

MAJx2_ASAP7_75t_L g389 ( 
.A(n_268),
.B(n_284),
.C(n_299),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_269),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_273),
.Y(n_282)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_279),
.Y(n_365)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_299),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVxp33_ASAP7_75t_L g593 ( 
.A(n_289),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_297),
.Y(n_511)
);

INVx5_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_303),
.Y(n_570)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_307),
.Y(n_572)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_317),
.B(n_348),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_327),
.C(n_346),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_318),
.B(n_597),
.Y(n_596)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_327),
.A2(n_328),
.B1(n_346),
.B2(n_598),
.Y(n_597)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_330),
.B1(n_337),
.B2(n_340),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_329),
.A2(n_340),
.B1(n_367),
.B2(n_368),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_329),
.A2(n_484),
.B1(n_485),
.B2(n_493),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_329),
.A2(n_330),
.B1(n_533),
.B2(n_562),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_336),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_336),
.Y(n_460)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_336),
.Y(n_463)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_336),
.Y(n_470)
);

BUFx2_ASAP7_75t_R g337 ( 
.A(n_338),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_338),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_339),
.Y(n_367)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_345),
.Y(n_376)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_345),
.Y(n_503)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_346),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_347),
.B(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_347),
.B(n_510),
.Y(n_509)
);

OAI21xp33_ASAP7_75t_SL g516 ( 
.A1(n_347),
.A2(n_509),
.B(n_517),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_347),
.B(n_559),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_349),
.A2(n_366),
.B1(n_377),
.B2(n_379),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_349),
.B(n_379),
.Y(n_409)
);

OAI32xp33_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_353),
.A3(n_357),
.B1(n_359),
.B2(n_365),
.Y(n_349)
);

OAI32xp33_ASAP7_75t_L g378 ( 
.A1(n_350),
.A2(n_353),
.A3(n_357),
.B1(n_359),
.B2(n_365),
.Y(n_378)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_SL g351 ( 
.A(n_352),
.Y(n_351)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx11_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_362),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_366),
.Y(n_379)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_372),
.Y(n_534)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_390),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_389),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_382),
.B(n_390),
.C(n_432),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_388),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_383),
.B(n_388),
.Y(n_417)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g386 ( 
.A(n_387),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_389),
.Y(n_432)
);

XNOR2x1_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_409),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_392),
.A2(n_393),
.B1(n_401),
.B2(n_402),
.Y(n_391)
);

MAJx2_ASAP7_75t_L g435 ( 
.A(n_392),
.B(n_409),
.C(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVxp33_ASAP7_75t_L g436 ( 
.A(n_402),
.Y(n_436)
);

INVx2_ASAP7_75t_SL g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

A2O1A1O1Ixp25_ASAP7_75t_L g605 ( 
.A1(n_410),
.A2(n_443),
.B(n_606),
.C(n_608),
.D(n_609),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_428),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_411),
.B(n_428),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_422),
.B(n_425),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_415),
.Y(n_412)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_413),
.Y(n_427)
);

INVxp33_ASAP7_75t_SL g426 ( 
.A(n_415),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_415),
.B(n_448),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_418),
.C(n_420),
.Y(n_415)
);

OAI22xp33_ASAP7_75t_SL g446 ( 
.A1(n_416),
.A2(n_417),
.B1(n_438),
.B2(n_442),
.Y(n_446)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_417),
.B(n_441),
.Y(n_440)
);

AO22x1_ASAP7_75t_L g438 ( 
.A1(n_418),
.A2(n_419),
.B1(n_420),
.B2(n_421),
.Y(n_438)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_423),
.B(n_427),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_433),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_431),
.B(n_433),
.C(n_607),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_437),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_435),
.B(n_445),
.C(n_446),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_438),
.A2(n_439),
.B1(n_440),
.B2(n_442),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_438),
.Y(n_442)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVxp33_ASAP7_75t_SL g445 ( 
.A(n_441),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_447),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_444),
.B(n_447),
.Y(n_608)
);

AOI21x1_ASAP7_75t_L g449 ( 
.A1(n_450),
.A2(n_600),
.B(n_604),
.Y(n_449)
);

OAI21x1_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_585),
.B(n_599),
.Y(n_450)
);

AOI21x1_ASAP7_75t_L g451 ( 
.A1(n_452),
.A2(n_549),
.B(n_584),
.Y(n_451)
);

OAI21x1_ASAP7_75t_L g452 ( 
.A1(n_453),
.A2(n_528),
.B(n_548),
.Y(n_452)
);

AOI22x1_ASAP7_75t_SL g453 ( 
.A1(n_454),
.A2(n_482),
.B1(n_526),
.B2(n_527),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_455),
.A2(n_474),
.B(n_481),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_473),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_456),
.B(n_473),
.Y(n_481)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_460),
.Y(n_492)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_461),
.Y(n_480)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_464),
.Y(n_484)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_471),
.Y(n_562)
);

INVx4_ASAP7_75t_SL g471 ( 
.A(n_472),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_476),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_477),
.B(n_480),
.Y(n_476)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_497),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_483),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_497),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_498),
.A2(n_499),
.B1(n_515),
.B2(n_525),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_498),
.B(n_525),
.Y(n_529)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_508),
.B1(n_512),
.B2(n_514),
.Y(n_499)
);

NAND2xp33_ASAP7_75t_SL g500 ( 
.A(n_501),
.B(n_504),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_502),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_515),
.Y(n_525)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_519),
.Y(n_557)
);

INVx5_ASAP7_75t_L g577 ( 
.A(n_519),
.Y(n_577)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_520),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_524),
.B(n_593),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_530),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_529),
.B(n_530),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_535),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_531),
.B(n_537),
.C(n_546),
.Y(n_550)
);

INVxp33_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_536),
.A2(n_537),
.B1(n_546),
.B2(n_547),
.Y(n_535)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_536),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_537),
.Y(n_547)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_539),
.Y(n_581)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_550),
.B(n_551),
.Y(n_549)
);

NOR2xp67_ASAP7_75t_SL g584 ( 
.A(n_550),
.B(n_551),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_552),
.B(n_565),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_552),
.B(n_573),
.C(n_583),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_553),
.A2(n_561),
.B1(n_563),
.B2(n_564),
.Y(n_552)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_553),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_553),
.B(n_564),
.Y(n_595)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_561),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_566),
.A2(n_573),
.B1(n_582),
.B2(n_583),
.Y(n_565)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_566),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_569),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_573),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_574),
.Y(n_591)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_577),
.Y(n_576)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

NOR2xp67_ASAP7_75t_L g585 ( 
.A(n_586),
.B(n_587),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_586),
.B(n_587),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_SL g587 ( 
.A(n_588),
.B(n_596),
.Y(n_587)
);

OA22x2_ASAP7_75t_L g588 ( 
.A1(n_589),
.A2(n_590),
.B1(n_594),
.B2(n_595),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_590),
.B(n_594),
.C(n_596),
.Y(n_603)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_601),
.B(n_603),
.Y(n_600)
);

NOR2x1_ASAP7_75t_L g604 ( 
.A(n_601),
.B(n_603),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_L g610 ( 
.A(n_611),
.B(n_634),
.Y(n_610)
);

NOR3xp33_ASAP7_75t_L g642 ( 
.A(n_611),
.B(n_635),
.C(n_643),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_R g611 ( 
.A(n_612),
.B(n_632),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g612 ( 
.A(n_613),
.B(n_629),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_613),
.B(n_629),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_614),
.B(n_616),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_617),
.B(n_625),
.Y(n_616)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_623),
.Y(n_622)
);

INVxp67_ASAP7_75t_SL g623 ( 
.A(n_624),
.Y(n_623)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_626),
.Y(n_628)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_633),
.Y(n_632)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_635),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_636),
.B(n_640),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_637),
.Y(n_636)
);

BUFx10_ASAP7_75t_L g637 ( 
.A(n_638),
.Y(n_637)
);

BUFx12f_ASAP7_75t_L g638 ( 
.A(n_639),
.Y(n_638)
);

INVxp67_ASAP7_75t_SL g641 ( 
.A(n_642),
.Y(n_641)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_644),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_645),
.Y(n_644)
);


endmodule