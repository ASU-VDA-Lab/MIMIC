module fake_ariane_1866_n_1971 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1971);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1971;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_212;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1910;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_205),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_149),
.Y(n_208)
);

BUFx2_ASAP7_75t_SL g209 ( 
.A(n_134),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_105),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_39),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_141),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_77),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_126),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_191),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_1),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_139),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_167),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_35),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_43),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_138),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_204),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_60),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_64),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_195),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_23),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_57),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_15),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_88),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_162),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_19),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_189),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_97),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_99),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_51),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_69),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_109),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_161),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_30),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_85),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_78),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_5),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_202),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_102),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_172),
.Y(n_246)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_5),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_54),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_56),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_180),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_17),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_168),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_30),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_18),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_96),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_44),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_200),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_106),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_187),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_132),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_81),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_49),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_64),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_192),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_74),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_153),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_197),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_41),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_36),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_117),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_166),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_1),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_158),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_128),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_193),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_179),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_40),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_131),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_4),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_116),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_177),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_137),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_38),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_27),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_186),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_4),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_121),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_206),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_58),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_147),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_49),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_136),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_56),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_68),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_157),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_40),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_151),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_79),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_199),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_188),
.Y(n_300)
);

INVxp67_ASAP7_75t_R g301 ( 
.A(n_21),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_10),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_39),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_140),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_113),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_16),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_83),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_154),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_17),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_32),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_120),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_115),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_65),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_201),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_95),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_51),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_181),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_26),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_20),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_129),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_69),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_35),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_175),
.Y(n_323)
);

BUFx10_ASAP7_75t_L g324 ( 
.A(n_58),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_190),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_82),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_164),
.Y(n_327)
);

BUFx10_ASAP7_75t_L g328 ( 
.A(n_11),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_114),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_46),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_87),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_152),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_171),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_101),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_75),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_29),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_107),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_93),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_110),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_26),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_41),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_16),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_6),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_44),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_50),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_144),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_142),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_57),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_13),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_65),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_48),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_135),
.Y(n_352)
);

BUFx10_ASAP7_75t_L g353 ( 
.A(n_169),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_183),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_163),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_198),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_176),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_184),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_34),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_3),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_6),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_32),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_86),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_150),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_130),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_66),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_68),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_174),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_23),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_194),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_123),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_143),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_19),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_24),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_133),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_108),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_54),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_111),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_94),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_18),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_21),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_63),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_50),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_47),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_25),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_53),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_90),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_203),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_160),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_45),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_148),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_10),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_7),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_92),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_60),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_73),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_55),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_48),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_196),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_8),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_52),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_14),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_42),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_155),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_122),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_59),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_112),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_119),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_22),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_62),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_84),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_385),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_247),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_247),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_247),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_247),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_225),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_359),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_245),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_260),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_247),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_247),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_261),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_247),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_271),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_247),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_385),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_254),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_254),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_254),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_254),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_213),
.B(n_0),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_254),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_280),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_314),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_343),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_343),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_343),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_333),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_338),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_343),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_343),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_344),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_346),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_344),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_344),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_358),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_344),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_344),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_324),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_365),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_388),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_221),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_389),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_227),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_391),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_232),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_228),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_232),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_324),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_336),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_324),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_336),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_265),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_360),
.Y(n_465)
);

INVxp33_ASAP7_75t_SL g466 ( 
.A(n_301),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_360),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_268),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_384),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_212),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_328),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_384),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_393),
.Y(n_473)
);

CKINVDCx14_ASAP7_75t_R g474 ( 
.A(n_331),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_269),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_328),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_393),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_272),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_279),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_208),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_303),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_369),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_208),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_217),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_217),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_234),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_222),
.B(n_0),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_256),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_328),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_410),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_262),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_231),
.B(n_2),
.Y(n_492)
);

INVxp33_ASAP7_75t_SL g493 ( 
.A(n_211),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_212),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_277),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_234),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_275),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_275),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_283),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_R g500 ( 
.A(n_257),
.B(n_125),
.Y(n_500)
);

INVxp33_ASAP7_75t_SL g501 ( 
.A(n_211),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_276),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_216),
.Y(n_503)
);

INVxp33_ASAP7_75t_L g504 ( 
.A(n_284),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_276),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_230),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_289),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_276),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_300),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_300),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_353),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_337),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_294),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_296),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_306),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_309),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_506),
.B(n_239),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_438),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_438),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_438),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_422),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_461),
.B(n_353),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_448),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_417),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_422),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_448),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_465),
.B(n_353),
.Y(n_527)
);

INVx6_ASAP7_75t_L g528 ( 
.A(n_506),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_418),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_448),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_413),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_413),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_414),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_470),
.B(n_238),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_414),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_415),
.Y(n_536)
);

INVx5_ASAP7_75t_L g537 ( 
.A(n_441),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_415),
.Y(n_538)
);

OA21x2_ASAP7_75t_L g539 ( 
.A1(n_416),
.A2(n_246),
.B(n_241),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_441),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_416),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_421),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_419),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_421),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_468),
.B(n_207),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_424),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_424),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_426),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_426),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_466),
.B(n_255),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_SL g551 ( 
.A(n_502),
.B(n_216),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_428),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_470),
.B(n_252),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_428),
.Y(n_554)
);

OA21x2_ASAP7_75t_L g555 ( 
.A1(n_429),
.A2(n_278),
.B(n_267),
.Y(n_555)
);

NAND2xp33_ASAP7_75t_L g556 ( 
.A(n_475),
.B(n_310),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_429),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_494),
.B(n_282),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_430),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_430),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_494),
.B(n_255),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_431),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_480),
.B(n_285),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_431),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_433),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_478),
.B(n_207),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_433),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_436),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_436),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_472),
.B(n_230),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_437),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_437),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_442),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_480),
.B(n_295),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_412),
.B(n_379),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_442),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_443),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_443),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g579 ( 
.A(n_450),
.B(n_263),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_445),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_445),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_446),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_446),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_449),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_503),
.B(n_293),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_449),
.Y(n_586)
);

NAND2x1p5_ASAP7_75t_L g587 ( 
.A(n_483),
.B(n_258),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_503),
.Y(n_588)
);

NAND2x1p5_ASAP7_75t_L g589 ( 
.A(n_483),
.B(n_258),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_427),
.B(n_379),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_484),
.Y(n_591)
);

OA21x2_ASAP7_75t_L g592 ( 
.A1(n_484),
.A2(n_317),
.B(n_315),
.Y(n_592)
);

AND3x2_ASAP7_75t_L g593 ( 
.A(n_462),
.B(n_352),
.C(n_337),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_485),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_485),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_486),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_486),
.Y(n_597)
);

INVx5_ASAP7_75t_L g598 ( 
.A(n_500),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_496),
.B(n_286),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_528),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_541),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_521),
.Y(n_602)
);

AND2x6_ASAP7_75t_L g603 ( 
.A(n_522),
.B(n_352),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_541),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_550),
.B(n_495),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_541),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_536),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_544),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_543),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_521),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_528),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_545),
.B(n_493),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_590),
.A2(n_487),
.B1(n_492),
.B2(n_302),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_528),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_588),
.Y(n_615)
);

INVx8_ASAP7_75t_L g616 ( 
.A(n_590),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_544),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_544),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_536),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_519),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_546),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_585),
.B(n_482),
.Y(n_622)
);

AO21x2_ASAP7_75t_L g623 ( 
.A1(n_546),
.A2(n_432),
.B(n_326),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_521),
.Y(n_624)
);

AO21x2_ASAP7_75t_L g625 ( 
.A1(n_546),
.A2(n_332),
.B(n_325),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_549),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_536),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_566),
.B(n_499),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_549),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_549),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_554),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_536),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_524),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_590),
.B(n_507),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_554),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_519),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_524),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_528),
.B(n_501),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_528),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_536),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_536),
.Y(n_641)
);

AND2x6_ASAP7_75t_L g642 ( 
.A(n_522),
.B(n_376),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_542),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_542),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_542),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_542),
.Y(n_646)
);

NAND3xp33_ASAP7_75t_L g647 ( 
.A(n_531),
.B(n_497),
.C(n_496),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_570),
.B(n_504),
.Y(n_648)
);

AND2x6_ASAP7_75t_L g649 ( 
.A(n_522),
.B(n_376),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_590),
.A2(n_561),
.B1(n_599),
.B2(n_592),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_527),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_590),
.A2(n_491),
.B1(n_319),
.B2(n_321),
.Y(n_652)
);

BUFx4f_ASAP7_75t_L g653 ( 
.A(n_592),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g654 ( 
.A(n_529),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_542),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_527),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_557),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_529),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_561),
.A2(n_330),
.B1(n_340),
.B2(n_291),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_542),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_588),
.B(n_474),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_557),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_551),
.Y(n_663)
);

AO22x2_ASAP7_75t_L g664 ( 
.A1(n_585),
.A2(n_471),
.B1(n_489),
.B2(n_497),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_561),
.A2(n_361),
.B1(n_366),
.B2(n_342),
.Y(n_665)
);

OAI22xp33_ASAP7_75t_SL g666 ( 
.A1(n_579),
.A2(n_476),
.B1(n_460),
.B2(n_224),
.Y(n_666)
);

OAI22xp33_ASAP7_75t_L g667 ( 
.A1(n_585),
.A2(n_514),
.B1(n_515),
.B2(n_513),
.Y(n_667)
);

BUFx10_ASAP7_75t_L g668 ( 
.A(n_575),
.Y(n_668)
);

BUFx10_ASAP7_75t_L g669 ( 
.A(n_575),
.Y(n_669)
);

AOI21x1_ASAP7_75t_L g670 ( 
.A1(n_531),
.A2(n_509),
.B(n_498),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_542),
.Y(n_671)
);

BUFx10_ASAP7_75t_L g672 ( 
.A(n_517),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_560),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_548),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_527),
.B(n_516),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_517),
.B(n_420),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_560),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_570),
.B(n_505),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_548),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_562),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_548),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_570),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_579),
.B(n_423),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_548),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_548),
.Y(n_685)
);

BUFx4f_ASAP7_75t_L g686 ( 
.A(n_592),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_562),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_548),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_599),
.B(n_453),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_548),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_561),
.A2(n_380),
.B1(n_382),
.B2(n_374),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_564),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_519),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_552),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_561),
.A2(n_392),
.B1(n_395),
.B2(n_386),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_L g696 ( 
.A(n_598),
.B(n_210),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_587),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_587),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_552),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_564),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_568),
.Y(n_701)
);

BUFx10_ASAP7_75t_L g702 ( 
.A(n_593),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_552),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_568),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_599),
.B(n_455),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_559),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_519),
.B(n_498),
.Y(n_707)
);

OR2x6_ASAP7_75t_L g708 ( 
.A(n_587),
.B(n_488),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_556),
.B(n_508),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_SL g710 ( 
.A(n_587),
.B(n_511),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_559),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_559),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_598),
.B(n_425),
.Y(n_713)
);

AND2x6_ASAP7_75t_L g714 ( 
.A(n_599),
.B(n_408),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_565),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_532),
.B(n_533),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_572),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_572),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_599),
.B(n_434),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_532),
.B(n_509),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_573),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_525),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_589),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_533),
.B(n_439),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_535),
.B(n_512),
.C(n_510),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_589),
.Y(n_726)
);

OAI22xp33_ASAP7_75t_L g727 ( 
.A1(n_589),
.A2(n_220),
.B1(n_377),
.B2(n_367),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_592),
.A2(n_401),
.B1(n_402),
.B2(n_403),
.Y(n_728)
);

BUFx6f_ASAP7_75t_SL g729 ( 
.A(n_594),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_565),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_565),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_567),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_573),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_576),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_535),
.Y(n_735)
);

OAI22xp33_ASAP7_75t_SL g736 ( 
.A1(n_589),
.A2(n_362),
.B1(n_237),
.B2(n_236),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_567),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_576),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_567),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_525),
.Y(n_740)
);

INVx4_ASAP7_75t_L g741 ( 
.A(n_539),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_593),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_582),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_571),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_582),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_571),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_583),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_571),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_583),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_538),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_538),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_735),
.Y(n_752)
);

NOR2xp67_ASAP7_75t_L g753 ( 
.A(n_609),
.B(n_452),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_682),
.B(n_598),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_735),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_682),
.B(n_598),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_602),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_616),
.B(n_668),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_616),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_609),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_616),
.B(n_668),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_R g762 ( 
.A(n_663),
.B(n_456),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_651),
.B(n_598),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_648),
.B(n_435),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_600),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_651),
.B(n_547),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_656),
.B(n_598),
.Y(n_767)
);

NOR3xp33_ASAP7_75t_L g768 ( 
.A(n_654),
.B(n_398),
.C(n_397),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_631),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_656),
.B(n_547),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_616),
.B(n_598),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_603),
.A2(n_596),
.B1(n_597),
.B2(n_594),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_648),
.B(n_440),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_603),
.B(n_534),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_668),
.B(n_525),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_622),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_675),
.B(n_553),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_668),
.B(n_525),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_669),
.B(n_553),
.Y(n_779)
);

NOR3xp33_ASAP7_75t_L g780 ( 
.A(n_667),
.B(n_224),
.C(n_220),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_603),
.B(n_558),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_669),
.B(n_634),
.Y(n_782)
);

NOR3xp33_ASAP7_75t_L g783 ( 
.A(n_633),
.B(n_236),
.C(n_229),
.Y(n_783)
);

NAND3xp33_ASAP7_75t_L g784 ( 
.A(n_724),
.B(n_237),
.C(n_229),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_615),
.B(n_444),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_669),
.B(n_558),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_635),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_635),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_603),
.B(n_596),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_669),
.B(n_525),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_603),
.B(n_597),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_637),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_603),
.B(n_591),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_658),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_657),
.Y(n_795)
);

OAI22xp33_ASAP7_75t_L g796 ( 
.A1(n_613),
.A2(n_563),
.B1(n_574),
.B2(n_409),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_603),
.B(n_591),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_672),
.B(n_563),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_642),
.B(n_591),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_642),
.B(n_574),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_610),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_642),
.B(n_525),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_642),
.A2(n_363),
.B1(n_250),
.B2(n_210),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_642),
.B(n_525),
.Y(n_804)
);

NOR3xp33_ASAP7_75t_L g805 ( 
.A(n_615),
.B(n_612),
.C(n_661),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_610),
.Y(n_806)
);

AO22x2_ASAP7_75t_L g807 ( 
.A1(n_683),
.A2(n_512),
.B1(n_510),
.B2(n_447),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_662),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_672),
.B(n_595),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_622),
.B(n_451),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_642),
.A2(n_649),
.B1(n_613),
.B2(n_714),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_600),
.Y(n_812)
);

INVx4_ASAP7_75t_L g813 ( 
.A(n_729),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_672),
.B(n_620),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_662),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_719),
.Y(n_816)
);

O2A1O1Ixp5_ASAP7_75t_L g817 ( 
.A1(n_632),
.A2(n_523),
.B(n_518),
.C(n_520),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_673),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_673),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_719),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_624),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_642),
.B(n_595),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_672),
.B(n_595),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_L g824 ( 
.A(n_714),
.B(n_750),
.Y(n_824)
);

NAND2xp33_ASAP7_75t_L g825 ( 
.A(n_714),
.B(n_214),
.Y(n_825)
);

OR2x2_ASAP7_75t_L g826 ( 
.A(n_678),
.B(n_454),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_649),
.B(n_595),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_626),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_677),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_677),
.Y(n_830)
);

OR2x6_ASAP7_75t_L g831 ( 
.A(n_742),
.B(n_457),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_650),
.A2(n_362),
.B1(n_240),
.B2(n_243),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_680),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_649),
.B(n_595),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_680),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_649),
.B(n_595),
.Y(n_836)
);

OR2x6_ASAP7_75t_L g837 ( 
.A(n_742),
.B(n_457),
.Y(n_837)
);

CKINVDCx16_ASAP7_75t_R g838 ( 
.A(n_709),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_687),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_649),
.B(n_518),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_649),
.B(n_638),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_714),
.A2(n_363),
.B1(n_244),
.B2(n_411),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_705),
.B(n_520),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_SL g844 ( 
.A1(n_710),
.A2(n_458),
.B1(n_464),
.B2(n_479),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_687),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_692),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_692),
.Y(n_847)
);

INVxp67_ASAP7_75t_R g848 ( 
.A(n_689),
.Y(n_848)
);

NOR3xp33_ASAP7_75t_L g849 ( 
.A(n_605),
.B(n_243),
.C(n_240),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_705),
.B(n_523),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_705),
.B(n_689),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_694),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_700),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_614),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_700),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_705),
.B(n_526),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_694),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_701),
.Y(n_858)
);

BUFx6f_ASAP7_75t_SL g859 ( 
.A(n_702),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_620),
.B(n_214),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_676),
.B(n_663),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_699),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_664),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_751),
.B(n_530),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_751),
.B(n_530),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_628),
.B(n_313),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_620),
.B(n_215),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_729),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_652),
.B(n_539),
.Y(n_869)
);

NAND2x1p5_ASAP7_75t_L g870 ( 
.A(n_697),
.B(n_592),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_697),
.B(n_539),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_699),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_698),
.B(n_539),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_653),
.A2(n_248),
.B(n_367),
.C(n_373),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_620),
.B(n_215),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_703),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_727),
.B(n_636),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_698),
.B(n_539),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_714),
.A2(n_378),
.B1(n_250),
.B2(n_244),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_723),
.B(n_235),
.Y(n_880)
);

INVxp67_ASAP7_75t_L g881 ( 
.A(n_664),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_723),
.B(n_264),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_636),
.B(n_219),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_702),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_701),
.Y(n_885)
);

OAI22xp33_ASAP7_75t_L g886 ( 
.A1(n_708),
.A2(n_248),
.B1(n_249),
.B2(n_251),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_636),
.B(n_316),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_726),
.B(n_394),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_726),
.B(n_219),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_706),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_664),
.Y(n_891)
);

INVx8_ASAP7_75t_L g892 ( 
.A(n_714),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_614),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_636),
.B(n_223),
.Y(n_894)
);

NOR3xp33_ASAP7_75t_L g895 ( 
.A(n_736),
.B(n_251),
.C(n_249),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_714),
.A2(n_242),
.B1(n_233),
.B2(n_226),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_693),
.B(n_223),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_693),
.B(n_226),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_653),
.A2(n_381),
.B(n_373),
.C(n_377),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_707),
.B(n_233),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_601),
.B(n_242),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_601),
.B(n_357),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_706),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_693),
.B(n_318),
.Y(n_904)
);

INVxp67_ASAP7_75t_SL g905 ( 
.A(n_740),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_604),
.B(n_357),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_604),
.B(n_606),
.Y(n_907)
);

OR2x2_ASAP7_75t_L g908 ( 
.A(n_659),
.B(n_481),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_702),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_711),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_611),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_664),
.B(n_490),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_702),
.B(n_459),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_R g914 ( 
.A(n_729),
.B(n_670),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_769),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_777),
.B(n_708),
.Y(n_916)
);

O2A1O1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_777),
.A2(n_736),
.B(n_716),
.C(n_720),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_798),
.B(n_666),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_817),
.A2(n_686),
.B(n_653),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_798),
.B(n_666),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_779),
.B(n_708),
.Y(n_921)
);

OR2x6_ASAP7_75t_L g922 ( 
.A(n_831),
.B(n_708),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_775),
.A2(n_693),
.B(n_722),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_796),
.A2(n_717),
.B(n_718),
.C(n_704),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_779),
.B(n_708),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_786),
.B(n_665),
.Y(n_926)
);

NOR2x1_ASAP7_75t_L g927 ( 
.A(n_813),
.B(n_713),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_765),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_786),
.B(n_691),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_776),
.B(n_695),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_877),
.A2(n_686),
.B(n_608),
.C(n_617),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_778),
.A2(n_722),
.B(n_641),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_782),
.B(n_741),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_907),
.A2(n_686),
.B(n_741),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_759),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_790),
.A2(n_641),
.B(n_632),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_782),
.B(n_741),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_796),
.A2(n_717),
.B(n_718),
.C(n_704),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_757),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_794),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_790),
.A2(n_645),
.B(n_643),
.Y(n_941)
);

AND2x6_ASAP7_75t_L g942 ( 
.A(n_811),
.B(n_606),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_759),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_823),
.A2(n_645),
.B(n_643),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_760),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_823),
.A2(n_660),
.B(n_646),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_766),
.B(n_728),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_851),
.B(n_741),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_787),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_788),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_757),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_877),
.B(n_740),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_813),
.B(n_611),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_766),
.A2(n_630),
.B(n_629),
.C(n_621),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_816),
.B(n_607),
.Y(n_955)
);

CKINVDCx6p67_ASAP7_75t_R g956 ( 
.A(n_792),
.Y(n_956)
);

NAND3xp33_ASAP7_75t_L g957 ( 
.A(n_805),
.B(n_725),
.C(n_647),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_809),
.A2(n_660),
.B(n_646),
.Y(n_958)
);

NAND2xp33_ASAP7_75t_L g959 ( 
.A(n_892),
.B(n_607),
.Y(n_959)
);

INVx2_ASAP7_75t_SL g960 ( 
.A(n_785),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_770),
.A2(n_617),
.B(n_608),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_820),
.B(n_607),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_848),
.A2(n_749),
.B1(n_721),
.B2(n_747),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_795),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_814),
.A2(n_674),
.B(n_671),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_886),
.B(n_740),
.Y(n_966)
);

AO21x1_ASAP7_75t_L g967 ( 
.A1(n_841),
.A2(n_621),
.B(n_618),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_770),
.A2(n_749),
.B1(n_721),
.B2(n_747),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_871),
.A2(n_629),
.B(n_618),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_913),
.B(n_630),
.Y(n_970)
);

NAND2x1_ASAP7_75t_L g971 ( 
.A(n_852),
.B(n_607),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_886),
.A2(n_733),
.B1(n_745),
.B2(n_734),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_831),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_763),
.A2(n_767),
.B(n_905),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_772),
.B(n_740),
.Y(n_975)
);

AOI21x1_ASAP7_75t_L g976 ( 
.A1(n_873),
.A2(n_734),
.B(n_733),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_887),
.B(n_623),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_887),
.B(n_623),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_SL g979 ( 
.A(n_753),
.B(n_647),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_808),
.Y(n_980)
);

AOI21x1_ASAP7_75t_L g981 ( 
.A1(n_878),
.A2(n_743),
.B(n_738),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_815),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_874),
.A2(n_738),
.B(n_743),
.C(n_745),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_838),
.B(n_619),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_874),
.A2(n_899),
.B(n_832),
.C(n_819),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_904),
.A2(n_623),
.B1(n_619),
.B2(n_644),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_904),
.B(n_625),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_754),
.A2(n_674),
.B(n_671),
.Y(n_988)
);

OAI21xp33_ASAP7_75t_L g989 ( 
.A1(n_899),
.A2(n_381),
.B(n_253),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_884),
.B(n_625),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_909),
.B(n_625),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_818),
.A2(n_655),
.B(n_640),
.C(n_681),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_756),
.A2(n_684),
.B(n_679),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_764),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_829),
.B(n_748),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_830),
.A2(n_655),
.B(n_640),
.C(n_681),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_833),
.B(n_748),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_835),
.B(n_711),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_758),
.B(n_740),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_831),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_839),
.B(n_712),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_810),
.B(n_459),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_845),
.A2(n_655),
.B1(n_619),
.B2(n_627),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_846),
.B(n_746),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_800),
.A2(n_684),
.B(n_679),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_821),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_847),
.B(n_746),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_773),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_758),
.B(n_619),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_853),
.B(n_744),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_837),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_860),
.A2(n_690),
.B(n_688),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_855),
.A2(n_885),
.B1(n_858),
.B2(n_843),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_789),
.A2(n_791),
.B(n_802),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_860),
.A2(n_690),
.B(n_688),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_867),
.A2(n_640),
.B(n_627),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_867),
.A2(n_640),
.B(n_627),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_761),
.B(n_627),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_837),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_804),
.A2(n_655),
.B(n_644),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_780),
.A2(n_644),
.B1(n_681),
.B2(n_685),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_875),
.A2(n_681),
.B(n_644),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_762),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_761),
.B(n_685),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_837),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_850),
.A2(n_685),
.B(n_696),
.Y(n_1026)
);

AOI21x1_ASAP7_75t_L g1027 ( 
.A1(n_822),
.A2(n_670),
.B(n_712),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_875),
.A2(n_685),
.B(n_639),
.Y(n_1028)
);

NOR3xp33_ASAP7_75t_L g1029 ( 
.A(n_784),
.B(n_725),
.C(n_341),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_880),
.B(n_715),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_866),
.A2(n_744),
.B(n_739),
.C(n_737),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_856),
.A2(n_739),
.B(n_730),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_882),
.B(n_715),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_888),
.B(n_737),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_864),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_883),
.A2(n_639),
.B(n_730),
.Y(n_1036)
);

AOI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_891),
.A2(n_732),
.B1(n_731),
.B2(n_555),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_866),
.A2(n_732),
.B(n_731),
.C(n_368),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_865),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_SL g1040 ( 
.A1(n_883),
.A2(n_356),
.B(n_355),
.C(n_354),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_826),
.B(n_463),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_SL g1042 ( 
.A1(n_894),
.A2(n_334),
.B(n_404),
.C(n_408),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_752),
.B(n_253),
.Y(n_1043)
);

AOI21xp33_ASAP7_75t_L g1044 ( 
.A1(n_774),
.A2(n_390),
.B(n_383),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_762),
.B(n_463),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_854),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_914),
.B(n_803),
.Y(n_1047)
);

AO21x1_ASAP7_75t_L g1048 ( 
.A1(n_870),
.A2(n_578),
.B(n_577),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_755),
.B(n_383),
.Y(n_1049)
);

INVx1_ASAP7_75t_SL g1050 ( 
.A(n_844),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_781),
.B(n_390),
.Y(n_1051)
);

NAND2x1p5_ASAP7_75t_L g1052 ( 
.A(n_868),
.B(n_854),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_868),
.B(n_364),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_863),
.B(n_396),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_765),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_869),
.A2(n_881),
.B1(n_895),
.B2(n_912),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_889),
.B(n_396),
.Y(n_1057)
);

NOR3xp33_ASAP7_75t_L g1058 ( 
.A(n_849),
.B(n_322),
.C(n_351),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_897),
.A2(n_555),
.B(n_364),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_861),
.Y(n_1060)
);

NOR3xp33_ASAP7_75t_L g1061 ( 
.A(n_783),
.B(n_350),
.C(n_349),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_765),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_900),
.B(n_400),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_914),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_901),
.B(n_400),
.Y(n_1065)
);

AO21x1_ASAP7_75t_L g1066 ( 
.A1(n_870),
.A2(n_577),
.B(n_584),
.Y(n_1066)
);

OAI21xp33_ASAP7_75t_L g1067 ( 
.A1(n_902),
.A2(n_409),
.B(n_406),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_890),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_897),
.A2(n_555),
.B(n_370),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_908),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_911),
.B(n_467),
.Y(n_1071)
);

NOR2xp67_ASAP7_75t_L g1072 ( 
.A(n_906),
.B(n_467),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_807),
.B(n_406),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_898),
.A2(n_555),
.B(n_372),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_807),
.B(n_345),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_898),
.A2(n_371),
.B(n_372),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_771),
.A2(n_371),
.B(n_375),
.Y(n_1077)
);

OAI21xp33_ASAP7_75t_SL g1078 ( 
.A1(n_842),
.A2(n_469),
.B(n_473),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_892),
.A2(n_348),
.B1(n_209),
.B2(n_375),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_824),
.A2(n_799),
.B(n_797),
.C(n_793),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_827),
.A2(n_584),
.B(n_581),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_903),
.A2(n_378),
.B(n_387),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_768),
.A2(n_577),
.B(n_581),
.C(n_580),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_859),
.B(n_399),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_903),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_825),
.A2(n_399),
.B(n_405),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_879),
.A2(n_578),
.B(n_581),
.C(n_580),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_892),
.A2(n_405),
.B1(n_407),
.B2(n_411),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_896),
.A2(n_407),
.B1(n_320),
.B2(n_259),
.Y(n_1089)
);

O2A1O1Ixp5_ASAP7_75t_L g1090 ( 
.A1(n_840),
.A2(n_580),
.B(n_540),
.C(n_477),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_834),
.A2(n_308),
.B(n_266),
.Y(n_1091)
);

AOI21x1_ASAP7_75t_L g1092 ( 
.A1(n_987),
.A2(n_836),
.B(n_910),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_994),
.B(n_469),
.Y(n_1093)
);

O2A1O1Ixp5_ASAP7_75t_L g1094 ( 
.A1(n_1048),
.A2(n_857),
.B(n_828),
.C(n_876),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_1023),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_R g1096 ( 
.A(n_945),
.B(n_859),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_939),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_916),
.A2(n_911),
.B1(n_893),
.B2(n_812),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_922),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1002),
.B(n_473),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_951),
.Y(n_1101)
);

INVx2_ASAP7_75t_SL g1102 ( 
.A(n_956),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_922),
.B(n_765),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1027),
.A2(n_872),
.B(n_862),
.Y(n_1104)
);

INVxp67_ASAP7_75t_L g1105 ( 
.A(n_940),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_1008),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_915),
.Y(n_1107)
);

NOR2xp67_ASAP7_75t_L g1108 ( 
.A(n_984),
.B(n_812),
.Y(n_1108)
);

INVxp67_ASAP7_75t_SL g1109 ( 
.A(n_921),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1035),
.B(n_1039),
.Y(n_1110)
);

OAI21xp33_ASAP7_75t_SL g1111 ( 
.A1(n_925),
.A2(n_801),
.B(n_806),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_926),
.B(n_929),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1050),
.A2(n_893),
.B1(n_812),
.B2(n_477),
.Y(n_1113)
);

AO32x2_ASAP7_75t_L g1114 ( 
.A1(n_968),
.A2(n_540),
.A3(n_586),
.B1(n_569),
.B2(n_893),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_918),
.B(n_812),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_R g1116 ( 
.A(n_960),
.B(n_893),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_SL g1117 ( 
.A1(n_1070),
.A2(n_305),
.B1(n_270),
.B2(n_273),
.Y(n_1117)
);

AND2x6_ASAP7_75t_L g1118 ( 
.A(n_963),
.B(n_218),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_972),
.A2(n_586),
.B1(n_569),
.B2(n_540),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_977),
.A2(n_311),
.B(n_274),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_918),
.B(n_2),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1006),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_SL g1123 ( 
.A1(n_1058),
.A2(n_962),
.B(n_955),
.C(n_983),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_SL g1124 ( 
.A1(n_1058),
.A2(n_3),
.B(n_7),
.C(n_8),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_984),
.B(n_281),
.Y(n_1125)
);

NOR3xp33_ASAP7_75t_L g1126 ( 
.A(n_920),
.B(n_287),
.C(n_288),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_947),
.A2(n_586),
.B1(n_569),
.B2(n_347),
.Y(n_1127)
);

OR2x2_ASAP7_75t_L g1128 ( 
.A(n_1041),
.B(n_569),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_979),
.B(n_290),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_920),
.A2(n_9),
.B(n_11),
.C(n_12),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_SL g1131 ( 
.A1(n_955),
.A2(n_9),
.B(n_12),
.C(n_13),
.Y(n_1131)
);

NOR2xp67_ASAP7_75t_L g1132 ( 
.A(n_1064),
.B(n_292),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_928),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_931),
.A2(n_323),
.B(n_298),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1045),
.B(n_14),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_930),
.B(n_15),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_978),
.A2(n_327),
.B(n_297),
.Y(n_1137)
);

INVxp67_ASAP7_75t_L g1138 ( 
.A(n_1060),
.Y(n_1138)
);

NAND2x1p5_ASAP7_75t_L g1139 ( 
.A(n_1046),
.B(n_569),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_933),
.B(n_299),
.Y(n_1140)
);

INVxp67_ASAP7_75t_SL g1141 ( 
.A(n_1064),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_SL g1142 ( 
.A(n_922),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1071),
.B(n_20),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_973),
.B(n_304),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1013),
.A2(n_586),
.B1(n_569),
.B2(n_339),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_1075),
.A2(n_586),
.B1(n_329),
.B2(n_335),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1071),
.B(n_949),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_973),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1000),
.B(n_1019),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_1000),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_950),
.B(n_22),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_964),
.A2(n_586),
.B1(n_312),
.B2(n_307),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_928),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_1011),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_934),
.A2(n_218),
.B(n_537),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1019),
.B(n_24),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_933),
.A2(n_218),
.B(n_537),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_980),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_1025),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_937),
.A2(n_974),
.B(n_919),
.Y(n_1160)
);

AND2x6_ASAP7_75t_L g1161 ( 
.A(n_928),
.B(n_218),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_937),
.A2(n_537),
.B(n_185),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_982),
.B(n_25),
.Y(n_1163)
);

NAND3xp33_ASAP7_75t_L g1164 ( 
.A(n_1029),
.B(n_537),
.C(n_28),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_959),
.A2(n_537),
.B(n_182),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1025),
.B(n_27),
.Y(n_1166)
);

OR2x6_ASAP7_75t_L g1167 ( 
.A(n_1052),
.B(n_28),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_R g1168 ( 
.A(n_1084),
.B(n_178),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_948),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1085),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_961),
.A2(n_537),
.B(n_173),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_1052),
.Y(n_1172)
);

AND2x2_ASAP7_75t_SL g1173 ( 
.A(n_1056),
.B(n_31),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_SL g1174 ( 
.A(n_1061),
.B(n_33),
.C(n_34),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1063),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1061),
.B(n_37),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_928),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_988),
.A2(n_170),
.B(n_159),
.Y(n_1178)
);

BUFx8_ASAP7_75t_L g1179 ( 
.A(n_953),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_993),
.A2(n_156),
.B(n_146),
.Y(n_1180)
);

INVxp67_ASAP7_75t_L g1181 ( 
.A(n_1084),
.Y(n_1181)
);

AO21x1_ASAP7_75t_L g1182 ( 
.A1(n_952),
.A2(n_145),
.B(n_127),
.Y(n_1182)
);

INVxp67_ASAP7_75t_L g1183 ( 
.A(n_1054),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_948),
.B(n_42),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_958),
.A2(n_124),
.B(n_118),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_962),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_970),
.B(n_43),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_942),
.B(n_45),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1046),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_953),
.B(n_46),
.Y(n_1190)
);

OR2x2_ASAP7_75t_L g1191 ( 
.A(n_1065),
.B(n_47),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1056),
.B(n_52),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1057),
.A2(n_53),
.B(n_55),
.C(n_59),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1062),
.B(n_61),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_924),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1067),
.B(n_66),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1062),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_942),
.B(n_67),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1055),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_917),
.A2(n_67),
.B(n_70),
.C(n_71),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1055),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_938),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_965),
.A2(n_89),
.B(n_103),
.Y(n_1203)
);

BUFx12f_ASAP7_75t_L g1204 ( 
.A(n_1055),
.Y(n_1204)
);

INVx1_ASAP7_75t_SL g1205 ( 
.A(n_942),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_957),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_942),
.B(n_76),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_1043),
.B(n_80),
.Y(n_1208)
);

AO32x1_ASAP7_75t_L g1209 ( 
.A1(n_1003),
.A2(n_91),
.A3(n_98),
.B1(n_100),
.B2(n_104),
.Y(n_1209)
);

A2O1A1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_985),
.A2(n_1044),
.B(n_989),
.C(n_1029),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_995),
.A2(n_997),
.B1(n_1001),
.B2(n_1004),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_999),
.A2(n_941),
.B(n_936),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_942),
.B(n_952),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_932),
.A2(n_923),
.B(n_944),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1055),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_946),
.A2(n_1018),
.B(n_1009),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1009),
.A2(n_1018),
.B(n_1024),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1024),
.A2(n_1026),
.B(n_1015),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1088),
.B(n_935),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1068),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_SL g1221 ( 
.A1(n_1073),
.A2(n_1079),
.B1(n_1049),
.B2(n_1051),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_954),
.A2(n_992),
.B(n_996),
.C(n_1053),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1090),
.A2(n_986),
.B(n_1069),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1047),
.B(n_1089),
.Y(n_1224)
);

OR2x6_ASAP7_75t_L g1225 ( 
.A(n_1047),
.B(n_927),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_966),
.B(n_1033),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_943),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1030),
.B(n_1034),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1072),
.B(n_1007),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_R g1230 ( 
.A(n_943),
.B(n_981),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1021),
.B(n_1076),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_990),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_998),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1012),
.A2(n_969),
.B(n_1016),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_971),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1078),
.B(n_991),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1010),
.B(n_1086),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_976),
.A2(n_1005),
.B(n_1066),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1038),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1083),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1017),
.A2(n_1022),
.B(n_1080),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_975),
.A2(n_1028),
.B(n_1036),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1037),
.B(n_1032),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1181),
.B(n_1040),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1105),
.B(n_1141),
.Y(n_1245)
);

INVx4_ASAP7_75t_L g1246 ( 
.A(n_1204),
.Y(n_1246)
);

OAI22x1_ASAP7_75t_L g1247 ( 
.A1(n_1192),
.A2(n_1224),
.B1(n_1121),
.B2(n_1190),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1103),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1160),
.A2(n_975),
.B(n_1020),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1110),
.B(n_1082),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1093),
.B(n_1037),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1107),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1210),
.A2(n_1090),
.B(n_1031),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1110),
.B(n_1042),
.Y(n_1254)
);

BUFx2_ASAP7_75t_R g1255 ( 
.A(n_1095),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1103),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1112),
.B(n_1014),
.Y(n_1257)
);

AO31x2_ASAP7_75t_L g1258 ( 
.A1(n_1211),
.A2(n_1059),
.A3(n_1074),
.B(n_1087),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1211),
.A2(n_1214),
.B(n_1171),
.Y(n_1259)
);

NAND3xp33_ASAP7_75t_L g1260 ( 
.A(n_1195),
.B(n_1077),
.C(n_1091),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_SL g1261 ( 
.A(n_1173),
.B(n_1081),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1099),
.B(n_1172),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1100),
.B(n_1159),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1162),
.A2(n_1234),
.B(n_1241),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1116),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1109),
.B(n_1233),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1096),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1158),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1190),
.B(n_1149),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1126),
.A2(n_1196),
.B1(n_1115),
.B2(n_1118),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1148),
.B(n_1150),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1133),
.Y(n_1272)
);

BUFx12f_ASAP7_75t_L g1273 ( 
.A(n_1102),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1232),
.B(n_1147),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1242),
.A2(n_1218),
.B(n_1238),
.Y(n_1275)
);

AO31x2_ASAP7_75t_L g1276 ( 
.A1(n_1243),
.A2(n_1127),
.A3(n_1182),
.B(n_1216),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1205),
.B(n_1108),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1237),
.A2(n_1184),
.B(n_1165),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1094),
.A2(n_1092),
.B(n_1223),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1184),
.A2(n_1140),
.B(n_1223),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_SL g1281 ( 
.A(n_1118),
.B(n_1205),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1231),
.A2(n_1145),
.B(n_1098),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1240),
.A2(n_1217),
.B(n_1222),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1187),
.A2(n_1226),
.B(n_1188),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1155),
.A2(n_1203),
.B(n_1178),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1187),
.A2(n_1188),
.B(n_1198),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1106),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1118),
.A2(n_1239),
.B1(n_1183),
.B2(n_1174),
.Y(n_1288)
);

A2O1A1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1130),
.A2(n_1135),
.B(n_1208),
.C(n_1164),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1198),
.A2(n_1119),
.B(n_1127),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1145),
.A2(n_1098),
.B(n_1123),
.Y(n_1291)
);

NAND2x1_ASAP7_75t_L g1292 ( 
.A(n_1177),
.B(n_1199),
.Y(n_1292)
);

AOI221x1_ASAP7_75t_L g1293 ( 
.A1(n_1195),
.A2(n_1202),
.B1(n_1206),
.B2(n_1169),
.C(n_1200),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1133),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1136),
.B(n_1154),
.Y(n_1295)
);

BUFx12f_ASAP7_75t_L g1296 ( 
.A(n_1179),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1180),
.A2(n_1185),
.B(n_1207),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1209),
.A2(n_1228),
.B(n_1157),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1220),
.Y(n_1299)
);

INVx3_ASAP7_75t_SL g1300 ( 
.A(n_1167),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_SL g1301 ( 
.A1(n_1219),
.A2(n_1124),
.B(n_1169),
.C(n_1202),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1207),
.A2(n_1119),
.B(n_1213),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1156),
.B(n_1166),
.Y(n_1303)
);

AO21x1_ASAP7_75t_L g1304 ( 
.A1(n_1134),
.A2(n_1206),
.B(n_1176),
.Y(n_1304)
);

AOI221xp5_ASAP7_75t_SL g1305 ( 
.A1(n_1175),
.A2(n_1193),
.B1(n_1163),
.B2(n_1151),
.C(n_1221),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1133),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1230),
.A2(n_1134),
.B(n_1137),
.Y(n_1307)
);

A2O1A1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1191),
.A2(n_1229),
.B(n_1120),
.C(n_1129),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1199),
.A2(n_1215),
.B(n_1139),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1118),
.A2(n_1097),
.B1(n_1170),
.B2(n_1101),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1111),
.A2(n_1186),
.B(n_1152),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1138),
.B(n_1144),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1209),
.A2(n_1125),
.B(n_1235),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1225),
.B(n_1122),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1179),
.A2(n_1167),
.B1(n_1117),
.B2(n_1143),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_1153),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1099),
.B(n_1189),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1152),
.A2(n_1128),
.B(n_1146),
.Y(n_1318)
);

AOI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1225),
.A2(n_1132),
.B(n_1167),
.Y(n_1319)
);

O2A1O1Ixp33_ASAP7_75t_SL g1320 ( 
.A1(n_1131),
.A2(n_1209),
.B(n_1227),
.C(n_1225),
.Y(n_1320)
);

NOR2xp67_ASAP7_75t_L g1321 ( 
.A(n_1153),
.B(n_1201),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1113),
.A2(n_1114),
.B(n_1161),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1153),
.B(n_1201),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1194),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1201),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1194),
.B(n_1197),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1114),
.A2(n_1161),
.B(n_1142),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1161),
.A2(n_1114),
.B(n_1168),
.Y(n_1328)
);

A2O1A1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1142),
.A2(n_1224),
.B(n_918),
.C(n_920),
.Y(n_1329)
);

AND2x2_ASAP7_75t_SL g1330 ( 
.A(n_1161),
.B(n_1173),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1160),
.A2(n_916),
.B(n_921),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1224),
.A2(n_918),
.B(n_920),
.C(n_777),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1104),
.A2(n_1212),
.B(n_1241),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1121),
.A2(n_916),
.B(n_931),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1160),
.A2(n_916),
.B(n_921),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1160),
.A2(n_916),
.B(n_921),
.Y(n_1336)
);

AO22x2_ASAP7_75t_L g1337 ( 
.A1(n_1192),
.A2(n_912),
.B1(n_1202),
.B2(n_1195),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_1204),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1096),
.Y(n_1339)
);

AO32x2_ASAP7_75t_L g1340 ( 
.A1(n_1195),
.A2(n_1202),
.A3(n_1206),
.B1(n_1169),
.B2(n_1211),
.Y(n_1340)
);

AOI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1224),
.A2(n_1173),
.B1(n_609),
.B2(n_637),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1093),
.B(n_764),
.Y(n_1342)
);

AO31x2_ASAP7_75t_L g1343 ( 
.A1(n_1236),
.A2(n_967),
.A3(n_1066),
.B(n_1048),
.Y(n_1343)
);

NAND3xp33_ASAP7_75t_L g1344 ( 
.A(n_1224),
.B(n_1202),
.C(n_1195),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_1095),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1173),
.A2(n_916),
.B1(n_1121),
.B2(n_877),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1160),
.A2(n_916),
.B(n_921),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1236),
.A2(n_967),
.A3(n_1066),
.B(n_1048),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1160),
.A2(n_916),
.B(n_921),
.Y(n_1349)
);

A2O1A1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1224),
.A2(n_918),
.B(n_920),
.C(n_777),
.Y(n_1350)
);

INVxp67_ASAP7_75t_L g1351 ( 
.A(n_1093),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1181),
.B(n_760),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1107),
.Y(n_1353)
);

CKINVDCx11_ASAP7_75t_R g1354 ( 
.A(n_1204),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1121),
.A2(n_916),
.B(n_931),
.Y(n_1355)
);

OA21x2_ASAP7_75t_L g1356 ( 
.A1(n_1160),
.A2(n_1238),
.B(n_1234),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1204),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1160),
.A2(n_916),
.B(n_921),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1160),
.A2(n_916),
.B(n_921),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1160),
.A2(n_916),
.B(n_921),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1096),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1104),
.A2(n_1212),
.B(n_1241),
.Y(n_1362)
);

AOI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1160),
.A2(n_1212),
.B(n_1241),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1160),
.A2(n_916),
.B(n_921),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1181),
.B(n_760),
.Y(n_1365)
);

O2A1O1Ixp33_ASAP7_75t_SL g1366 ( 
.A1(n_1123),
.A2(n_758),
.B(n_761),
.C(n_916),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1112),
.B(n_1110),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1104),
.A2(n_1212),
.B(n_1241),
.Y(n_1368)
);

AO31x2_ASAP7_75t_L g1369 ( 
.A1(n_1236),
.A2(n_967),
.A3(n_1066),
.B(n_1048),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1104),
.A2(n_1212),
.B(n_1241),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1096),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1173),
.A2(n_916),
.B1(n_1121),
.B2(n_877),
.Y(n_1372)
);

AO21x1_ASAP7_75t_L g1373 ( 
.A1(n_1224),
.A2(n_1121),
.B(n_1184),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1160),
.A2(n_916),
.B(n_921),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1104),
.A2(n_1212),
.B(n_1241),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1160),
.A2(n_1238),
.B(n_1234),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1181),
.B(n_760),
.Y(n_1377)
);

CKINVDCx16_ASAP7_75t_R g1378 ( 
.A(n_1096),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1159),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1181),
.B(n_760),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1093),
.B(n_764),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1096),
.Y(n_1382)
);

NOR2xp67_ASAP7_75t_L g1383 ( 
.A(n_1105),
.B(n_760),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1104),
.A2(n_1212),
.B(n_1241),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1107),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1095),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1121),
.A2(n_916),
.B(n_931),
.Y(n_1387)
);

AO32x2_ASAP7_75t_L g1388 ( 
.A1(n_1195),
.A2(n_1202),
.A3(n_1206),
.B1(n_1169),
.B2(n_1211),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1121),
.A2(n_916),
.B(n_931),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1107),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1093),
.B(n_776),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1104),
.A2(n_1212),
.B(n_1241),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1181),
.B(n_760),
.Y(n_1393)
);

INVx4_ASAP7_75t_L g1394 ( 
.A(n_1204),
.Y(n_1394)
);

OAI21xp33_ASAP7_75t_L g1395 ( 
.A1(n_1121),
.A2(n_777),
.B(n_609),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1093),
.B(n_776),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1160),
.A2(n_1238),
.B(n_1234),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1181),
.B(n_916),
.Y(n_1398)
);

INVxp67_ASAP7_75t_SL g1399 ( 
.A(n_1141),
.Y(n_1399)
);

CKINVDCx11_ASAP7_75t_R g1400 ( 
.A(n_1296),
.Y(n_1400)
);

NAND2x1p5_ASAP7_75t_L g1401 ( 
.A(n_1262),
.B(n_1265),
.Y(n_1401)
);

OAI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1341),
.A2(n_1274),
.B1(n_1315),
.B2(n_1270),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1337),
.A2(n_1344),
.B1(n_1330),
.B2(n_1372),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1252),
.Y(n_1404)
);

INVx6_ASAP7_75t_L g1405 ( 
.A(n_1378),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_SL g1406 ( 
.A1(n_1337),
.A2(n_1344),
.B1(n_1346),
.B2(n_1372),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1346),
.A2(n_1247),
.B1(n_1304),
.B2(n_1381),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_SL g1408 ( 
.A1(n_1300),
.A2(n_1352),
.B1(n_1365),
.B2(n_1377),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1332),
.A2(n_1350),
.B1(n_1303),
.B2(n_1395),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1261),
.A2(n_1281),
.B1(n_1290),
.B2(n_1328),
.Y(n_1410)
);

INVx6_ASAP7_75t_L g1411 ( 
.A(n_1338),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1268),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1342),
.A2(n_1251),
.B1(n_1373),
.B2(n_1261),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1353),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1288),
.A2(n_1284),
.B1(n_1351),
.B2(n_1290),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1329),
.A2(n_1289),
.B1(n_1399),
.B2(n_1282),
.Y(n_1416)
);

INVx6_ASAP7_75t_L g1417 ( 
.A(n_1338),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1284),
.A2(n_1286),
.B1(n_1355),
.B2(n_1334),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1294),
.Y(n_1419)
);

INVx6_ASAP7_75t_L g1420 ( 
.A(n_1338),
.Y(n_1420)
);

BUFx4f_ASAP7_75t_SL g1421 ( 
.A(n_1345),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1385),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1390),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1286),
.A2(n_1387),
.B1(n_1334),
.B2(n_1355),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_1256),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1387),
.A2(n_1389),
.B1(n_1244),
.B2(n_1328),
.Y(n_1426)
);

OAI21xp33_ASAP7_75t_L g1427 ( 
.A1(n_1280),
.A2(n_1291),
.B(n_1308),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_1267),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1389),
.A2(n_1396),
.B1(n_1391),
.B2(n_1281),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1339),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1398),
.A2(n_1318),
.B1(n_1367),
.B2(n_1266),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1379),
.B(n_1271),
.Y(n_1432)
);

AOI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1380),
.A2(n_1393),
.B1(n_1312),
.B2(n_1245),
.Y(n_1433)
);

OAI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1293),
.A2(n_1340),
.B1(n_1388),
.B2(n_1254),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1318),
.A2(n_1266),
.B1(n_1311),
.B2(n_1269),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1311),
.A2(n_1340),
.B1(n_1388),
.B2(n_1283),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1379),
.B(n_1314),
.Y(n_1437)
);

INVx6_ASAP7_75t_L g1438 ( 
.A(n_1357),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1354),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1314),
.B(n_1295),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1340),
.A2(n_1388),
.B1(n_1283),
.B2(n_1250),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1256),
.Y(n_1442)
);

CKINVDCx11_ASAP7_75t_R g1443 ( 
.A(n_1273),
.Y(n_1443)
);

INVx4_ASAP7_75t_L g1444 ( 
.A(n_1371),
.Y(n_1444)
);

CKINVDCx11_ASAP7_75t_R g1445 ( 
.A(n_1386),
.Y(n_1445)
);

CKINVDCx11_ASAP7_75t_R g1446 ( 
.A(n_1357),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1382),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1307),
.A2(n_1253),
.B1(n_1324),
.B2(n_1257),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1255),
.Y(n_1449)
);

INVx3_ASAP7_75t_L g1450 ( 
.A(n_1294),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1361),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1265),
.B(n_1287),
.Y(n_1452)
);

CKINVDCx20_ASAP7_75t_R g1453 ( 
.A(n_1357),
.Y(n_1453)
);

CKINVDCx11_ASAP7_75t_R g1454 ( 
.A(n_1246),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1323),
.Y(n_1455)
);

OAI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1326),
.A2(n_1253),
.B1(n_1360),
.B2(n_1331),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1248),
.B(n_1262),
.Y(n_1457)
);

CKINVDCx20_ASAP7_75t_R g1458 ( 
.A(n_1246),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_1306),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1394),
.B(n_1383),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1394),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1306),
.Y(n_1462)
);

BUFx4f_ASAP7_75t_SL g1463 ( 
.A(n_1316),
.Y(n_1463)
);

NAND2x1p5_ASAP7_75t_L g1464 ( 
.A(n_1277),
.B(n_1321),
.Y(n_1464)
);

AO22x1_ASAP7_75t_L g1465 ( 
.A1(n_1317),
.A2(n_1272),
.B1(n_1323),
.B2(n_1325),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1319),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1305),
.B(n_1335),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1260),
.A2(n_1259),
.B1(n_1374),
.B2(n_1364),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1305),
.B(n_1309),
.Y(n_1469)
);

CKINVDCx11_ASAP7_75t_R g1470 ( 
.A(n_1292),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1307),
.A2(n_1260),
.B1(n_1310),
.B2(n_1358),
.Y(n_1471)
);

INVx4_ASAP7_75t_L g1472 ( 
.A(n_1356),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1336),
.B(n_1359),
.Y(n_1473)
);

OR2x6_ASAP7_75t_L g1474 ( 
.A(n_1327),
.B(n_1322),
.Y(n_1474)
);

INVx8_ASAP7_75t_L g1475 ( 
.A(n_1301),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1343),
.B(n_1348),
.Y(n_1476)
);

CKINVDCx20_ASAP7_75t_R g1477 ( 
.A(n_1313),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1302),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1347),
.A2(n_1349),
.B1(n_1298),
.B2(n_1278),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1249),
.A2(n_1264),
.B1(n_1297),
.B2(n_1397),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1376),
.A2(n_1397),
.B1(n_1279),
.B2(n_1285),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1363),
.A2(n_1376),
.B1(n_1366),
.B2(n_1320),
.Y(n_1482)
);

BUFx10_ASAP7_75t_L g1483 ( 
.A(n_1348),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1275),
.A2(n_1368),
.B1(n_1384),
.B2(n_1375),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1333),
.A2(n_1362),
.B1(n_1370),
.B2(n_1392),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1276),
.A2(n_1337),
.B1(n_1173),
.B2(n_1344),
.Y(n_1486)
);

INVx6_ASAP7_75t_L g1487 ( 
.A(n_1369),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1258),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1258),
.Y(n_1489)
);

CKINVDCx6p67_ASAP7_75t_R g1490 ( 
.A(n_1276),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1338),
.Y(n_1491)
);

OAI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1344),
.A2(n_1341),
.B1(n_1293),
.B2(n_1261),
.Y(n_1492)
);

BUFx6f_ASAP7_75t_L g1493 ( 
.A(n_1256),
.Y(n_1493)
);

BUFx10_ASAP7_75t_L g1494 ( 
.A(n_1267),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1337),
.A2(n_1173),
.B1(n_1344),
.B2(n_1330),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1337),
.A2(n_1173),
.B1(n_1344),
.B2(n_1330),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1341),
.A2(n_1344),
.B1(n_1350),
.B2(n_1332),
.Y(n_1497)
);

BUFx3_ASAP7_75t_L g1498 ( 
.A(n_1296),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_SL g1499 ( 
.A1(n_1337),
.A2(n_1173),
.B1(n_1330),
.B2(n_1344),
.Y(n_1499)
);

BUFx12f_ASAP7_75t_L g1500 ( 
.A(n_1354),
.Y(n_1500)
);

INVx6_ASAP7_75t_L g1501 ( 
.A(n_1378),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1341),
.A2(n_1344),
.B1(n_1350),
.B2(n_1332),
.Y(n_1502)
);

INVx4_ASAP7_75t_L g1503 ( 
.A(n_1267),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1296),
.Y(n_1504)
);

BUFx8_ASAP7_75t_SL g1505 ( 
.A(n_1345),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1341),
.A2(n_1344),
.B1(n_1350),
.B2(n_1332),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1267),
.Y(n_1507)
);

CKINVDCx11_ASAP7_75t_R g1508 ( 
.A(n_1296),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_SL g1509 ( 
.A1(n_1337),
.A2(n_1173),
.B1(n_1330),
.B2(n_1344),
.Y(n_1509)
);

OAI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1344),
.A2(n_1341),
.B1(n_1293),
.B2(n_1261),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_SL g1511 ( 
.A1(n_1337),
.A2(n_1173),
.B1(n_1330),
.B2(n_1344),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1294),
.Y(n_1512)
);

OAI22x1_ASAP7_75t_L g1513 ( 
.A1(n_1341),
.A2(n_1300),
.B1(n_1315),
.B2(n_1344),
.Y(n_1513)
);

CKINVDCx11_ASAP7_75t_R g1514 ( 
.A(n_1296),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1299),
.Y(n_1515)
);

CKINVDCx20_ASAP7_75t_R g1516 ( 
.A(n_1378),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1337),
.A2(n_1173),
.B1(n_1344),
.B2(n_1330),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1296),
.Y(n_1518)
);

CKINVDCx9p33_ASAP7_75t_R g1519 ( 
.A(n_1245),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1341),
.A2(n_1344),
.B1(n_1350),
.B2(n_1332),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1337),
.A2(n_1173),
.B1(n_1344),
.B2(n_1330),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1337),
.A2(n_1173),
.B1(n_1344),
.B2(n_1330),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1341),
.A2(n_1344),
.B1(n_1350),
.B2(n_1332),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1299),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1341),
.A2(n_1344),
.B1(n_1350),
.B2(n_1332),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1263),
.B(n_1342),
.Y(n_1526)
);

OAI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1344),
.A2(n_1341),
.B1(n_1293),
.B2(n_1261),
.Y(n_1527)
);

BUFx12f_ASAP7_75t_L g1528 ( 
.A(n_1354),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1436),
.B(n_1406),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1476),
.B(n_1436),
.Y(n_1530)
);

AO31x2_ASAP7_75t_L g1531 ( 
.A1(n_1489),
.A2(n_1482),
.A3(n_1468),
.B(n_1488),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1480),
.A2(n_1479),
.B(n_1481),
.Y(n_1532)
);

OA21x2_ASAP7_75t_L g1533 ( 
.A1(n_1479),
.A2(n_1427),
.B(n_1480),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1404),
.Y(n_1534)
);

CKINVDCx12_ASAP7_75t_R g1535 ( 
.A(n_1408),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1437),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1487),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1487),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_SL g1539 ( 
.A(n_1402),
.B(n_1492),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1412),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1414),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1432),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1422),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1423),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1474),
.B(n_1466),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1406),
.A2(n_1521),
.B1(n_1522),
.B2(n_1517),
.Y(n_1546)
);

OAI221xp5_ASAP7_75t_L g1547 ( 
.A1(n_1499),
.A2(n_1511),
.B1(n_1509),
.B2(n_1426),
.C(n_1415),
.Y(n_1547)
);

OA21x2_ASAP7_75t_L g1548 ( 
.A1(n_1481),
.A2(n_1473),
.B(n_1471),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1474),
.B(n_1469),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1474),
.B(n_1457),
.Y(n_1550)
);

AOI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1467),
.A2(n_1416),
.B(n_1497),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1483),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1483),
.Y(n_1553)
);

NAND3xp33_ASAP7_75t_L g1554 ( 
.A(n_1502),
.B(n_1523),
.C(n_1520),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1431),
.B(n_1526),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1515),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1478),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1431),
.B(n_1440),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1485),
.A2(n_1484),
.B(n_1471),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1524),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1434),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1434),
.Y(n_1562)
);

CKINVDCx20_ASAP7_75t_R g1563 ( 
.A(n_1505),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1441),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1441),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_1401),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1455),
.Y(n_1567)
);

OAI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1506),
.A2(n_1525),
.B(n_1424),
.Y(n_1568)
);

OAI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1424),
.A2(n_1510),
.B(n_1527),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1403),
.B(n_1486),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1403),
.B(n_1486),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1490),
.Y(n_1572)
);

OA21x2_ASAP7_75t_L g1573 ( 
.A1(n_1448),
.A2(n_1426),
.B(n_1484),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1418),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1418),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1472),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1456),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1435),
.B(n_1415),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1456),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1448),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1499),
.B(n_1509),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1435),
.B(n_1413),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1477),
.Y(n_1583)
);

OAI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1492),
.A2(n_1527),
.B(n_1510),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1409),
.B(n_1429),
.Y(n_1585)
);

AND2x2_ASAP7_75t_SL g1586 ( 
.A(n_1495),
.B(n_1496),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1519),
.Y(n_1587)
);

INVx4_ASAP7_75t_L g1588 ( 
.A(n_1475),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1511),
.B(n_1495),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1410),
.Y(n_1590)
);

OR2x2_ASAP7_75t_SL g1591 ( 
.A(n_1405),
.B(n_1501),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1519),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1475),
.Y(n_1593)
);

INVxp33_ASAP7_75t_L g1594 ( 
.A(n_1452),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1410),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1429),
.B(n_1407),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1465),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1496),
.B(n_1521),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1517),
.B(n_1522),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1407),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1433),
.B(n_1413),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1459),
.B(n_1462),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1485),
.Y(n_1603)
);

BUFx3_ASAP7_75t_L g1604 ( 
.A(n_1463),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1419),
.Y(n_1605)
);

NOR2xp67_ASAP7_75t_SL g1606 ( 
.A(n_1500),
.B(n_1528),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1462),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1419),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1513),
.B(n_1450),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1512),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1425),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1442),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1442),
.Y(n_1613)
);

A2O1A1Ixp33_ASAP7_75t_L g1614 ( 
.A1(n_1584),
.A2(n_1449),
.B(n_1491),
.C(n_1460),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1540),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1554),
.A2(n_1516),
.B1(n_1458),
.B2(n_1463),
.Y(n_1616)
);

AO32x2_ASAP7_75t_L g1617 ( 
.A1(n_1546),
.A2(n_1503),
.A3(n_1444),
.B1(n_1417),
.B2(n_1420),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1569),
.A2(n_1464),
.B(n_1442),
.Y(n_1618)
);

BUFx12f_ASAP7_75t_L g1619 ( 
.A(n_1591),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1583),
.B(n_1491),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1583),
.B(n_1445),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1594),
.B(n_1446),
.Y(n_1622)
);

AND2x2_ASAP7_75t_SL g1623 ( 
.A(n_1581),
.B(n_1493),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1568),
.B(n_1438),
.Y(n_1624)
);

AO32x2_ASAP7_75t_L g1625 ( 
.A1(n_1566),
.A2(n_1444),
.A3(n_1503),
.B1(n_1417),
.B2(n_1420),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1550),
.B(n_1518),
.Y(n_1626)
);

A2O1A1Ixp33_ASAP7_75t_L g1627 ( 
.A1(n_1547),
.A2(n_1453),
.B(n_1498),
.C(n_1504),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1540),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1536),
.B(n_1438),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1586),
.A2(n_1443),
.B1(n_1514),
.B2(n_1400),
.Y(n_1630)
);

AOI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1539),
.A2(n_1439),
.B1(n_1451),
.B2(n_1420),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1549),
.B(n_1542),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1541),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1551),
.B(n_1592),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1543),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1549),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1549),
.B(n_1587),
.Y(n_1637)
);

A2O1A1Ixp33_ASAP7_75t_L g1638 ( 
.A1(n_1581),
.A2(n_1461),
.B(n_1447),
.C(n_1470),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1550),
.B(n_1545),
.Y(n_1639)
);

INVx2_ASAP7_75t_SL g1640 ( 
.A(n_1602),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1587),
.B(n_1602),
.Y(n_1641)
);

OAI211xp5_ASAP7_75t_L g1642 ( 
.A1(n_1551),
.A2(n_1454),
.B(n_1508),
.C(n_1428),
.Y(n_1642)
);

AOI221xp5_ASAP7_75t_L g1643 ( 
.A1(n_1561),
.A2(n_1507),
.B1(n_1430),
.B2(n_1464),
.C(n_1411),
.Y(n_1643)
);

CKINVDCx11_ASAP7_75t_R g1644 ( 
.A(n_1563),
.Y(n_1644)
);

OAI21x1_ASAP7_75t_SL g1645 ( 
.A1(n_1588),
.A2(n_1601),
.B(n_1585),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1567),
.B(n_1421),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1531),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1555),
.B(n_1421),
.Y(n_1648)
);

O2A1O1Ixp5_ASAP7_75t_L g1649 ( 
.A1(n_1578),
.A2(n_1494),
.B(n_1562),
.C(n_1561),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1556),
.Y(n_1650)
);

OAI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1574),
.A2(n_1575),
.B(n_1577),
.Y(n_1651)
);

OA21x2_ASAP7_75t_L g1652 ( 
.A1(n_1559),
.A2(n_1532),
.B(n_1579),
.Y(n_1652)
);

OA21x2_ASAP7_75t_L g1653 ( 
.A1(n_1559),
.A2(n_1579),
.B(n_1577),
.Y(n_1653)
);

OAI211xp5_ASAP7_75t_L g1654 ( 
.A1(n_1574),
.A2(n_1575),
.B(n_1529),
.C(n_1596),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1586),
.A2(n_1589),
.B1(n_1529),
.B2(n_1595),
.Y(n_1655)
);

NAND3xp33_ASAP7_75t_L g1656 ( 
.A(n_1562),
.B(n_1533),
.C(n_1572),
.Y(n_1656)
);

A2O1A1Ixp33_ASAP7_75t_L g1657 ( 
.A1(n_1589),
.A2(n_1582),
.B(n_1599),
.C(n_1598),
.Y(n_1657)
);

A2O1A1Ixp33_ASAP7_75t_L g1658 ( 
.A1(n_1582),
.A2(n_1598),
.B(n_1599),
.C(n_1590),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1607),
.B(n_1534),
.Y(n_1659)
);

A2O1A1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1590),
.A2(n_1595),
.B(n_1571),
.C(n_1570),
.Y(n_1660)
);

OAI211xp5_ASAP7_75t_SL g1661 ( 
.A1(n_1603),
.A2(n_1610),
.B(n_1605),
.C(n_1608),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1560),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1609),
.B(n_1557),
.Y(n_1663)
);

CKINVDCx14_ASAP7_75t_R g1664 ( 
.A(n_1604),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1609),
.B(n_1557),
.Y(n_1665)
);

A2O1A1Ixp33_ASAP7_75t_L g1666 ( 
.A1(n_1570),
.A2(n_1571),
.B(n_1600),
.C(n_1580),
.Y(n_1666)
);

A2O1A1Ixp33_ASAP7_75t_L g1667 ( 
.A1(n_1600),
.A2(n_1580),
.B(n_1558),
.C(n_1530),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1611),
.B(n_1612),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1613),
.B(n_1544),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1613),
.B(n_1544),
.Y(n_1670)
);

A2O1A1Ixp33_ASAP7_75t_L g1671 ( 
.A1(n_1530),
.A2(n_1564),
.B(n_1565),
.C(n_1603),
.Y(n_1671)
);

OAI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1533),
.A2(n_1605),
.B(n_1610),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1659),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1615),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1628),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1632),
.B(n_1548),
.Y(n_1676)
);

INVxp67_ASAP7_75t_SL g1677 ( 
.A(n_1634),
.Y(n_1677)
);

AOI21x1_ASAP7_75t_L g1678 ( 
.A1(n_1647),
.A2(n_1552),
.B(n_1553),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1642),
.B(n_1664),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1633),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1635),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1664),
.B(n_1535),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1655),
.A2(n_1623),
.B1(n_1651),
.B2(n_1656),
.Y(n_1683)
);

INVxp67_ASAP7_75t_L g1684 ( 
.A(n_1646),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1663),
.B(n_1548),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1627),
.A2(n_1588),
.B1(n_1591),
.B2(n_1593),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1639),
.B(n_1552),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1623),
.A2(n_1573),
.B1(n_1597),
.B2(n_1537),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1669),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1629),
.B(n_1548),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1625),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1650),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1665),
.B(n_1573),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1662),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1630),
.A2(n_1573),
.B1(n_1597),
.B2(n_1538),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1670),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1641),
.B(n_1533),
.Y(n_1697)
);

INVx1_ASAP7_75t_SL g1698 ( 
.A(n_1644),
.Y(n_1698)
);

BUFx2_ASAP7_75t_L g1699 ( 
.A(n_1625),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1668),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1639),
.B(n_1636),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1636),
.B(n_1553),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1640),
.B(n_1637),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1653),
.B(n_1531),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1636),
.B(n_1576),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1672),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1644),
.B(n_1606),
.Y(n_1707)
);

INVxp67_ASAP7_75t_L g1708 ( 
.A(n_1648),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1625),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1685),
.B(n_1693),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1683),
.A2(n_1657),
.B1(n_1660),
.B2(n_1658),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1677),
.B(n_1652),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1691),
.Y(n_1713)
);

OAI221xp5_ASAP7_75t_SL g1714 ( 
.A1(n_1691),
.A2(n_1658),
.B1(n_1660),
.B2(n_1654),
.C(n_1666),
.Y(n_1714)
);

AO21x2_ASAP7_75t_L g1715 ( 
.A1(n_1704),
.A2(n_1667),
.B(n_1666),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1706),
.B(n_1652),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1698),
.Y(n_1717)
);

AOI21x1_ASAP7_75t_L g1718 ( 
.A1(n_1678),
.A2(n_1606),
.B(n_1645),
.Y(n_1718)
);

INVx4_ASAP7_75t_L g1719 ( 
.A(n_1699),
.Y(n_1719)
);

INVx3_ASAP7_75t_L g1720 ( 
.A(n_1705),
.Y(n_1720)
);

BUFx2_ASAP7_75t_L g1721 ( 
.A(n_1699),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1685),
.B(n_1652),
.Y(n_1722)
);

NOR3xp33_ASAP7_75t_SL g1723 ( 
.A(n_1707),
.B(n_1616),
.C(n_1638),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1709),
.B(n_1617),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1674),
.Y(n_1725)
);

INVxp67_ASAP7_75t_L g1726 ( 
.A(n_1709),
.Y(n_1726)
);

NOR3xp33_ASAP7_75t_SL g1727 ( 
.A(n_1679),
.B(n_1638),
.C(n_1627),
.Y(n_1727)
);

INVx5_ASAP7_75t_SL g1728 ( 
.A(n_1702),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1674),
.Y(n_1729)
);

AOI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1695),
.A2(n_1624),
.B1(n_1631),
.B2(n_1619),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1675),
.Y(n_1731)
);

AOI221xp5_ASAP7_75t_L g1732 ( 
.A1(n_1697),
.A2(n_1667),
.B1(n_1671),
.B2(n_1649),
.C(n_1624),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1676),
.B(n_1617),
.Y(n_1733)
);

NOR2x1_ASAP7_75t_L g1734 ( 
.A(n_1682),
.B(n_1661),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_SL g1735 ( 
.A(n_1686),
.B(n_1614),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1675),
.Y(n_1736)
);

AOI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1688),
.A2(n_1619),
.B1(n_1643),
.B2(n_1618),
.Y(n_1737)
);

BUFx3_ASAP7_75t_L g1738 ( 
.A(n_1702),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1676),
.B(n_1617),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1705),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1703),
.B(n_1617),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1703),
.B(n_1701),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_1680),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1743),
.B(n_1681),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1733),
.B(n_1700),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1726),
.B(n_1689),
.Y(n_1746)
);

INVx3_ASAP7_75t_L g1747 ( 
.A(n_1728),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1743),
.B(n_1681),
.Y(n_1748)
);

NOR3xp33_ASAP7_75t_L g1749 ( 
.A(n_1714),
.B(n_1614),
.C(n_1678),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1725),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1715),
.Y(n_1751)
);

BUFx3_ASAP7_75t_L g1752 ( 
.A(n_1717),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1715),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1738),
.B(n_1740),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1725),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1733),
.B(n_1673),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1729),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1729),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1715),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1731),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1731),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1715),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1713),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1736),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1715),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1739),
.B(n_1708),
.Y(n_1766)
);

NOR2x1_ASAP7_75t_L g1767 ( 
.A(n_1734),
.B(n_1621),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1726),
.B(n_1696),
.Y(n_1768)
);

INVx6_ASAP7_75t_L g1769 ( 
.A(n_1719),
.Y(n_1769)
);

INVxp67_ASAP7_75t_L g1770 ( 
.A(n_1734),
.Y(n_1770)
);

NOR3xp33_ASAP7_75t_SL g1771 ( 
.A(n_1714),
.B(n_1692),
.C(n_1694),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1739),
.B(n_1684),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1739),
.B(n_1690),
.Y(n_1773)
);

BUFx2_ASAP7_75t_L g1774 ( 
.A(n_1719),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1738),
.B(n_1687),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1713),
.B(n_1696),
.Y(n_1776)
);

AND2x4_ASAP7_75t_L g1777 ( 
.A(n_1720),
.B(n_1687),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1771),
.B(n_1724),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1750),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1767),
.B(n_1710),
.Y(n_1780)
);

INVxp67_ASAP7_75t_L g1781 ( 
.A(n_1770),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1751),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1750),
.Y(n_1783)
);

AOI32xp33_ASAP7_75t_L g1784 ( 
.A1(n_1767),
.A2(n_1749),
.A3(n_1711),
.B1(n_1724),
.B2(n_1735),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1755),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1773),
.B(n_1710),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1755),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1768),
.B(n_1713),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1751),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1747),
.B(n_1721),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1747),
.B(n_1721),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1771),
.B(n_1724),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1757),
.Y(n_1793)
);

INVxp33_ASAP7_75t_L g1794 ( 
.A(n_1752),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1757),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1751),
.Y(n_1796)
);

AOI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1749),
.A2(n_1711),
.B1(n_1735),
.B2(n_1732),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1772),
.B(n_1710),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1772),
.B(n_1741),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1772),
.B(n_1741),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1758),
.Y(n_1801)
);

BUFx2_ASAP7_75t_L g1802 ( 
.A(n_1770),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1753),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1775),
.B(n_1741),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1775),
.B(n_1721),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1773),
.B(n_1719),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1758),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1775),
.B(n_1742),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1760),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1753),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1760),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1773),
.B(n_1722),
.Y(n_1812)
);

INVxp67_ASAP7_75t_SL g1813 ( 
.A(n_1763),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1761),
.Y(n_1814)
);

NAND2x1p5_ASAP7_75t_L g1815 ( 
.A(n_1747),
.B(n_1718),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1753),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1775),
.B(n_1742),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1766),
.B(n_1742),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1768),
.B(n_1716),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1747),
.B(n_1719),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1746),
.B(n_1716),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1763),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1761),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1764),
.Y(n_1824)
);

AOI21xp33_ASAP7_75t_L g1825 ( 
.A1(n_1784),
.A2(n_1762),
.B(n_1759),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1797),
.B(n_1766),
.Y(n_1826)
);

NOR3xp33_ASAP7_75t_L g1827 ( 
.A(n_1802),
.B(n_1718),
.C(n_1759),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1788),
.B(n_1776),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1822),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1797),
.B(n_1766),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1818),
.B(n_1754),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1822),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1779),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1779),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1783),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1786),
.B(n_1754),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1802),
.B(n_1756),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1788),
.B(n_1778),
.Y(n_1838)
);

INVxp33_ASAP7_75t_L g1839 ( 
.A(n_1794),
.Y(n_1839)
);

OAI21xp33_ASAP7_75t_L g1840 ( 
.A1(n_1784),
.A2(n_1727),
.B(n_1746),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1783),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1778),
.A2(n_1792),
.B1(n_1732),
.B2(n_1737),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1781),
.B(n_1756),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1781),
.B(n_1792),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1786),
.B(n_1754),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1812),
.B(n_1776),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1786),
.B(n_1798),
.Y(n_1847)
);

NOR3xp33_ASAP7_75t_L g1848 ( 
.A(n_1813),
.B(n_1762),
.C(n_1759),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1798),
.B(n_1756),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1813),
.B(n_1818),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1780),
.B(n_1754),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1780),
.B(n_1777),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1790),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1806),
.B(n_1745),
.Y(n_1854)
);

INVx1_ASAP7_75t_SL g1855 ( 
.A(n_1790),
.Y(n_1855)
);

NAND3xp33_ASAP7_75t_L g1856 ( 
.A(n_1790),
.B(n_1727),
.C(n_1774),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1808),
.B(n_1752),
.Y(n_1857)
);

INVx1_ASAP7_75t_SL g1858 ( 
.A(n_1790),
.Y(n_1858)
);

HB1xp67_ASAP7_75t_L g1859 ( 
.A(n_1785),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1791),
.B(n_1774),
.Y(n_1860)
);

NAND3xp33_ASAP7_75t_L g1861 ( 
.A(n_1791),
.B(n_1787),
.C(n_1785),
.Y(n_1861)
);

INVxp67_ASAP7_75t_L g1862 ( 
.A(n_1857),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1839),
.B(n_1752),
.Y(n_1863)
);

NAND3xp33_ASAP7_75t_SL g1864 ( 
.A(n_1840),
.B(n_1842),
.C(n_1830),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1836),
.B(n_1808),
.Y(n_1865)
);

NAND4xp75_ASAP7_75t_L g1866 ( 
.A(n_1844),
.B(n_1723),
.C(n_1765),
.D(n_1762),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1826),
.B(n_1806),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1859),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1839),
.B(n_1806),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1855),
.B(n_1858),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1836),
.B(n_1817),
.Y(n_1871)
);

AOI222xp33_ASAP7_75t_L g1872 ( 
.A1(n_1843),
.A2(n_1765),
.B1(n_1800),
.B2(n_1799),
.C1(n_1722),
.C2(n_1712),
.Y(n_1872)
);

INVx3_ASAP7_75t_L g1873 ( 
.A(n_1831),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1833),
.Y(n_1874)
);

AOI21x1_ASAP7_75t_L g1875 ( 
.A1(n_1860),
.A2(n_1791),
.B(n_1820),
.Y(n_1875)
);

INVxp67_ASAP7_75t_SL g1876 ( 
.A(n_1857),
.Y(n_1876)
);

INVx2_ASAP7_75t_SL g1877 ( 
.A(n_1853),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1838),
.B(n_1799),
.Y(n_1878)
);

OAI22xp33_ASAP7_75t_L g1879 ( 
.A1(n_1838),
.A2(n_1719),
.B1(n_1812),
.B2(n_1765),
.Y(n_1879)
);

AOI21xp33_ASAP7_75t_L g1880 ( 
.A1(n_1825),
.A2(n_1835),
.B(n_1834),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1841),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1829),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1845),
.B(n_1817),
.Y(n_1883)
);

OAI211xp5_ASAP7_75t_SL g1884 ( 
.A1(n_1860),
.A2(n_1723),
.B(n_1821),
.C(n_1819),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1845),
.B(n_1804),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1831),
.B(n_1804),
.Y(n_1886)
);

NOR2xp67_ASAP7_75t_SL g1887 ( 
.A(n_1856),
.B(n_1604),
.Y(n_1887)
);

OAI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1847),
.A2(n_1769),
.B1(n_1800),
.B2(n_1820),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1873),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1874),
.Y(n_1890)
);

OAI21xp5_ASAP7_75t_L g1891 ( 
.A1(n_1866),
.A2(n_1827),
.B(n_1861),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1881),
.Y(n_1892)
);

INVx1_ASAP7_75t_SL g1893 ( 
.A(n_1873),
.Y(n_1893)
);

INVxp67_ASAP7_75t_L g1894 ( 
.A(n_1863),
.Y(n_1894)
);

OAI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1866),
.A2(n_1831),
.B1(n_1837),
.B2(n_1849),
.Y(n_1895)
);

OAI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1862),
.A2(n_1850),
.B1(n_1769),
.B2(n_1854),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1886),
.B(n_1851),
.Y(n_1897)
);

AOI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1864),
.A2(n_1884),
.B1(n_1887),
.B2(n_1878),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1882),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1882),
.Y(n_1900)
);

XNOR2x1_ASAP7_75t_L g1901 ( 
.A(n_1870),
.B(n_1815),
.Y(n_1901)
);

AOI32xp33_ASAP7_75t_L g1902 ( 
.A1(n_1879),
.A2(n_1848),
.A3(n_1791),
.B1(n_1851),
.B2(n_1852),
.Y(n_1902)
);

OAI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1875),
.A2(n_1853),
.B(n_1815),
.Y(n_1903)
);

INVx3_ASAP7_75t_L g1904 ( 
.A(n_1873),
.Y(n_1904)
);

INVxp67_ASAP7_75t_L g1905 ( 
.A(n_1876),
.Y(n_1905)
);

HB1xp67_ASAP7_75t_L g1906 ( 
.A(n_1877),
.Y(n_1906)
);

AOI22xp5_ASAP7_75t_SL g1907 ( 
.A1(n_1868),
.A2(n_1815),
.B1(n_1820),
.B2(n_1832),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1887),
.B(n_1828),
.Y(n_1908)
);

INVxp67_ASAP7_75t_L g1909 ( 
.A(n_1877),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1905),
.B(n_1867),
.Y(n_1910)
);

HB1xp67_ASAP7_75t_L g1911 ( 
.A(n_1906),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1906),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1909),
.Y(n_1913)
);

BUFx2_ASAP7_75t_L g1914 ( 
.A(n_1904),
.Y(n_1914)
);

INVxp67_ASAP7_75t_SL g1915 ( 
.A(n_1905),
.Y(n_1915)
);

OA22x2_ASAP7_75t_L g1916 ( 
.A1(n_1891),
.A2(n_1869),
.B1(n_1886),
.B2(n_1888),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1893),
.B(n_1828),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1909),
.Y(n_1918)
);

OAI21xp33_ASAP7_75t_L g1919 ( 
.A1(n_1898),
.A2(n_1871),
.B(n_1865),
.Y(n_1919)
);

OAI31xp33_ASAP7_75t_SL g1920 ( 
.A1(n_1895),
.A2(n_1880),
.A3(n_1883),
.B(n_1865),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1889),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1904),
.B(n_1885),
.Y(n_1922)
);

AOI211xp5_ASAP7_75t_SL g1923 ( 
.A1(n_1913),
.A2(n_1894),
.B(n_1908),
.C(n_1896),
.Y(n_1923)
);

AOI322xp5_ASAP7_75t_L g1924 ( 
.A1(n_1915),
.A2(n_1900),
.A3(n_1899),
.B1(n_1894),
.B2(n_1890),
.C1(n_1892),
.C2(n_1897),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1911),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1914),
.B(n_1915),
.Y(n_1926)
);

NAND4xp25_ASAP7_75t_L g1927 ( 
.A(n_1920),
.B(n_1910),
.C(n_1918),
.D(n_1912),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1911),
.B(n_1885),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1917),
.B(n_1902),
.Y(n_1929)
);

NAND4xp25_ASAP7_75t_SL g1930 ( 
.A(n_1922),
.B(n_1872),
.C(n_1903),
.D(n_1883),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1921),
.B(n_1871),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1916),
.B(n_1852),
.Y(n_1932)
);

NAND4xp75_ASAP7_75t_L g1933 ( 
.A(n_1916),
.B(n_1901),
.C(n_1907),
.D(n_1805),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1919),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1922),
.B(n_1805),
.Y(n_1935)
);

OAI22xp5_ASAP7_75t_L g1936 ( 
.A1(n_1933),
.A2(n_1846),
.B1(n_1875),
.B2(n_1821),
.Y(n_1936)
);

OAI221xp5_ASAP7_75t_L g1937 ( 
.A1(n_1927),
.A2(n_1929),
.B1(n_1932),
.B2(n_1926),
.C(n_1934),
.Y(n_1937)
);

AOI221xp5_ASAP7_75t_SL g1938 ( 
.A1(n_1927),
.A2(n_1824),
.B1(n_1823),
.B2(n_1787),
.C(n_1793),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1928),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1925),
.Y(n_1940)
);

NAND2x1_ASAP7_75t_L g1941 ( 
.A(n_1935),
.B(n_1820),
.Y(n_1941)
);

NAND4xp25_ASAP7_75t_L g1942 ( 
.A(n_1937),
.B(n_1923),
.C(n_1924),
.D(n_1931),
.Y(n_1942)
);

AOI221xp5_ASAP7_75t_L g1943 ( 
.A1(n_1936),
.A2(n_1930),
.B1(n_1782),
.B2(n_1789),
.C(n_1816),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1938),
.B(n_1793),
.Y(n_1944)
);

AOI221xp5_ASAP7_75t_L g1945 ( 
.A1(n_1940),
.A2(n_1810),
.B1(n_1803),
.B2(n_1782),
.C(n_1796),
.Y(n_1945)
);

OAI221xp5_ASAP7_75t_SL g1946 ( 
.A1(n_1939),
.A2(n_1819),
.B1(n_1737),
.B2(n_1730),
.C(n_1789),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1941),
.Y(n_1947)
);

AOI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1936),
.A2(n_1815),
.B1(n_1769),
.B2(n_1816),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1947),
.Y(n_1949)
);

XNOR2xp5_ASAP7_75t_L g1950 ( 
.A(n_1942),
.B(n_1622),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1944),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1948),
.B(n_1745),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1945),
.Y(n_1953)
);

NOR3xp33_ASAP7_75t_L g1954 ( 
.A(n_1943),
.B(n_1789),
.C(n_1782),
.Y(n_1954)
);

OAI211xp5_ASAP7_75t_SL g1955 ( 
.A1(n_1951),
.A2(n_1946),
.B(n_1824),
.C(n_1823),
.Y(n_1955)
);

NAND4xp25_ASAP7_75t_L g1956 ( 
.A(n_1949),
.B(n_1730),
.C(n_1814),
.D(n_1811),
.Y(n_1956)
);

AOI21xp33_ASAP7_75t_SL g1957 ( 
.A1(n_1950),
.A2(n_1801),
.B(n_1795),
.Y(n_1957)
);

XOR2xp5_ASAP7_75t_L g1958 ( 
.A(n_1956),
.B(n_1951),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1958),
.Y(n_1959)
);

OAI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1959),
.A2(n_1955),
.B(n_1953),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1959),
.Y(n_1961)
);

OAI22xp5_ASAP7_75t_L g1962 ( 
.A1(n_1961),
.A2(n_1957),
.B1(n_1952),
.B2(n_1954),
.Y(n_1962)
);

OAI22xp5_ASAP7_75t_SL g1963 ( 
.A1(n_1960),
.A2(n_1769),
.B1(n_1814),
.B2(n_1811),
.Y(n_1963)
);

AOI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1962),
.A2(n_1801),
.B(n_1795),
.Y(n_1964)
);

OAI22xp5_ASAP7_75t_L g1965 ( 
.A1(n_1963),
.A2(n_1809),
.B1(n_1807),
.B2(n_1769),
.Y(n_1965)
);

OAI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1964),
.A2(n_1807),
.B1(n_1809),
.B2(n_1810),
.Y(n_1966)
);

AO21x1_ASAP7_75t_L g1967 ( 
.A1(n_1965),
.A2(n_1803),
.B(n_1796),
.Y(n_1967)
);

AO21x2_ASAP7_75t_L g1968 ( 
.A1(n_1967),
.A2(n_1803),
.B(n_1796),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1968),
.Y(n_1969)
);

OAI221xp5_ASAP7_75t_R g1970 ( 
.A1(n_1969),
.A2(n_1966),
.B1(n_1816),
.B2(n_1810),
.C(n_1748),
.Y(n_1970)
);

AOI211xp5_ASAP7_75t_L g1971 ( 
.A1(n_1970),
.A2(n_1620),
.B(n_1626),
.C(n_1744),
.Y(n_1971)
);


endmodule