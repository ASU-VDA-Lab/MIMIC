module fake_jpeg_5248_n_33 (n_3, n_2, n_1, n_0, n_4, n_5, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_33;

wire n_13;
wire n_21;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_SL g12 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_12),
.B(n_13),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_6),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_13)
);

AOI22xp33_ASAP7_75t_L g14 ( 
.A1(n_11),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_8),
.B(n_5),
.Y(n_15)
);

AND2x6_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_11),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_8),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_15),
.B1(n_12),
.B2(n_13),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_20),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_22),
.C(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_17),
.C(n_15),
.Y(n_25)
);

BUFx12f_ASAP7_75t_SL g26 ( 
.A(n_25),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_23),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_29),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_9),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_28),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_26),
.B(n_9),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_10),
.B(n_30),
.Y(n_33)
);


endmodule