module fake_ibex_1331_n_6672 (n_151, n_1084, n_85, n_599, n_778, n_822, n_1042, n_507, n_743, n_1060, n_540, n_754, n_395, n_1104, n_1011, n_84, n_64, n_992, n_1148, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_1041, n_688, n_130, n_1090, n_177, n_1110, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_1097, n_9, n_1079, n_1031, n_1143, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_972, n_981, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_1067, n_255, n_175, n_586, n_773, n_994, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_962, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_1080, n_1162, n_957, n_1015, n_678, n_663, n_969, n_194, n_249, n_334, n_1125, n_634, n_733, n_961, n_991, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_1034, n_1152, n_371, n_974, n_1036, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_1018, n_1044, n_1106, n_1129, n_40, n_90, n_17, n_74, n_449, n_1131, n_547, n_176, n_1134, n_727, n_1138, n_58, n_1077, n_43, n_216, n_996, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_1045, n_753, n_645, n_500, n_747, n_963, n_1147, n_542, n_114, n_236, n_900, n_34, n_376, n_1098, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_1096, n_105, n_187, n_667, n_884, n_1061, n_1, n_154, n_682, n_850, n_182, n_196, n_1140, n_326, n_327, n_879, n_89, n_1056, n_50, n_723, n_144, n_170, n_270, n_1144, n_346, n_383, n_113, n_886, n_840, n_1010, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_1029, n_859, n_259, n_276, n_339, n_470, n_770, n_965, n_210, n_348, n_1109, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_989, n_373, n_1051, n_854, n_1008, n_458, n_244, n_73, n_1053, n_1112, n_343, n_310, n_714, n_1076, n_1032, n_936, n_703, n_426, n_323, n_469, n_829, n_1099, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_967, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_1055, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_1103, n_1161, n_121, n_527, n_893, n_590, n_1025, n_465, n_1057, n_1068, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_1013, n_982, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_1024, n_13, n_637, n_1141, n_122, n_523, n_116, n_694, n_787, n_977, n_1075, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_1130, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_1081, n_215, n_1153, n_279, n_49, n_1037, n_374, n_235, n_464, n_538, n_669, n_838, n_987, n_1155, n_750, n_1021, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_1117, n_30, n_1101, n_518, n_367, n_221, n_1052, n_852, n_789, n_1133, n_880, n_654, n_1083, n_656, n_1014, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_1023, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_1001, n_156, n_570, n_126, n_1116, n_623, n_585, n_1030, n_1094, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_1082, n_222, n_1137, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_980, n_454, n_1070, n_1074, n_777, n_1017, n_295, n_730, n_331, n_1120, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_968, n_619, n_1089, n_536, n_1124, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_1064, n_1071, n_207, n_922, n_438, n_851, n_993, n_1012, n_1028, n_689, n_960, n_1022, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_1151, n_145, n_65, n_1135, n_973, n_1146, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_999, n_1038, n_1092, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_1009, n_635, n_979, n_844, n_1066, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_1020, n_847, n_830, n_1062, n_1142, n_1004, n_473, n_1027, n_445, n_629, n_335, n_413, n_1072, n_82, n_263, n_1069, n_27, n_573, n_353, n_966, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_1007, n_1126, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_1006, n_402, n_725, n_180, n_369, n_976, n_596, n_201, n_699, n_14, n_1063, n_351, n_368, n_456, n_834, n_257, n_77, n_998, n_935, n_869, n_1115, n_925, n_718, n_801, n_918, n_1054, n_44, n_672, n_1100, n_1039, n_722, n_401, n_1046, n_553, n_554, n_1078, n_1043, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_1049, n_1086, n_763, n_1158, n_745, n_329, n_1149, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_1065, n_592, n_986, n_495, n_762, n_410, n_905, n_308, n_975, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_1160, n_512, n_615, n_950, n_685, n_1026, n_283, n_366, n_397, n_111, n_803, n_894, n_1033, n_1118, n_692, n_36, n_627, n_990, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_1087, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_971, n_101, n_190, n_906, n_138, n_650, n_776, n_1114, n_409, n_1093, n_582, n_978, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_1019, n_1059, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_1107, n_223, n_381, n_1073, n_1108, n_525, n_815, n_919, n_780, n_535, n_1002, n_382, n_502, n_681, n_633, n_1111, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_1128, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_997, n_833, n_1145, n_217, n_324, n_391, n_831, n_537, n_1113, n_728, n_78, n_805, n_670, n_820, n_20, n_1132, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_1164, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_1016, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_1139, n_870, n_46, n_284, n_811, n_1047, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_1040, n_476, n_792, n_461, n_575, n_313, n_1159, n_1119, n_903, n_1154, n_519, n_345, n_408, n_119, n_1085, n_361, n_1095, n_455, n_1136, n_419, n_774, n_72, n_1048, n_319, n_1091, n_195, n_885, n_513, n_212, n_588, n_877, n_1121, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_1088, n_896, n_97, n_197, n_528, n_181, n_1005, n_131, n_123, n_1102, n_631, n_683, n_260, n_620, n_794, n_836, n_1150, n_462, n_302, n_450, n_443, n_686, n_985, n_572, n_1165, n_867, n_983, n_1003, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_970, n_491, n_1122, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_1058, n_1105, n_107, n_1163, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_964, n_424, n_565, n_916, n_823, n_1123, n_701, n_271, n_995, n_241, n_68, n_503, n_292, n_807, n_984, n_394, n_79, n_1000, n_81, n_35, n_364, n_687, n_895, n_988, n_159, n_202, n_231, n_298, n_587, n_1035, n_760, n_1157, n_751, n_806, n_1127, n_932, n_160, n_657, n_764, n_184, n_1156, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_1050, n_6672);

input n_151;
input n_1084;
input n_85;
input n_599;
input n_778;
input n_822;
input n_1042;
input n_507;
input n_743;
input n_1060;
input n_540;
input n_754;
input n_395;
input n_1104;
input n_1011;
input n_84;
input n_64;
input n_992;
input n_1148;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_1041;
input n_688;
input n_130;
input n_1090;
input n_177;
input n_1110;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_1097;
input n_9;
input n_1079;
input n_1031;
input n_1143;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_972;
input n_981;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_1067;
input n_255;
input n_175;
input n_586;
input n_773;
input n_994;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_962;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_1080;
input n_1162;
input n_957;
input n_1015;
input n_678;
input n_663;
input n_969;
input n_194;
input n_249;
input n_334;
input n_1125;
input n_634;
input n_733;
input n_961;
input n_991;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_1034;
input n_1152;
input n_371;
input n_974;
input n_1036;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_1018;
input n_1044;
input n_1106;
input n_1129;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_1131;
input n_547;
input n_176;
input n_1134;
input n_727;
input n_1138;
input n_58;
input n_1077;
input n_43;
input n_216;
input n_996;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_1045;
input n_753;
input n_645;
input n_500;
input n_747;
input n_963;
input n_1147;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_1098;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_1096;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1061;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_1140;
input n_326;
input n_327;
input n_879;
input n_89;
input n_1056;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_1144;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_1010;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_1029;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_965;
input n_210;
input n_348;
input n_1109;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_989;
input n_373;
input n_1051;
input n_854;
input n_1008;
input n_458;
input n_244;
input n_73;
input n_1053;
input n_1112;
input n_343;
input n_310;
input n_714;
input n_1076;
input n_1032;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_1099;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_967;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_1055;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_1103;
input n_1161;
input n_121;
input n_527;
input n_893;
input n_590;
input n_1025;
input n_465;
input n_1057;
input n_1068;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_1013;
input n_982;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_1024;
input n_13;
input n_637;
input n_1141;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_977;
input n_1075;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_1130;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_1081;
input n_215;
input n_1153;
input n_279;
input n_49;
input n_1037;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_987;
input n_1155;
input n_750;
input n_1021;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_1117;
input n_30;
input n_1101;
input n_518;
input n_367;
input n_221;
input n_1052;
input n_852;
input n_789;
input n_1133;
input n_880;
input n_654;
input n_1083;
input n_656;
input n_1014;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_1023;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_1001;
input n_156;
input n_570;
input n_126;
input n_1116;
input n_623;
input n_585;
input n_1030;
input n_1094;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_1082;
input n_222;
input n_1137;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_980;
input n_454;
input n_1070;
input n_1074;
input n_777;
input n_1017;
input n_295;
input n_730;
input n_331;
input n_1120;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_968;
input n_619;
input n_1089;
input n_536;
input n_1124;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_1064;
input n_1071;
input n_207;
input n_922;
input n_438;
input n_851;
input n_993;
input n_1012;
input n_1028;
input n_689;
input n_960;
input n_1022;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_1151;
input n_145;
input n_65;
input n_1135;
input n_973;
input n_1146;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_999;
input n_1038;
input n_1092;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_1009;
input n_635;
input n_979;
input n_844;
input n_1066;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_1020;
input n_847;
input n_830;
input n_1062;
input n_1142;
input n_1004;
input n_473;
input n_1027;
input n_445;
input n_629;
input n_335;
input n_413;
input n_1072;
input n_82;
input n_263;
input n_1069;
input n_27;
input n_573;
input n_353;
input n_966;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_1007;
input n_1126;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_1006;
input n_402;
input n_725;
input n_180;
input n_369;
input n_976;
input n_596;
input n_201;
input n_699;
input n_14;
input n_1063;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_998;
input n_935;
input n_869;
input n_1115;
input n_925;
input n_718;
input n_801;
input n_918;
input n_1054;
input n_44;
input n_672;
input n_1100;
input n_1039;
input n_722;
input n_401;
input n_1046;
input n_553;
input n_554;
input n_1078;
input n_1043;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_1049;
input n_1086;
input n_763;
input n_1158;
input n_745;
input n_329;
input n_1149;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_1065;
input n_592;
input n_986;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_975;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_1160;
input n_512;
input n_615;
input n_950;
input n_685;
input n_1026;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_1033;
input n_1118;
input n_692;
input n_36;
input n_627;
input n_990;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_1087;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_971;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_1114;
input n_409;
input n_1093;
input n_582;
input n_978;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_1019;
input n_1059;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_1107;
input n_223;
input n_381;
input n_1073;
input n_1108;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_1002;
input n_382;
input n_502;
input n_681;
input n_633;
input n_1111;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_1128;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_997;
input n_833;
input n_1145;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_1113;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_1132;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_1164;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_1016;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_1139;
input n_870;
input n_46;
input n_284;
input n_811;
input n_1047;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_1040;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_1159;
input n_1119;
input n_903;
input n_1154;
input n_519;
input n_345;
input n_408;
input n_119;
input n_1085;
input n_361;
input n_1095;
input n_455;
input n_1136;
input n_419;
input n_774;
input n_72;
input n_1048;
input n_319;
input n_1091;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_1121;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_1088;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_1005;
input n_131;
input n_123;
input n_1102;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_1150;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_985;
input n_572;
input n_1165;
input n_867;
input n_983;
input n_1003;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_970;
input n_491;
input n_1122;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_1058;
input n_1105;
input n_107;
input n_1163;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_964;
input n_424;
input n_565;
input n_916;
input n_823;
input n_1123;
input n_701;
input n_271;
input n_995;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_984;
input n_394;
input n_79;
input n_1000;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_988;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_1035;
input n_760;
input n_1157;
input n_751;
input n_806;
input n_1127;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_1156;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;
input n_1050;

output n_6672;

wire n_4557;
wire n_6210;
wire n_5285;
wire n_6516;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_4983;
wire n_3548;
wire n_5647;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_6537;
wire n_3319;
wire n_3915;
wire n_5002;
wire n_5155;
wire n_5130;
wire n_4204;
wire n_5899;
wire n_6259;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_5827;
wire n_4805;
wire n_1765;
wire n_2392;
wire n_5008;
wire n_6183;
wire n_3280;
wire n_6616;
wire n_4371;
wire n_4601;
wire n_6035;
wire n_5858;
wire n_5879;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_6567;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_3570;
wire n_5760;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_2506;
wire n_6229;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_6639;
wire n_1730;
wire n_5243;
wire n_3479;
wire n_5587;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_5667;
wire n_2343;
wire n_5615;
wire n_1480;
wire n_6327;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_6256;
wire n_4423;
wire n_5517;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_5962;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_6658;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_6286;
wire n_3472;
wire n_5922;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_5931;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_6159;
wire n_6517;
wire n_4801;
wire n_6005;
wire n_3639;
wire n_5809;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_5588;
wire n_4569;
wire n_5404;
wire n_3671;
wire n_1778;
wire n_2839;
wire n_4998;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_5505;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_6530;
wire n_4510;
wire n_5658;
wire n_4567;
wire n_5151;
wire n_2362;
wire n_5478;
wire n_2822;
wire n_1306;
wire n_5994;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_6602;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_5037;
wire n_5878;
wire n_5716;
wire n_1960;
wire n_6562;
wire n_3979;
wire n_3714;
wire n_6534;
wire n_6629;
wire n_2844;
wire n_6192;
wire n_3565;
wire n_5304;
wire n_3883;
wire n_5866;
wire n_5941;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_5882;
wire n_1316;
wire n_1562;
wire n_6102;
wire n_4854;
wire n_3769;
wire n_6456;
wire n_1445;
wire n_6026;
wire n_2147;
wire n_5591;
wire n_6083;
wire n_2253;
wire n_4479;
wire n_5381;
wire n_3858;
wire n_4173;
wire n_6486;
wire n_5261;
wire n_5895;
wire n_5944;
wire n_6328;
wire n_5673;
wire n_4422;
wire n_5743;
wire n_1865;
wire n_5033;
wire n_6491;
wire n_4842;
wire n_4786;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_6219;
wire n_5075;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_6241;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_3780;
wire n_5571;
wire n_1653;
wire n_1375;
wire n_6254;
wire n_6066;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_5241;
wire n_3060;
wire n_5129;
wire n_4124;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_5191;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_2412;
wire n_2783;
wire n_5259;
wire n_3293;
wire n_2550;
wire n_5913;
wire n_6302;
wire n_6580;
wire n_5266;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_5580;
wire n_6078;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_5660;
wire n_5955;
wire n_1209;
wire n_5419;
wire n_3732;
wire n_6070;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_6625;
wire n_2389;
wire n_5612;
wire n_6408;
wire n_6638;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_2782;
wire n_4258;
wire n_4290;
wire n_1549;
wire n_1531;
wire n_2919;
wire n_6019;
wire n_4577;
wire n_1424;
wire n_2444;
wire n_2625;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_6485;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_5987;
wire n_6421;
wire n_6009;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_6114;
wire n_4823;
wire n_5195;
wire n_5541;
wire n_6081;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_5609;
wire n_5904;
wire n_4757;
wire n_5254;
wire n_6334;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_5423;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_6606;
wire n_1504;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_5732;
wire n_5141;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_6178;
wire n_3950;
wire n_5252;
wire n_6209;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_1271;
wire n_6011;
wire n_3416;
wire n_3147;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_5238;
wire n_6533;
wire n_3859;
wire n_6540;
wire n_4489;
wire n_3455;
wire n_1591;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_1409;
wire n_2744;
wire n_3524;
wire n_6085;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_5502;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_5288;
wire n_2264;
wire n_1987;
wire n_5749;
wire n_1244;
wire n_3365;
wire n_4974;
wire n_4725;
wire n_6431;
wire n_1932;
wire n_3775;
wire n_6196;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_6377;
wire n_3300;
wire n_5920;
wire n_5969;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_1218;
wire n_4572;
wire n_5705;
wire n_4374;
wire n_6146;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_3218;
wire n_2880;
wire n_5887;
wire n_5948;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3222;
wire n_3529;
wire n_6124;
wire n_3352;
wire n_4180;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_5199;
wire n_1207;
wire n_1735;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_4199;
wire n_6061;
wire n_5099;
wire n_1210;
wire n_6136;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_1201;
wire n_5859;
wire n_1246;
wire n_5258;
wire n_4231;
wire n_6187;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_6402;
wire n_2549;
wire n_4325;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_6305;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_6128;
wire n_2361;
wire n_4128;
wire n_5213;
wire n_6469;
wire n_5354;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_1963;
wire n_1418;
wire n_2552;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_4114;
wire n_1776;
wire n_6113;
wire n_3544;
wire n_5049;
wire n_1279;
wire n_4209;
wire n_3692;
wire n_5163;
wire n_1408;
wire n_5707;
wire n_3913;
wire n_3535;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_2954;
wire n_6379;
wire n_2046;
wire n_6454;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_4424;
wire n_6570;
wire n_1465;
wire n_6071;
wire n_4674;
wire n_6450;
wire n_1232;
wire n_2715;
wire n_6270;
wire n_4679;
wire n_6065;
wire n_1345;
wire n_4456;
wire n_5574;
wire n_1590;
wire n_2133;
wire n_3553;
wire n_5081;
wire n_6332;
wire n_6345;
wire n_1471;
wire n_3441;
wire n_5385;
wire n_4559;
wire n_5336;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_5668;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_5310;
wire n_4145;
wire n_6507;
wire n_1627;
wire n_3880;
wire n_5192;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_5206;
wire n_2010;
wire n_2733;
wire n_6120;
wire n_3796;
wire n_5719;
wire n_6544;
wire n_5157;
wire n_1836;
wire n_6384;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_4894;
wire n_5892;
wire n_5216;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_4321;
wire n_5375;
wire n_2418;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_4416;
wire n_5998;
wire n_4024;
wire n_5521;
wire n_3975;
wire n_3164;
wire n_6314;
wire n_1448;
wire n_3034;
wire n_6605;
wire n_5433;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_6349;
wire n_3759;
wire n_4777;
wire n_4800;
wire n_3629;
wire n_5573;
wire n_5620;
wire n_4117;
wire n_6527;
wire n_2884;
wire n_3383;
wire n_3687;
wire n_6626;
wire n_4154;
wire n_3459;
wire n_6105;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_5330;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_2654;
wire n_5729;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_1426;
wire n_2365;
wire n_6528;
wire n_2245;
wire n_3877;
wire n_5083;
wire n_3260;
wire n_6463;
wire n_2776;
wire n_2630;
wire n_6348;
wire n_1967;
wire n_5801;
wire n_3834;
wire n_5579;
wire n_1378;
wire n_3257;
wire n_2459;
wire n_6652;
wire n_2439;
wire n_1430;
wire n_5365;
wire n_2450;
wire n_6459;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_5263;
wire n_4851;
wire n_4963;
wire n_3387;
wire n_6126;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_6115;
wire n_3428;
wire n_5959;
wire n_6282;
wire n_2427;
wire n_5017;
wire n_5938;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_5292;
wire n_2422;
wire n_6277;
wire n_5190;
wire n_1679;
wire n_2342;
wire n_5926;
wire n_2755;
wire n_6531;
wire n_2301;
wire n_1578;
wire n_2712;
wire n_5316;
wire n_4314;
wire n_6502;
wire n_2788;
wire n_2089;
wire n_1857;
wire n_1997;
wire n_3314;
wire n_5135;
wire n_1349;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_6646;
wire n_1546;
wire n_6394;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_5840;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_6439;
wire n_6084;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_4858;
wire n_1914;
wire n_3833;
wire n_5833;
wire n_3339;
wire n_3673;
wire n_5792;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_5617;
wire n_1340;
wire n_2562;
wire n_6191;
wire n_3269;
wire n_5491;
wire n_2223;
wire n_5024;
wire n_3876;
wire n_4971;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_5696;
wire n_1816;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_6044;
wire n_4339;
wire n_5493;
wire n_4085;
wire n_3190;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_5406;
wire n_1754;
wire n_3686;
wire n_6595;
wire n_2679;
wire n_4028;
wire n_5704;
wire n_1517;
wire n_5973;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_5555;
wire n_1895;
wire n_1860;
wire n_5727;
wire n_5770;
wire n_1763;
wire n_3912;
wire n_5169;
wire n_1607;
wire n_2959;
wire n_2380;
wire n_2420;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_5274;
wire n_2516;
wire n_2031;
wire n_1348;
wire n_1191;
wire n_4099;
wire n_3899;
wire n_6153;
wire n_4729;
wire n_5957;
wire n_1617;
wire n_2639;
wire n_5323;
wire n_3099;
wire n_6412;
wire n_4745;
wire n_4057;
wire n_2410;
wire n_3206;
wire n_2633;
wire n_2049;
wire n_6245;
wire n_2113;
wire n_1690;
wire n_6553;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_6543;
wire n_5566;
wire n_6185;
wire n_5342;
wire n_4603;
wire n_4300;
wire n_3277;
wire n_2758;
wire n_5787;
wire n_4417;
wire n_5967;
wire n_1550;
wire n_1169;
wire n_6224;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_5843;
wire n_2194;
wire n_6072;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_1901;
wire n_5332;
wire n_6073;
wire n_3096;
wire n_6097;
wire n_1278;
wire n_2059;
wire n_5553;
wire n_4730;
wire n_5763;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_1603;
wire n_5864;
wire n_5227;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_5352;
wire n_4583;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_5370;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_4282;
wire n_5600;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_3650;
wire n_5014;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_6591;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_5824;
wire n_6280;
wire n_5472;
wire n_5950;
wire n_3739;
wire n_2825;
wire n_4338;
wire n_5546;
wire n_6222;
wire n_5972;
wire n_4985;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_5924;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_6656;
wire n_2366;
wire n_6318;
wire n_6200;
wire n_4919;
wire n_4200;
wire n_4111;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_4803;
wire n_1878;
wire n_1374;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_6637;
wire n_4666;
wire n_5752;
wire n_1242;
wire n_2810;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_5233;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_5977;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_5968;
wire n_2871;
wire n_2764;
wire n_5713;
wire n_3648;
wire n_3234;
wire n_6577;
wire n_4058;
wire n_6268;
wire n_5403;
wire n_4611;
wire n_5527;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_5831;
wire n_1459;
wire n_4032;
wire n_6032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_5048;
wire n_5671;
wire n_6129;
wire n_1303;
wire n_1994;
wire n_6058;
wire n_1526;
wire n_4268;
wire n_3236;
wire n_2367;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_5834;
wire n_1257;
wire n_6641;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_5951;
wire n_4895;
wire n_5480;
wire n_3354;
wire n_4069;
wire n_5289;
wire n_3373;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_6556;
wire n_4778;
wire n_4789;
wire n_2703;
wire n_6152;
wire n_2574;
wire n_5492;
wire n_1887;
wire n_6106;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_5260;
wire n_6416;
wire n_5069;
wire n_2364;
wire n_2641;
wire n_4751;
wire n_5930;
wire n_5309;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_5782;
wire n_2228;
wire n_4474;
wire n_5646;
wire n_1518;
wire n_4350;
wire n_5327;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_2266;
wire n_4473;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_5927;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_5019;
wire n_4891;
wire n_2394;
wire n_1572;
wire n_1245;
wire n_4867;
wire n_2929;
wire n_6346;
wire n_4911;
wire n_5414;
wire n_1329;
wire n_2409;
wire n_6403;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_6172;
wire n_3742;
wire n_6004;
wire n_3532;
wire n_6347;
wire n_6482;
wire n_5280;
wire n_5466;
wire n_5469;
wire n_6483;
wire n_4686;
wire n_6358;
wire n_4682;
wire n_5750;
wire n_5305;
wire n_2914;
wire n_1833;
wire n_6598;
wire n_5186;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_6499;
wire n_6215;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_3700;
wire n_5180;
wire n_6594;
wire n_6233;
wire n_4733;
wire n_5368;
wire n_6338;
wire n_5757;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_6621;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_6053;
wire n_2734;
wire n_1166;
wire n_5267;
wire n_6020;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_6432;
wire n_6426;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4797;
wire n_4962;
wire n_5397;
wire n_2596;
wire n_1488;
wire n_1379;
wire n_2972;
wire n_1721;
wire n_3606;
wire n_5232;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_5890;
wire n_4644;
wire n_4412;
wire n_6068;
wire n_5802;
wire n_4266;
wire n_5815;
wire n_5605;
wire n_2982;
wire n_2634;
wire n_3124;
wire n_5384;
wire n_6550;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_5664;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_5863;
wire n_1230;
wire n_3622;
wire n_5276;
wire n_3857;
wire n_6042;
wire n_2357;
wire n_5197;
wire n_4354;
wire n_5320;
wire n_2937;
wire n_3728;
wire n_5087;
wire n_5265;
wire n_4401;
wire n_4727;
wire n_6265;
wire n_4296;
wire n_5312;
wire n_5534;
wire n_2967;
wire n_3005;
wire n_4627;
wire n_5107;
wire n_4309;
wire n_4027;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_6452;
wire n_2802;
wire n_4728;
wire n_2279;
wire n_1536;
wire n_1719;
wire n_5281;
wire n_4046;
wire n_2961;
wire n_6458;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_1736;
wire n_6176;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_6092;
wire n_3675;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_5025;
wire n_4539;
wire n_1205;
wire n_5575;
wire n_2969;
wire n_6052;
wire n_5753;
wire n_3550;
wire n_5401;
wire n_5509;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_6468;
wire n_1414;
wire n_5506;
wire n_6063;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_5417;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_5015;
wire n_5372;
wire n_1675;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_6418;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_3662;
wire n_6344;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_5995;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_5253;
wire n_3789;
wire n_6308;
wire n_2174;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_6662;
wire n_6461;
wire n_1674;
wire n_6304;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_6617;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_5937;
wire n_2978;
wire n_5291;
wire n_3502;
wire n_5460;
wire n_3935;
wire n_5379;
wire n_1854;
wire n_2804;
wire n_5390;
wire n_5691;
wire n_4926;
wire n_5043;
wire n_6549;
wire n_4688;
wire n_5097;
wire n_5675;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_6179;
wire n_1930;
wire n_5577;
wire n_1234;
wire n_4881;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_3255;
wire n_1652;
wire n_2183;
wire n_6607;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_5181;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_5745;
wire n_4421;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_5893;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_5067;
wire n_3904;
wire n_4378;
wire n_6455;
wire n_3729;
wire n_5637;
wire n_3484;
wire n_2485;
wire n_5614;
wire n_4477;
wire n_5177;
wire n_5643;
wire n_2179;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_5695;
wire n_3726;
wire n_5438;
wire n_4277;
wire n_4431;
wire n_4771;
wire n_4652;
wire n_4970;
wire n_5179;
wire n_3804;
wire n_1908;
wire n_6457;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_5683;
wire n_3566;
wire n_6564;
wire n_2820;
wire n_2311;
wire n_5701;
wire n_4403;
wire n_3242;
wire n_6566;
wire n_1654;
wire n_6428;
wire n_5774;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_2537;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_4437;
wire n_3856;
wire n_6496;
wire n_5394;
wire n_1292;
wire n_5462;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_5428;
wire n_4491;
wire n_4672;
wire n_5001;
wire n_2421;
wire n_3237;
wire n_6095;
wire n_1970;
wire n_3946;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_6150;
wire n_3926;
wire n_3688;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_4267;
wire n_5933;
wire n_4723;
wire n_2269;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_5874;
wire n_5104;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_5964;
wire n_5551;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_5319;
wire n_5543;
wire n_4721;
wire n_2663;
wire n_3882;
wire n_2595;
wire n_5723;
wire n_5621;
wire n_5386;
wire n_4433;
wire n_5133;
wire n_5056;
wire n_3030;
wire n_5631;
wire n_5983;
wire n_5796;
wire n_4503;
wire n_6232;
wire n_3917;
wire n_3679;
wire n_4517;
wire n_6021;
wire n_3221;
wire n_3210;
wire n_4511;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_5405;
wire n_6389;
wire n_3795;
wire n_6055;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_5848;
wire n_5221;
wire n_1301;
wire n_5997;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_5122;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_5439;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_6351;
wire n_4610;
wire n_6441;
wire n_5854;
wire n_4067;
wire n_4997;
wire n_5906;
wire n_4393;
wire n_5205;
wire n_3777;
wire n_5916;
wire n_5993;
wire n_4553;
wire n_5240;
wire n_3961;
wire n_1520;
wire n_2509;
wire n_5714;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_6476;
wire n_5828;
wire n_6276;
wire n_5907;
wire n_5284;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_6669;
wire n_5357;
wire n_4994;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_6040;
wire n_2257;
wire n_4856;
wire n_5088;
wire n_5250;
wire n_1467;
wire n_6388;
wire n_3217;
wire n_2511;
wire n_5461;
wire n_6298;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_3573;
wire n_3563;
wire n_4993;
wire n_3510;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_5958;
wire n_5619;
wire n_1709;
wire n_6655;
wire n_6541;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_6460;
wire n_3241;
wire n_2746;
wire n_5471;
wire n_2256;
wire n_5210;
wire n_2445;
wire n_1980;
wire n_3583;
wire n_4987;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_6295;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_4992;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_5273;
wire n_4177;
wire n_1888;
wire n_6497;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_5877;
wire n_6535;
wire n_5457;
wire n_5482;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_6090;
wire n_3720;
wire n_1196;
wire n_1182;
wire n_4074;
wire n_5237;
wire n_5360;
wire n_3633;
wire n_1731;
wire n_5596;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_5625;
wire n_4037;
wire n_4582;
wire n_5539;
wire n_3426;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_3448;
wire n_3788;
wire n_6164;
wire n_6211;
wire n_2076;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_6117;
wire n_6563;
wire n_1312;
wire n_5844;
wire n_6470;
wire n_6448;
wire n_3684;
wire n_6667;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_6018;
wire n_6094;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_4973;
wire n_2829;
wire n_4966;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_5362;
wire n_6236;
wire n_6208;
wire n_5294;
wire n_6197;
wire n_3263;
wire n_4501;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_6552;
wire n_1421;
wire n_4922;
wire n_6237;
wire n_5089;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_2390;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_6653;
wire n_3098;
wire n_6449;
wire n_1711;
wire n_3069;
wire n_5465;
wire n_3107;
wire n_5488;
wire n_4134;
wire n_4131;
wire n_6539;
wire n_4330;
wire n_5832;
wire n_2176;
wire n_2805;
wire n_5165;
wire n_2319;
wire n_5678;
wire n_3757;
wire n_5811;
wire n_1933;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_5234;
wire n_3787;
wire n_5140;
wire n_3445;
wire n_2080;
wire n_5655;
wire n_5514;
wire n_2554;
wire n_6130;
wire n_1676;
wire n_5020;
wire n_5225;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_4462;
wire n_6560;
wire n_2787;
wire n_4540;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_4979;
wire n_3503;
wire n_2441;
wire n_4063;
wire n_4362;
wire n_5318;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_5946;
wire n_6131;
wire n_3394;
wire n_6207;
wire n_5942;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_4965;
wire n_1522;
wire n_2523;
wire n_6326;
wire n_3488;
wire n_6365;
wire n_2832;
wire n_4991;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_5242;
wire n_2142;
wire n_6519;
wire n_3703;
wire n_5116;
wire n_6635;
wire n_4554;
wire n_1260;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_6155;
wire n_5953;
wire n_2600;
wire n_3952;
wire n_1171;
wire n_6151;
wire n_6074;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_4734;
wire n_5947;
wire n_6661;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_6370;
wire n_1729;
wire n_5563;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_5194;
wire n_4579;
wire n_5628;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_6262;
wire n_2398;
wire n_1593;
wire n_1775;
wire n_6361;
wire n_2570;
wire n_4025;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_2469;
wire n_6024;
wire n_3074;
wire n_4640;
wire n_5790;
wire n_6523;
wire n_5746;
wire n_5883;
wire n_5630;
wire n_3136;
wire n_3108;
wire n_2395;
wire n_6062;
wire n_4059;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_4878;
wire n_3718;
wire n_1832;
wire n_2376;
wire n_3398;
wire n_6252;
wire n_5193;
wire n_2170;
wire n_6407;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_5153;
wire n_6235;
wire n_5369;
wire n_3238;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_5007;
wire n_4717;
wire n_4052;
wire n_6447;
wire n_2463;
wire n_6434;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_3378;
wire n_5689;
wire n_3350;
wire n_6391;
wire n_5399;
wire n_4873;
wire n_6630;
wire n_6631;
wire n_3936;
wire n_1560;
wire n_5513;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_5891;
wire n_1925;
wire n_6489;
wire n_1251;
wire n_6657;
wire n_3090;
wire n_1247;
wire n_5030;
wire n_3816;
wire n_5755;
wire n_5098;
wire n_4636;
wire n_5408;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_2765;
wire n_4278;
wire n_6165;
wire n_6263;
wire n_6481;
wire n_4609;
wire n_5148;
wire n_4822;
wire n_2936;
wire n_2985;
wire n_3106;
wire n_6597;
wire n_4030;
wire n_4276;
wire n_6238;
wire n_4612;
wire n_1667;
wire n_6272;
wire n_5454;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_5650;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_5656;
wire n_6647;
wire n_2584;
wire n_4381;
wire n_5183;
wire n_2442;
wire n_5072;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_5146;
wire n_5131;
wire n_1894;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_4699;
wire n_5803;
wire n_1331;
wire n_1223;
wire n_5754;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_5018;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_2238;
wire n_4924;
wire n_6398;
wire n_5786;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_6366;
wire n_1294;
wire n_1351;
wire n_5035;
wire n_5425;
wire n_1380;
wire n_6036;
wire n_3336;
wire n_6104;
wire n_1291;
wire n_5742;
wire n_5901;
wire n_3763;
wire n_4284;
wire n_5943;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_6253;
wire n_1830;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_5499;
wire n_1662;
wire n_3443;
wire n_5143;
wire n_3029;
wire n_4135;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_5302;
wire n_1660;
wire n_5640;
wire n_4000;
wire n_5841;
wire n_5011;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_6242;
wire n_6660;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_6414;
wire n_1962;
wire n_5296;
wire n_5159;
wire n_1952;
wire n_1624;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_2075;
wire n_4816;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_6029;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_5798;
wire n_2309;
wire n_2274;
wire n_6278;
wire n_5096;
wire n_6480;
wire n_6443;
wire n_3712;
wire n_5805;
wire n_5171;
wire n_2143;
wire n_4637;
wire n_4976;
wire n_4021;
wire n_5351;
wire n_2739;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_6157;
wire n_6453;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_4855;
wire n_5851;
wire n_4643;
wire n_5217;
wire n_6030;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_5767;
wire n_4287;
wire n_2809;
wire n_6615;
wire n_3921;
wire n_3480;
wire n_1494;
wire n_2060;
wire n_2214;
wire n_1726;
wire n_5751;
wire n_1241;
wire n_5929;
wire n_2589;
wire n_5928;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_5862;
wire n_5869;
wire n_1238;
wire n_3959;
wire n_4288;
wire n_2452;
wire n_6274;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_5201;
wire n_1644;
wire n_4586;
wire n_6190;
wire n_3860;
wire n_5353;
wire n_1871;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2818;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_5444;
wire n_4905;
wire n_6100;
wire n_1457;
wire n_3172;
wire n_2159;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_3637;
wire n_3393;
wire n_5772;
wire n_1261;
wire n_5520;
wire n_3327;
wire n_5277;
wire n_5900;
wire n_3647;
wire n_6240;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_1956;
wire n_5779;
wire n_5569;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_6498;
wire n_1669;
wire n_6247;
wire n_5109;
wire n_1885;
wire n_1989;
wire n_5837;
wire n_5402;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_4344;
wire n_1342;
wire n_6574;
wire n_2756;
wire n_4408;
wire n_1175;
wire n_5473;
wire n_1221;
wire n_3875;
wire n_5113;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2567;
wire n_5645;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_5102;
wire n_6258;
wire n_6139;
wire n_5167;
wire n_4565;
wire n_5562;
wire n_1451;
wire n_4663;
wire n_2471;
wire n_5666;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_1622;
wire n_2757;
wire n_3121;
wire n_2121;
wire n_4515;
wire n_1893;
wire n_5639;
wire n_5607;
wire n_2278;
wire n_2433;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_6169;
wire n_1507;
wire n_5914;
wire n_1206;
wire n_3576;
wire n_5275;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_2130;
wire n_4862;
wire n_5114;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_3122;
wire n_3012;
wire n_5005;
wire n_5004;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_4597;
wire n_1812;
wire n_5090;
wire n_4574;
wire n_4242;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_3820;
wire n_5395;
wire n_6494;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_5489;
wire n_2316;
wire n_5649;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2911;
wire n_1828;
wire n_1389;
wire n_6380;
wire n_5791;
wire n_1798;
wire n_5559;
wire n_4562;
wire n_1584;
wire n_5009;
wire n_6034;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_6526;
wire n_4986;
wire n_4453;
wire n_1366;
wire n_1187;
wire n_3173;
wire n_6212;
wire n_4281;
wire n_4332;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_6111;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_5295;
wire n_6427;
wire n_4310;
wire n_3752;
wire n_2637;
wire n_5047;
wire n_5504;
wire n_5076;
wire n_3543;
wire n_5693;
wire n_3655;
wire n_3791;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_6520;
wire n_4906;
wire n_4257;
wire n_5712;
wire n_4516;
wire n_2913;
wire n_5028;
wire n_2254;
wire n_1381;
wire n_1597;
wire n_1486;
wire n_6444;
wire n_5622;
wire n_4196;
wire n_5255;
wire n_2371;
wire n_6362;
wire n_3898;
wire n_3366;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_6648;
wire n_2408;
wire n_4961;
wire n_6330;
wire n_5013;
wire n_2140;
wire n_6622;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_5348;
wire n_6405;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_5251;
wire n_5036;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_6488;
wire n_4342;
wire n_5554;
wire n_2671;
wire n_3296;
wire n_5919;
wire n_5978;
wire n_6220;
wire n_1390;
wire n_2775;
wire n_3223;
wire n_2005;
wire n_2811;
wire n_1758;
wire n_2848;
wire n_6087;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_5702;
wire n_3207;
wire n_5450;
wire n_5806;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_5071;
wire n_5308;
wire n_5982;
wire n_6590;
wire n_3036;
wire n_5012;
wire n_5376;
wire n_6501;
wire n_5778;
wire n_4207;
wire n_1760;
wire n_5208;
wire n_6396;
wire n_2173;
wire n_2824;
wire n_4038;
wire n_5503;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_3046;
wire n_6551;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_5644;
wire n_6368;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_4532;
wire n_5235;
wire n_5062;
wire n_6309;
wire n_3332;
wire n_5161;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_5016;
wire n_2702;
wire n_3922;
wire n_2791;
wire n_1450;
wire n_2092;
wire n_6248;
wire n_5996;
wire n_3189;
wire n_2797;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_4442;
wire n_5700;
wire n_2168;
wire n_1442;
wire n_4689;
wire n_2886;
wire n_5699;
wire n_6287;
wire n_6022;
wire n_1968;
wire n_6579;
wire n_4018;
wire n_2609;
wire n_6633;
wire n_4613;
wire n_5940;
wire n_6614;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_3261;
wire n_5324;
wire n_6547;
wire n_5421;
wire n_3861;
wire n_5175;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_5820;
wire n_3463;
wire n_2559;
wire n_6589;
wire n_4188;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_5340;
wire n_3738;
wire n_1640;
wire n_5694;
wire n_5022;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_6297;
wire n_5245;
wire n_5651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_6367;
wire n_6198;
wire n_1355;
wire n_5364;
wire n_5459;
wire n_4534;
wire n_3635;
wire n_3270;
wire n_5168;
wire n_4590;
wire n_4602;
wire n_5510;
wire n_5329;
wire n_6251;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_6583;
wire n_3418;
wire n_2614;
wire n_5581;
wire n_1780;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_5812;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_3482;
wire n_2282;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_5711;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_3615;
wire n_5970;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_5570;
wire n_1743;
wire n_6310;
wire n_1506;
wire n_5061;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_5550;
wire n_4773;
wire n_3853;
wire n_2512;
wire n_4449;
wire n_5219;
wire n_6618;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_5132;
wire n_4883;
wire n_6249;
wire n_3559;
wire n_5184;
wire n_6440;
wire n_5747;
wire n_6575;
wire n_4943;
wire n_5821;
wire n_2498;
wire n_4630;
wire n_3812;
wire n_6584;
wire n_2017;
wire n_1227;
wire n_5326;
wire n_3750;
wire n_5909;
wire n_6050;
wire n_3838;
wire n_5868;
wire n_1954;
wire n_4749;
wire n_2687;
wire n_3456;
wire n_6643;
wire n_6569;
wire n_3132;
wire n_5618;
wire n_6596;
wire n_4159;
wire n_4372;
wire n_5528;
wire n_4731;
wire n_4004;
wire n_1684;
wire n_4353;
wire n_5593;
wire n_3334;
wire n_3819;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_5740;
wire n_1233;
wire n_5108;
wire n_3653;
wire n_4360;
wire n_6123;
wire n_4897;
wire n_2139;
wire n_3693;
wire n_5477;
wire n_5934;
wire n_5218;
wire n_2943;
wire n_5272;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_6273;
wire n_5464;
wire n_6548;
wire n_6420;
wire n_6474;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_5688;
wire n_6141;
wire n_1829;
wire n_1338;
wire n_6234;
wire n_1327;
wire n_5204;
wire n_5400;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_6311;
wire n_2565;
wire n_4201;
wire n_6634;
wire n_6288;
wire n_1636;
wire n_1687;
wire n_5303;
wire n_4584;
wire n_3184;
wire n_6290;
wire n_5804;
wire n_4155;
wire n_3890;
wire n_5519;
wire n_5023;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_1258;
wire n_2208;
wire n_1344;
wire n_5971;
wire n_2198;
wire n_1929;
wire n_5095;
wire n_1680;
wire n_1195;
wire n_5902;
wire n_4304;
wire n_4821;
wire n_4975;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_5064;
wire n_6478;
wire n_3641;
wire n_5203;
wire n_5065;
wire n_4887;
wire n_5436;
wire n_3996;
wire n_6056;
wire n_2873;
wire n_1576;
wire n_6466;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_5314;
wire n_5044;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_6228;
wire n_1841;
wire n_5886;
wire n_2685;
wire n_5344;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_5173;
wire n_5585;
wire n_3722;
wire n_5981;
wire n_3802;
wire n_5343;
wire n_5783;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_5515;
wire n_4806;
wire n_2116;
wire n_5784;
wire n_5337;
wire n_3592;
wire n_5545;
wire n_1645;
wire n_3186;
wire n_6393;
wire n_6375;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_5209;
wire n_1269;
wire n_2773;
wire n_2906;
wire n_3097;
wire n_5495;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_6424;
wire n_3822;
wire n_1276;
wire n_1637;
wire n_2900;
wire n_5799;
wire n_6296;
wire n_3765;
wire n_2216;
wire n_5888;
wire n_4259;
wire n_1620;
wire n_5196;
wire n_5086;
wire n_6025;
wire n_6168;
wire n_3518;
wire n_5885;
wire n_2022;
wire n_3967;
wire n_2373;
wire n_2275;
wire n_1853;
wire n_5398;
wire n_5434;
wire n_5797;
wire n_2899;
wire n_5830;
wire n_5896;
wire n_3351;
wire n_2008;
wire n_5052;
wire n_2859;
wire n_5952;
wire n_6003;
wire n_2564;
wire n_5110;
wire n_5918;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_5808;
wire n_6119;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_5212;
wire n_6525;
wire n_1764;
wire n_1250;
wire n_1190;
wire n_5733;
wire n_4598;
wire n_3259;
wire n_5483;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_3779;
wire n_3203;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_5278;
wire n_2114;
wire n_6204;
wire n_1609;
wire n_5522;
wire n_3530;
wire n_5584;
wire n_4548;
wire n_1803;
wire n_5264;
wire n_6321;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_6337;
wire n_4999;
wire n_5328;
wire n_2660;
wire n_5447;
wire n_5029;
wire n_5127;
wire n_5006;
wire n_5679;
wire n_4604;
wire n_5123;
wire n_6160;
wire n_3467;
wire n_6156;
wire n_4240;
wire n_2219;
wire n_6116;
wire n_4522;
wire n_1387;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_6267;
wire n_2539;
wire n_1701;
wire n_5236;
wire n_5239;
wire n_5307;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_6561;
wire n_2529;
wire n_4103;
wire n_4126;
wire n_4710;
wire n_5576;
wire n_3282;
wire n_5144;
wire n_2708;
wire n_5164;
wire n_6557;
wire n_2748;
wire n_5359;
wire n_6503;
wire n_5925;
wire n_2224;
wire n_5526;
wire n_5810;
wire n_2233;
wire n_2499;
wire n_6333;
wire n_5172;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_5126;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_5999;
wire n_5147;
wire n_5407;
wire n_1553;
wire n_3542;
wire n_5536;
wire n_6002;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_6140;
wire n_5903;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_6336;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_5849;
wire n_6663;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_2101;
wire n_5378;
wire n_3626;
wire n_2599;
wire n_4571;
wire n_5389;
wire n_6166;
wire n_3171;
wire n_6170;
wire n_1733;
wire n_6257;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_6620;
wire n_4930;
wire n_5345;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_5138;
wire n_3153;
wire n_6202;
wire n_1189;
wire n_4995;
wire n_6529;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_3232;
wire n_5228;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_5629;
wire n_5945;
wire n_4205;
wire n_6161;
wire n_3790;
wire n_6147;
wire n_2404;
wire n_5601;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_6554;
wire n_3640;
wire n_2821;
wire n_4768;
wire n_6133;
wire n_6109;
wire n_6585;
wire n_5985;
wire n_5665;
wire n_5435;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_6436;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_2063;
wire n_3082;
wire n_5709;
wire n_4504;
wire n_5176;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_5003;
wire n_2852;
wire n_2132;
wire n_5567;
wire n_1236;
wire n_3412;
wire n_5765;
wire n_1712;
wire n_6409;
wire n_4537;
wire n_5771;
wire n_5271;
wire n_1184;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_5068;
wire n_4184;
wire n_2468;
wire n_5078;
wire n_3248;
wire n_2606;
wire n_5980;
wire n_4826;
wire n_4337;
wire n_2152;
wire n_5073;
wire n_5420;
wire n_6386;
wire n_5599;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_5508;
wire n_2779;
wire n_2547;
wire n_6473;
wire n_1748;
wire n_2935;
wire n_5084;
wire n_6651;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_3568;
wire n_5789;
wire n_4876;
wire n_5322;
wire n_6490;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_6558;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_2300;
wire n_6500;
wire n_5590;
wire n_5638;
wire n_4747;
wire n_5152;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_5497;
wire n_2481;
wire n_4409;
wire n_5361;
wire n_1264;
wire n_2808;
wire n_5010;
wire n_6363;
wire n_3396;
wire n_6007;
wire n_2102;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_5117;
wire n_2977;
wire n_1682;
wire n_6142;
wire n_3599;
wire n_6244;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_6369;
wire n_6518;
wire n_5050;
wire n_5608;
wire n_5610;
wire n_4152;
wire n_1352;
wire n_5125;
wire n_2328;
wire n_6578;
wire n_4587;
wire n_6118;
wire n_6429;
wire n_6158;
wire n_2332;
wire n_1628;
wire n_1773;
wire n_3580;
wire n_2369;
wire n_5474;
wire n_3584;
wire n_4500;
wire n_5845;
wire n_1395;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_6049;
wire n_2419;
wire n_6671;
wire n_5794;
wire n_5299;
wire n_2807;
wire n_4047;
wire n_5905;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_5202;
wire n_5170;
wire n_5724;
wire n_6610;
wire n_1523;
wire n_1756;
wire n_6108;
wire n_2241;
wire n_2458;
wire n_3032;
wire n_3401;
wire n_5042;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_6382;
wire n_5662;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_6576;
wire n_1875;
wire n_1615;
wire n_3719;
wire n_5334;
wire n_5595;
wire n_6260;
wire n_5244;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_5692;
wire n_2908;
wire n_4561;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_5728;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_6148;
wire n_6404;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_6217;
wire n_6324;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_2903;
wire n_3659;
wire n_5795;
wire n_4496;
wire n_6048;
wire n_1528;
wire n_3840;
wire n_5889;
wire n_5856;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_5722;
wire n_2464;
wire n_1413;
wire n_5498;
wire n_2925;
wire n_2270;
wire n_5034;
wire n_5725;
wire n_1706;
wire n_1592;
wire n_6110;
wire n_1461;
wire n_2695;
wire n_6300;
wire n_5657;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_5282;
wire n_5511;
wire n_2414;
wire n_5736;
wire n_5642;
wire n_6624;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_4175;
wire n_4458;
wire n_6001;
wire n_3955;
wire n_3158;
wire n_3657;
wire n_5776;
wire n_5826;
wire n_2684;
wire n_2205;
wire n_2875;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_5932;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_6088;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_6239;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_6091;
wire n_4316;
wire n_5453;
wire n_3328;
wire n_2763;
wire n_5136;
wire n_6352;
wire n_2761;
wire n_4020;
wire n_5494;
wire n_6101;
wire n_1920;
wire n_4306;
wire n_6319;
wire n_2997;
wire n_3735;
wire n_2127;
wire n_6188;
wire n_5718;
wire n_5634;
wire n_3028;
wire n_3228;
wire n_5079;
wire n_3706;
wire n_6395;
wire n_1432;
wire n_3322;
wire n_1174;
wire n_6037;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_3784;
wire n_4142;
wire n_6206;
wire n_4621;
wire n_3016;
wire n_1629;
wire n_5706;
wire n_2694;
wire n_6177;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_5496;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_4007;
wire n_3960;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_5606;
wire n_6322;
wire n_1225;
wire n_2346;
wire n_4695;
wire n_2180;
wire n_3376;
wire n_6313;
wire n_5989;
wire n_2617;
wire n_5870;
wire n_4163;
wire n_2831;
wire n_6504;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_5530;
wire n_4498;
wire n_2240;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_5424;
wire n_5230;
wire n_2086;
wire n_4832;
wire n_5229;
wire n_3666;
wire n_6374;
wire n_1839;
wire n_5160;
wire n_2555;
wire n_2330;
wire n_1587;
wire n_6356;
wire n_6640;
wire n_5313;
wire n_2108;
wire n_6462;
wire n_5333;
wire n_5207;
wire n_2535;
wire n_5158;
wire n_2945;
wire n_5154;
wire n_3057;
wire n_4319;
wire n_3760;
wire n_5721;
wire n_1396;
wire n_1923;
wire n_1224;
wire n_5654;
wire n_2196;
wire n_5860;
wire n_1538;
wire n_3773;
wire n_5884;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_2437;
wire n_2351;
wire n_1889;
wire n_5839;
wire n_2688;
wire n_4990;
wire n_3302;
wire n_1673;
wire n_5058;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_6231;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_3645;
wire n_5823;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_6401;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_6521;
wire n_4849;
wire n_5101;
wire n_5532;
wire n_4366;
wire n_6582;
wire n_4139;
wire n_1270;
wire n_5297;
wire n_4340;
wire n_1476;
wire n_2027;
wire n_5611;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_6623;
wire n_1880;
wire n_6225;
wire n_1642;
wire n_5744;
wire n_2447;
wire n_3358;
wire n_5538;
wire n_2894;
wire n_5249;
wire n_5669;
wire n_2587;
wire n_1605;
wire n_6134;
wire n_2099;
wire n_1202;
wire n_5793;
wire n_3410;
wire n_4900;
wire n_6493;
wire n_6364;
wire n_5715;
wire n_6665;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_5966;
wire n_2299;
wire n_2078;
wire n_6284;
wire n_3709;
wire n_3011;
wire n_5383;
wire n_6649;
wire n_5775;
wire n_2315;
wire n_3623;
wire n_6230;
wire n_5558;
wire n_2157;
wire n_6546;
wire n_3446;
wire n_5547;
wire n_5572;
wire n_5659;
wire n_5223;
wire n_6555;
wire n_1770;
wire n_4167;
wire n_6010;
wire n_3058;
wire n_4334;
wire n_6331;
wire n_2211;
wire n_6047;
wire n_5708;
wire n_6532;
wire n_5817;
wire n_3384;
wire n_4698;
wire n_2225;
wire n_1411;
wire n_5867;
wire n_1501;
wire n_5636;
wire n_5106;
wire n_5800;
wire n_5257;
wire n_4397;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_5371;
wire n_6524;
wire n_4229;
wire n_4294;
wire n_1919;
wire n_4351;
wire n_6226;
wire n_2893;
wire n_6281;
wire n_2009;
wire n_6514;
wire n_5731;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_3871;
wire n_2388;
wire n_3112;
wire n_5623;
wire n_5921;
wire n_6082;
wire n_3413;
wire n_4580;
wire n_2624;
wire n_1813;
wire n_4581;
wire n_4618;
wire n_5178;
wire n_6609;
wire n_5853;
wire n_5898;
wire n_5198;
wire n_2898;
wire n_5437;
wire n_6627;
wire n_2519;
wire n_2231;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_5053;
wire n_1256;
wire n_4670;
wire n_6162;
wire n_5592;
wire n_5484;
wire n_6650;
wire n_4982;
wire n_5418;
wire n_6079;
wire n_6013;
wire n_5432;
wire n_1769;
wire n_5270;
wire n_1372;
wire n_1847;
wire n_5166;
wire n_5358;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_1586;
wire n_3497;
wire n_5156;
wire n_6592;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_5548;
wire n_5687;
wire n_3561;
wire n_2543;
wire n_6512;
wire n_2992;
wire n_1541;
wire n_6008;
wire n_6522;
wire n_4907;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_5822;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_5758;
wire n_1939;
wire n_5366;
wire n_4053;
wire n_5392;
wire n_4279;
wire n_3937;
wire n_6400;
wire n_3303;
wire n_5115;
wire n_5046;
wire n_5139;
wire n_4555;
wire n_5829;
wire n_5686;
wire n_5735;
wire n_3549;
wire n_1481;
wire n_6613;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_5674;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1361;
wire n_5039;
wire n_6538;
wire n_1693;
wire n_2081;
wire n_5341;
wire n_2993;
wire n_5032;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_5041;
wire n_6505;
wire n_3989;
wire n_6581;
wire n_5565;
wire n_6350;
wire n_4752;
wire n_4546;
wire n_3918;
wire n_6378;
wire n_3191;
wire n_3051;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_4415;
wire n_2487;
wire n_3343;
wire n_3163;
wire n_6243;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_6484;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_6573;
wire n_6419;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_5448;
wire n_4263;
wire n_3725;
wire n_5974;
wire n_5852;
wire n_6143;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_5085;
wire n_4335;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_6112;
wire n_6138;
wire n_3009;
wire n_4471;
wire n_3297;
wire n_1168;
wire n_5500;
wire n_6045;
wire n_5293;
wire n_6203;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_6568;
wire n_4547;
wire n_4836;
wire n_5458;
wire n_3545;
wire n_4193;
wire n_5670;
wire n_1336;
wire n_6433;
wire n_6023;
wire n_1358;
wire n_3318;
wire n_5684;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_4984;
wire n_1532;
wire n_5624;
wire n_3430;
wire n_1685;
wire n_5325;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_6167;
wire n_6189;
wire n_5059;
wire n_1462;
wire n_5825;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_5586;
wire n_1398;
wire n_5222;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_6335;
wire n_5741;
wire n_1692;
wire n_5875;
wire n_4796;
wire n_6312;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_5045;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_6611;
wire n_5038;
wire n_5769;
wire n_3837;
wire n_4841;
wire n_6213;
wire n_3076;
wire n_6264;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_5703;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2653;
wire n_2855;
wire n_6301;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_5501;
wire n_6216;
wire n_2331;
wire n_1600;
wire n_5894;
wire n_4701;
wire n_5248;
wire n_5872;
wire n_4088;
wire n_2136;
wire n_5443;
wire n_6193;
wire n_1913;
wire n_3056;
wire n_4208;
wire n_5363;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_6588;
wire n_4589;
wire n_3924;
wire n_1915;
wire n_2534;
wire n_5908;
wire n_4972;
wire n_5597;
wire n_4617;
wire n_3311;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_3613;
wire n_1383;
wire n_2057;
wire n_5984;
wire n_6385;
wire n_5533;
wire n_1822;
wire n_6051;
wire n_1804;
wire n_1581;
wire n_5387;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_1851;
wire n_1755;
wire n_5589;
wire n_4702;
wire n_1341;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_5380;
wire n_2262;
wire n_5134;
wire n_1333;
wire n_4506;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_6015;
wire n_4329;
wire n_6435;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_6411;
wire n_4327;
wire n_5954;
wire n_5412;
wire n_2656;
wire n_6323;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_5174;
wire n_4465;
wire n_6174;
wire n_2544;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_5468;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_4075;
wire n_5429;
wire n_3593;
wire n_6586;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_5269;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_3768;
wire n_4224;
wire n_4868;
wire n_5124;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_3181;
wire n_3644;
wire n_5287;
wire n_4387;
wire n_5865;
wire n_2368;
wire n_6437;
wire n_4896;
wire n_2065;
wire n_2901;
wire n_5583;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_4798;
wire n_2201;
wire n_1582;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_3610;
wire n_5416;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_5373;
wire n_4967;
wire n_6067;
wire n_5377;
wire n_2290;
wire n_6479;
wire n_3272;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_5350;
wire n_6279;
wire n_4668;
wire n_2383;
wire n_5632;
wire n_2640;
wire n_1492;
wire n_6425;
wire n_1478;
wire n_1796;
wire n_3569;
wire n_2374;
wire n_1614;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_5290;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_5120;
wire n_2230;
wire n_5535;
wire n_3033;
wire n_2151;
wire n_5382;
wire n_6354;
wire n_4912;
wire n_6320;
wire n_1971;
wire n_5759;
wire n_2479;
wire n_4914;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_6612;
wire n_6376;
wire n_2571;
wire n_5479;
wire n_6006;
wire n_5598;
wire n_6132;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_5578;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_6089;
wire n_5211;
wire n_1668;
wire n_5861;
wire n_6417;
wire n_1681;
wire n_4031;
wire n_4120;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_5092;
wire n_1945;
wire n_5182;
wire n_5430;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_4840;
wire n_2354;
wire n_5956;
wire n_6027;
wire n_6477;
wire n_4311;
wire n_5766;
wire n_6269;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_5094;
wire n_6275;
wire n_3264;
wire n_3204;
wire n_6390;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_6306;
wire n_3881;
wire n_1910;
wire n_5446;
wire n_1606;
wire n_5315;
wire n_3711;
wire n_2164;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_6122;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_6175;
wire n_5279;
wire n_6506;
wire n_4650;
wire n_6415;
wire n_2280;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_3809;
wire n_1999;
wire n_3810;
wire n_5103;
wire n_5835;
wire n_4968;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_5311;
wire n_2283;
wire n_2806;
wire n_6184;
wire n_2813;
wire n_5268;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_6285;
wire n_5773;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_5451;
wire n_5452;
wire n_2145;
wire n_2122;
wire n_6644;
wire n_1588;
wire n_2579;
wire n_2876;
wire n_6670;
wire n_3301;
wire n_2370;
wire n_5321;
wire n_5215;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_4513;
wire n_5635;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_5356;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_5150;
wire n_2826;
wire n_2112;
wire n_6180;
wire n_5613;
wire n_6137;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_6410;
wire n_5063;
wire n_4671;
wire n_1326;
wire n_6046;
wire n_4981;
wire n_1799;
wire n_1689;
wire n_1304;
wire n_6465;
wire n_5653;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_5788;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_2722;
wire n_5057;
wire n_3618;
wire n_2727;
wire n_5560;
wire n_2719;
wire n_2213;
wire n_5476;
wire n_3521;
wire n_6121;
wire n_2723;
wire n_6077;
wire n_4054;
wire n_1569;
wire n_6000;
wire n_6205;
wire n_4012;
wire n_5582;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_5935;
wire n_6201;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_5697;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_5119;
wire n_2292;
wire n_6471;
wire n_3560;
wire n_5813;
wire n_1742;
wire n_1818;
wire n_5100;
wire n_3847;
wire n_2203;
wire n_5427;
wire n_4909;
wire n_2693;
wire n_2281;
wire n_3202;
wire n_5467;
wire n_2646;
wire n_5346;
wire n_3887;
wire n_3800;
wire n_4435;
wire n_1235;
wire n_6329;
wire n_4755;
wire n_6355;
wire n_3827;
wire n_6145;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_5633;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_5726;
wire n_2890;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_5415;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_5445;
wire n_6446;
wire n_4996;
wire n_4136;
wire n_5040;
wire n_4358;
wire n_2857;
wire n_5031;
wire n_1360;
wire n_5814;
wire n_5374;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_4156;
wire n_3754;
wire n_6057;
wire n_5818;
wire n_2416;
wire n_2962;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_6221;
wire n_5876;
wire n_5529;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_5317;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_5490;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_5897;
wire n_5331;
wire n_6107;
wire n_4655;
wire n_6080;
wire n_1634;
wire n_5556;
wire n_1452;
wire n_4953;
wire n_6339;
wire n_4570;
wire n_5391;
wire n_5431;
wire n_3966;
wire n_4293;
wire n_6371;
wire n_6014;
wire n_1577;
wire n_1700;
wire n_4122;
wire n_4542;
wire n_5021;
wire n_2819;
wire n_5456;
wire n_5523;
wire n_1985;
wire n_4740;
wire n_3007;
wire n_1487;
wire n_6373;
wire n_1237;
wire n_4230;
wire n_2741;
wire n_4333;
wire n_5231;
wire n_5512;
wire n_6406;
wire n_3436;
wire n_6223;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_1884;
wire n_6632;
wire n_2717;
wire n_1589;
wire n_5720;
wire n_4527;
wire n_2877;
wire n_5881;
wire n_1996;
wire n_5857;
wire n_5256;
wire n_3964;
wire n_3110;
wire n_5717;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_1792;
wire n_6654;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_5561;
wire n_1877;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_5487;
wire n_4407;
wire n_5961;
wire n_5077;
wire n_5214;
wire n_1249;
wire n_3468;
wire n_2006;
wire n_1990;
wire n_5413;
wire n_3680;
wire n_6227;
wire n_3624;
wire n_6098;
wire n_4989;
wire n_2467;
wire n_5066;
wire n_4292;
wire n_3145;
wire n_5682;
wire n_2662;
wire n_3872;
wire n_5602;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_6163;
wire n_1464;
wire n_1566;
wire n_6565;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_6601;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_2999;
wire n_3331;
wire n_2910;
wire n_4414;
wire n_2294;
wire n_2295;
wire n_4977;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_6076;
wire n_5347;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_3554;
wire n_6199;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_1935;
wire n_5568;
wire n_3367;
wire n_2785;
wire n_5060;
wire n_4929;
wire n_5121;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_5756;
wire n_5162;
wire n_5224;
wire n_2160;
wire n_2991;
wire n_2699;
wire n_6513;
wire n_6214;
wire n_1436;
wire n_4137;
wire n_1485;
wire n_2239;
wire n_6289;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_4215;
wire n_4315;
wire n_6559;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3797;
wire n_3281;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2934;
wire n_6430;
wire n_4042;
wire n_5663;
wire n_2525;
wire n_5552;
wire n_4624;
wire n_6043;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_5672;
wire n_4958;
wire n_5051;
wire n_4297;
wire n_5367;
wire n_5339;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_5000;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_3646;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_5226;
wire n_2095;
wire n_2486;
wire n_5819;
wire n_5855;
wire n_2521;
wire n_5388;
wire n_1574;
wire n_6608;
wire n_6186;
wire n_4764;
wire n_4899;
wire n_6283;
wire n_6445;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_6372;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_3167;
wire n_5188;
wire n_2986;
wire n_4969;
wire n_2400;
wire n_6467;
wire n_6144;
wire n_5681;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_6291;
wire n_1357;
wire n_6593;
wire n_4566;
wire n_5262;
wire n_2794;
wire n_6542;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_5604;
wire n_2990;
wire n_2923;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_5910;
wire n_1315;
wire n_4647;
wire n_2340;
wire n_6125;
wire n_2117;
wire n_5990;
wire n_1328;
wire n_4837;
wire n_6218;
wire n_3638;
wire n_2106;
wire n_5880;
wire n_5685;
wire n_6515;
wire n_6619;
wire n_6060;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_6664;
wire n_5992;
wire n_5105;
wire n_5807;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_5449;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_6599;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_2524;
wire n_3927;
wire n_1941;
wire n_5338;
wire n_5070;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_5842;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_6173;
wire n_4133;
wire n_6093;
wire n_3985;
wire n_6099;
wire n_5939;
wire n_5481;
wire n_5187;
wire n_5762;
wire n_3252;
wire n_2578;
wire n_5486;
wire n_5426;
wire n_2745;
wire n_2110;
wire n_6031;
wire n_6064;
wire n_3747;
wire n_1323;
wire n_5846;
wire n_6033;
wire n_3710;
wire n_1429;
wire n_6316;
wire n_3209;
wire n_2026;
wire n_5537;
wire n_3588;
wire n_5220;
wire n_6341;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_3632;
wire n_5200;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_5816;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1458;
wire n_1694;
wire n_2271;
wire n_2356;
wire n_5676;
wire n_5463;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_4980;
wire n_2187;
wire n_2105;
wire n_5780;
wire n_2642;
wire n_5485;
wire n_5737;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_6571;
wire n_2384;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_6039;
wire n_5355;
wire n_4048;
wire n_4084;
wire n_5149;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_5185;
wire n_2849;
wire n_6509;
wire n_6642;
wire n_5847;
wire n_5091;
wire n_5936;
wire n_1177;
wire n_3292;
wire n_6442;
wire n_6636;
wire n_3940;
wire n_6475;
wire n_2502;
wire n_5396;
wire n_4860;
wire n_4438;
wire n_5300;
wire n_3290;
wire n_3585;
wire n_2878;
wire n_1810;
wire n_6342;
wire n_3047;
wire n_2610;
wire n_5917;
wire n_5306;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_2698;
wire n_3930;
wire n_4149;
wire n_5518;
wire n_5531;
wire n_1259;
wire n_4101;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_6012;
wire n_4383;
wire n_2709;
wire n_5074;
wire n_6492;
wire n_2244;
wire n_6387;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_5246;
wire n_2665;
wire n_5544;
wire n_3063;
wire n_4543;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_5652;
wire n_5409;
wire n_2581;
wire n_6271;
wire n_5540;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_2255;
wire n_1820;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_6149;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_2153;
wire n_5777;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_6545;
wire n_4434;
wire n_2737;
wire n_5557;
wire n_1406;
wire n_3591;
wire n_6054;
wire n_2137;
wire n_5442;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_5549;
wire n_3139;
wire n_4715;
wire n_6250;
wire n_4222;
wire n_5730;
wire n_2206;
wire n_3734;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_5054;
wire n_5349;
wire n_1167;
wire n_3231;
wire n_6423;
wire n_6659;
wire n_3138;
wire n_6303;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_4988;
wire n_5128;
wire n_3454;
wire n_6668;
wire n_6299;
wire n_4143;
wire n_5027;
wire n_4410;
wire n_5026;
wire n_5189;
wire n_1718;
wire n_3229;
wire n_2546;
wire n_4741;
wire n_6383;
wire n_5516;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_3649;
wire n_1838;
wire n_3824;
wire n_3439;
wire n_5525;
wire n_1513;
wire n_5836;
wire n_5677;
wire n_6182;
wire n_6510;
wire n_1788;
wire n_5764;
wire n_2348;
wire n_6171;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_5768;
wire n_6353;
wire n_6472;
wire n_2248;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_6360;
wire n_3846;
wire n_4328;
wire n_5142;
wire n_1433;
wire n_5082;
wire n_1907;
wire n_3994;
wire n_5911;
wire n_5118;
wire n_2135;
wire n_5781;
wire n_5739;
wire n_6666;
wire n_6075;
wire n_5145;
wire n_4487;
wire n_5111;
wire n_4148;
wire n_3066;
wire n_6135;
wire n_2869;
wire n_6422;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_6266;
wire n_5748;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_5734;
wire n_2667;
wire n_6317;
wire n_6059;
wire n_5247;
wire n_1565;
wire n_2325;
wire n_6041;
wire n_3346;
wire n_5411;
wire n_5422;
wire n_3391;
wire n_1542;
wire n_1547;
wire n_5991;
wire n_1362;
wire n_6343;
wire n_4178;
wire n_4324;
wire n_3288;
wire n_2518;
wire n_6069;
wire n_3045;
wire n_3014;
wire n_5475;
wire n_6511;
wire n_1951;
wire n_1330;
wire n_5850;
wire n_6307;
wire n_5440;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_5641;
wire n_1861;
wire n_1564;
wire n_2593;
wire n_1623;
wire n_6413;
wire n_6603;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_6255;
wire n_4761;
wire n_6294;
wire n_2021;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_3342;
wire n_5441;
wire n_2939;
wire n_6587;
wire n_4036;
wire n_5055;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_6487;
wire n_1892;
wire n_5761;
wire n_6195;
wire n_2061;
wire n_6038;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_5976;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_5871;
wire n_2827;
wire n_5680;
wire n_3278;
wire n_2701;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_6086;
wire n_5915;
wire n_5524;
wire n_5112;
wire n_3042;
wire n_5542;
wire n_5627;
wire n_2561;
wire n_5785;
wire n_2491;
wire n_6438;
wire n_5298;
wire n_4363;
wire n_5564;
wire n_5603;
wire n_3551;
wire n_3992;
wire n_4147;
wire n_6451;
wire n_4811;
wire n_6495;
wire n_5093;
wire n_5710;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_5986;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_5137;
wire n_1759;
wire n_2096;
wire n_5912;
wire n_2296;
wire n_6194;
wire n_1911;
wire n_6381;
wire n_2870;
wire n_4869;
wire n_6397;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_6628;
wire n_5283;
wire n_1419;
wire n_4738;
wire n_6604;
wire n_1193;
wire n_2928;
wire n_3380;
wire n_3557;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_5286;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_5626;
wire n_4086;
wire n_5410;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_3286;
wire n_2668;
wire n_1386;
wire n_2931;
wire n_2492;
wire n_5960;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_5988;
wire n_1499;
wire n_5838;
wire n_2155;
wire n_3938;
wire n_6103;
wire n_6016;
wire n_3114;
wire n_3905;
wire n_1661;
wire n_6261;
wire n_1965;
wire n_5616;
wire n_1757;
wire n_6399;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_6181;
wire n_3053;
wire n_5965;
wire n_3894;
wire n_6645;
wire n_2407;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2453;
wire n_2560;
wire n_6572;
wire n_4544;
wire n_4418;
wire n_4595;
wire n_2770;
wire n_2704;
wire n_6246;
wire n_1762;
wire n_4944;
wire n_4468;
wire n_5923;
wire n_6357;
wire n_6508;
wire n_6536;
wire n_3421;
wire n_4950;
wire n_3247;
wire n_1454;
wire n_4108;
wire n_4594;
wire n_6359;
wire n_5949;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_5738;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_6096;
wire n_4921;
wire n_1819;
wire n_4863;
wire n_2670;
wire n_1745;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_5080;
wire n_5975;
wire n_1791;
wire n_5301;
wire n_6464;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_6017;
wire n_5507;
wire n_6340;
wire n_3749;
wire n_5470;
wire n_6315;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_6392;
wire n_4280;
wire n_2285;
wire n_5979;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_5648;
wire n_1665;
wire n_5335;
wire n_5594;
wire n_3417;
wire n_2725;
wire n_1482;
wire n_4782;
wire n_5393;
wire n_5661;
wire n_4978;
wire n_6292;
wire n_5690;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_6154;
wire n_5963;
wire n_6293;
wire n_1417;
wire n_5455;
wire n_3536;
wire n_1346;
wire n_5873;
wire n_2834;
wire n_6127;
wire n_1272;
wire n_2497;
wire n_3040;
wire n_6028;
wire n_6325;
wire n_1410;
wire n_6600;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_2743;
wire n_5698;
wire n_4662;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_941),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_946),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_1025),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_666),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_331),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_744),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_1072),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_882),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_28),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_165),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_678),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_742),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_167),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_463),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_291),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_544),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_831),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_799),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_841),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_514),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_906),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1133),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_210),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_44),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_627),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_821),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_519),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1061),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1129),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_752),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1038),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_38),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1088),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_398),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1124),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_362),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1026),
.Y(n_1202)
);

CKINVDCx14_ASAP7_75t_R g1203 ( 
.A(n_1105),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_649),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1035),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_622),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_814),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_314),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_664),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_128),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_619),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_416),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1090),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_882),
.Y(n_1214)
);

INVx1_ASAP7_75t_SL g1215 ( 
.A(n_400),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_579),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1130),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_80),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_1070),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1139),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_951),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_71),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_59),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1089),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_157),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_142),
.Y(n_1226)
);

CKINVDCx20_ASAP7_75t_R g1227 ( 
.A(n_96),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_899),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_1092),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_391),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_771),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_1111),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_164),
.Y(n_1233)
);

CKINVDCx16_ASAP7_75t_R g1234 ( 
.A(n_381),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1058),
.Y(n_1235)
);

CKINVDCx16_ASAP7_75t_R g1236 ( 
.A(n_145),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1021),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_581),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_592),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_390),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_991),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_573),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_403),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_381),
.Y(n_1244)
);

INVxp67_ASAP7_75t_L g1245 ( 
.A(n_129),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_676),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_736),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1123),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1094),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_1139),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_442),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_186),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_380),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_164),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1151),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1163),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_472),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_524),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_648),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_639),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_100),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_542),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_952),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1116),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1118),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_399),
.Y(n_1266)
);

CKINVDCx20_ASAP7_75t_R g1267 ( 
.A(n_1165),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_479),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_309),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1027),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_35),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_812),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_232),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_308),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_932),
.Y(n_1275)
);

INVxp67_ASAP7_75t_L g1276 ( 
.A(n_220),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_305),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_231),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_1114),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_511),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_416),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_13),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_1000),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_564),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_781),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_463),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_246),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_15),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_692),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_907),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_927),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_503),
.Y(n_1292)
);

INVx1_ASAP7_75t_SL g1293 ( 
.A(n_1095),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_289),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1082),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_941),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_736),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_812),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_443),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1135),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_726),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1005),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_72),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_255),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_741),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_449),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_767),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_992),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_732),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_279),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_26),
.Y(n_1311)
);

BUFx10_ASAP7_75t_L g1312 ( 
.A(n_896),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_514),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_745),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_8),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_1140),
.Y(n_1316)
);

INVx1_ASAP7_75t_SL g1317 ( 
.A(n_295),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_53),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_412),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_177),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_165),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_55),
.Y(n_1322)
);

BUFx3_ASAP7_75t_L g1323 ( 
.A(n_195),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_297),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_998),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_855),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1135),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1075),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1151),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_30),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_787),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_711),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_853),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_222),
.Y(n_1334)
);

INVxp67_ASAP7_75t_SL g1335 ( 
.A(n_228),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_605),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1066),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_648),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_758),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_799),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_671),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_679),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_836),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_739),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_535),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_804),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_151),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_317),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1098),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_317),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_595),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_423),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1117),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_889),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_177),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_984),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_45),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_756),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_540),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_996),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_177),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_166),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_216),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_353),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1136),
.Y(n_1365)
);

INVx1_ASAP7_75t_SL g1366 ( 
.A(n_649),
.Y(n_1366)
);

CKINVDCx14_ASAP7_75t_R g1367 ( 
.A(n_231),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1021),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_307),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1091),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_891),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_123),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_530),
.Y(n_1373)
);

BUFx10_ASAP7_75t_L g1374 ( 
.A(n_1048),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_995),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_184),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_103),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_183),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1104),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1107),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_846),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_84),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1096),
.Y(n_1383)
);

BUFx2_ASAP7_75t_SL g1384 ( 
.A(n_1099),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_364),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_919),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_238),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_315),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_328),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_696),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_738),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_382),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_432),
.Y(n_1393)
);

CKINVDCx20_ASAP7_75t_R g1394 ( 
.A(n_13),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_734),
.Y(n_1395)
);

CKINVDCx20_ASAP7_75t_R g1396 ( 
.A(n_1031),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_49),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1077),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1108),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_236),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_453),
.Y(n_1401)
);

INVx1_ASAP7_75t_SL g1402 ( 
.A(n_412),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_994),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_962),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_993),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_398),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_143),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_377),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_5),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_297),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1067),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1137),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_428),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_968),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_564),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_887),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_872),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1028),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1161),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_109),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_984),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_843),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_733),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_167),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_735),
.Y(n_1425)
);

CKINVDCx16_ASAP7_75t_R g1426 ( 
.A(n_520),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1128),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1138),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_661),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_207),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1006),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_228),
.Y(n_1432)
);

BUFx10_ASAP7_75t_L g1433 ( 
.A(n_810),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_932),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_107),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1010),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_200),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_213),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_911),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_647),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_949),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_635),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_225),
.Y(n_1443)
);

INVx1_ASAP7_75t_SL g1444 ( 
.A(n_985),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1091),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_952),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1159),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1079),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_909),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_317),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_453),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_481),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_682),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_60),
.Y(n_1454)
);

CKINVDCx20_ASAP7_75t_R g1455 ( 
.A(n_55),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_315),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_687),
.Y(n_1457)
);

CKINVDCx20_ASAP7_75t_R g1458 ( 
.A(n_183),
.Y(n_1458)
);

CKINVDCx20_ASAP7_75t_R g1459 ( 
.A(n_935),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_900),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1112),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_332),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_689),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_979),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1120),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_180),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_1110),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_492),
.Y(n_1468)
);

BUFx3_ASAP7_75t_L g1469 ( 
.A(n_446),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_729),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_285),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_673),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_1159),
.Y(n_1473)
);

CKINVDCx20_ASAP7_75t_R g1474 ( 
.A(n_233),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_555),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_895),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_423),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_439),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1004),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_112),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1109),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_233),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_283),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_10),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_674),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_9),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_761),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_957),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1121),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_499),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1132),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_698),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_927),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_183),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_74),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_587),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_3),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1028),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_469),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_885),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_593),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_674),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1083),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_154),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_692),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_337),
.Y(n_1506)
);

BUFx10_ASAP7_75t_L g1507 ( 
.A(n_909),
.Y(n_1507)
);

BUFx6f_ASAP7_75t_L g1508 ( 
.A(n_128),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_99),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_684),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_489),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1093),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1157),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_197),
.Y(n_1514)
);

BUFx8_ASAP7_75t_SL g1515 ( 
.A(n_48),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_37),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_834),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_222),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_789),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_289),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_9),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_10),
.Y(n_1522)
);

CKINVDCx16_ASAP7_75t_R g1523 ( 
.A(n_1053),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_988),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_208),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_628),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_415),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_454),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_448),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_792),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_925),
.Y(n_1531)
);

BUFx10_ASAP7_75t_L g1532 ( 
.A(n_399),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1104),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_616),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_657),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_942),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_932),
.Y(n_1537)
);

BUFx10_ASAP7_75t_L g1538 ( 
.A(n_117),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_719),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1088),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_782),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_34),
.Y(n_1542)
);

INVx1_ASAP7_75t_SL g1543 ( 
.A(n_564),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_963),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_1115),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_635),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_803),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1081),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_323),
.Y(n_1549)
);

BUFx8_ASAP7_75t_SL g1550 ( 
.A(n_953),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1089),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_911),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_318),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_864),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_969),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1125),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_206),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_179),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_257),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1078),
.Y(n_1560)
);

CKINVDCx20_ASAP7_75t_R g1561 ( 
.A(n_304),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1146),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1074),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_62),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_719),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_880),
.Y(n_1566)
);

BUFx10_ASAP7_75t_L g1567 ( 
.A(n_362),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_622),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_77),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_392),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_637),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_705),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1087),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_910),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_537),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_670),
.Y(n_1576)
);

CKINVDCx20_ASAP7_75t_R g1577 ( 
.A(n_141),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_555),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_387),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_133),
.Y(n_1580)
);

BUFx5_ASAP7_75t_L g1581 ( 
.A(n_465),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1128),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_555),
.Y(n_1583)
);

BUFx5_ASAP7_75t_L g1584 ( 
.A(n_980),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_405),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_692),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_629),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1133),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_556),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_917),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_345),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_703),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1026),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_388),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_571),
.Y(n_1595)
);

BUFx6f_ASAP7_75t_L g1596 ( 
.A(n_526),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1141),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_129),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1074),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_184),
.Y(n_1600)
);

CKINVDCx14_ASAP7_75t_R g1601 ( 
.A(n_25),
.Y(n_1601)
);

INVx2_ASAP7_75t_SL g1602 ( 
.A(n_1116),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_92),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_380),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_233),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_412),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_837),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_140),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1085),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_886),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_562),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_408),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_283),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_865),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_513),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_55),
.Y(n_1616)
);

BUFx6f_ASAP7_75t_L g1617 ( 
.A(n_199),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_359),
.Y(n_1618)
);

CKINVDCx16_ASAP7_75t_R g1619 ( 
.A(n_105),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_612),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_638),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_422),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1103),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1065),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_1084),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_727),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_347),
.Y(n_1627)
);

INVx1_ASAP7_75t_SL g1628 ( 
.A(n_678),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_717),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_913),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_452),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1097),
.Y(n_1632)
);

CKINVDCx20_ASAP7_75t_R g1633 ( 
.A(n_948),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_179),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_713),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_559),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_235),
.Y(n_1637)
);

CKINVDCx16_ASAP7_75t_R g1638 ( 
.A(n_1121),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1154),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_71),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_660),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_714),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_707),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_338),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1101),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_629),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_253),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_915),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_966),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_987),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_173),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_619),
.Y(n_1652)
);

CKINVDCx20_ASAP7_75t_R g1653 ( 
.A(n_341),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_69),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_838),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_1100),
.Y(n_1656)
);

BUFx10_ASAP7_75t_L g1657 ( 
.A(n_312),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_181),
.Y(n_1658)
);

BUFx10_ASAP7_75t_L g1659 ( 
.A(n_1053),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_62),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_755),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1106),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1127),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_253),
.Y(n_1664)
);

CKINVDCx20_ASAP7_75t_R g1665 ( 
.A(n_940),
.Y(n_1665)
);

INVxp67_ASAP7_75t_L g1666 ( 
.A(n_781),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_457),
.Y(n_1667)
);

CKINVDCx20_ASAP7_75t_R g1668 ( 
.A(n_1099),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_526),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_784),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_324),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_529),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_631),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_559),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1165),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_885),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_237),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_764),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_221),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_742),
.Y(n_1680)
);

BUFx3_ASAP7_75t_L g1681 ( 
.A(n_225),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_563),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_174),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_268),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_299),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_1067),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_640),
.Y(n_1687)
);

BUFx6f_ASAP7_75t_L g1688 ( 
.A(n_995),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_207),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_678),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_556),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_82),
.Y(n_1692)
);

CKINVDCx16_ASAP7_75t_R g1693 ( 
.A(n_1128),
.Y(n_1693)
);

INVxp67_ASAP7_75t_L g1694 ( 
.A(n_488),
.Y(n_1694)
);

INVx2_ASAP7_75t_SL g1695 ( 
.A(n_1003),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_873),
.Y(n_1696)
);

BUFx2_ASAP7_75t_L g1697 ( 
.A(n_1156),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_148),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_944),
.Y(n_1699)
);

BUFx3_ASAP7_75t_L g1700 ( 
.A(n_748),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_348),
.Y(n_1701)
);

INVx2_ASAP7_75t_SL g1702 ( 
.A(n_1064),
.Y(n_1702)
);

BUFx3_ASAP7_75t_L g1703 ( 
.A(n_326),
.Y(n_1703)
);

CKINVDCx20_ASAP7_75t_R g1704 ( 
.A(n_834),
.Y(n_1704)
);

BUFx3_ASAP7_75t_L g1705 ( 
.A(n_127),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_233),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_1019),
.Y(n_1707)
);

CKINVDCx20_ASAP7_75t_R g1708 ( 
.A(n_108),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_195),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_148),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_560),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_516),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_872),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_288),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_138),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_314),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_713),
.Y(n_1717)
);

INVxp67_ASAP7_75t_SL g1718 ( 
.A(n_194),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1113),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_0),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_471),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_633),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_1022),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_754),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_902),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1119),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_511),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_543),
.Y(n_1728)
);

CKINVDCx20_ASAP7_75t_R g1729 ( 
.A(n_1052),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_991),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_1046),
.Y(n_1731)
);

BUFx6f_ASAP7_75t_L g1732 ( 
.A(n_878),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_1126),
.Y(n_1733)
);

INVx1_ASAP7_75t_SL g1734 ( 
.A(n_619),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_467),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_223),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1102),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_385),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_625),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_346),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_880),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_378),
.Y(n_1742)
);

CKINVDCx20_ASAP7_75t_R g1743 ( 
.A(n_1073),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_592),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_209),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_174),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_569),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_1016),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_231),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_181),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_419),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_290),
.Y(n_1752)
);

CKINVDCx20_ASAP7_75t_R g1753 ( 
.A(n_204),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_94),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1058),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_900),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1111),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_556),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_750),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_673),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_842),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_41),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_576),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_889),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_479),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_41),
.Y(n_1766)
);

CKINVDCx16_ASAP7_75t_R g1767 ( 
.A(n_220),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_463),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_671),
.Y(n_1769)
);

BUFx10_ASAP7_75t_L g1770 ( 
.A(n_123),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_1156),
.Y(n_1771)
);

CKINVDCx14_ASAP7_75t_R g1772 ( 
.A(n_1096),
.Y(n_1772)
);

BUFx10_ASAP7_75t_L g1773 ( 
.A(n_225),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_271),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_1129),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_1103),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_644),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1065),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_693),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_109),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_782),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_1051),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_935),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_803),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_158),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_431),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_1023),
.Y(n_1787)
);

BUFx10_ASAP7_75t_L g1788 ( 
.A(n_567),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_428),
.Y(n_1789)
);

INVxp33_ASAP7_75t_SL g1790 ( 
.A(n_524),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_1033),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1137),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_116),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_1135),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_802),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_320),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_380),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_345),
.Y(n_1798)
);

BUFx8_ASAP7_75t_SL g1799 ( 
.A(n_1018),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1099),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_1073),
.Y(n_1801)
);

BUFx3_ASAP7_75t_L g1802 ( 
.A(n_877),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_440),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_680),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_279),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_450),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_36),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_625),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_1063),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_595),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_632),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_323),
.Y(n_1812)
);

CKINVDCx20_ASAP7_75t_R g1813 ( 
.A(n_537),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_149),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_373),
.Y(n_1815)
);

CKINVDCx20_ASAP7_75t_R g1816 ( 
.A(n_1066),
.Y(n_1816)
);

BUFx3_ASAP7_75t_L g1817 ( 
.A(n_1134),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_85),
.Y(n_1818)
);

BUFx6f_ASAP7_75t_L g1819 ( 
.A(n_650),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_433),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_875),
.Y(n_1821)
);

CKINVDCx20_ASAP7_75t_R g1822 ( 
.A(n_293),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_239),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_814),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_738),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_774),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_846),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_888),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_451),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_1086),
.Y(n_1830)
);

BUFx6f_ASAP7_75t_L g1831 ( 
.A(n_1131),
.Y(n_1831)
);

CKINVDCx20_ASAP7_75t_R g1832 ( 
.A(n_639),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1108),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_788),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_1071),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_92),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1069),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_379),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1068),
.Y(n_1839)
);

CKINVDCx20_ASAP7_75t_R g1840 ( 
.A(n_490),
.Y(n_1840)
);

INVx1_ASAP7_75t_SL g1841 ( 
.A(n_1109),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_359),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_1080),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_469),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_206),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_827),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_690),
.Y(n_1847)
);

BUFx6f_ASAP7_75t_L g1848 ( 
.A(n_249),
.Y(n_1848)
);

INVx2_ASAP7_75t_SL g1849 ( 
.A(n_229),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_909),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_269),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_639),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1149),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_571),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_152),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_72),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1003),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_848),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_1015),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_1161),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_818),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_894),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_883),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_12),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_800),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_15),
.Y(n_1866)
);

CKINVDCx16_ASAP7_75t_R g1867 ( 
.A(n_90),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_231),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1122),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_141),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_325),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_95),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_126),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_68),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_378),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_826),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_887),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_611),
.Y(n_1878)
);

CKINVDCx20_ASAP7_75t_R g1879 ( 
.A(n_844),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_1076),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_480),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_396),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_948),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_239),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_32),
.Y(n_1885)
);

INVxp33_ASAP7_75t_L g1886 ( 
.A(n_1515),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1538),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1581),
.Y(n_1888)
);

INVxp33_ASAP7_75t_SL g1889 ( 
.A(n_1397),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1538),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_1515),
.Y(n_1891)
);

INVxp33_ASAP7_75t_L g1892 ( 
.A(n_1173),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1538),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1770),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1770),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_1367),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_1367),
.Y(n_1897)
);

INVxp67_ASAP7_75t_L g1898 ( 
.A(n_1323),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1770),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1773),
.Y(n_1900)
);

INVxp33_ASAP7_75t_L g1901 ( 
.A(n_1761),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1773),
.Y(n_1902)
);

INVxp33_ASAP7_75t_SL g1903 ( 
.A(n_1828),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_1601),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1773),
.Y(n_1905)
);

CKINVDCx20_ASAP7_75t_R g1906 ( 
.A(n_1601),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1175),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1178),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1210),
.Y(n_1909)
);

CKINVDCx14_ASAP7_75t_R g1910 ( 
.A(n_1203),
.Y(n_1910)
);

BUFx2_ASAP7_75t_L g1911 ( 
.A(n_1223),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1252),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1254),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1321),
.Y(n_1914)
);

CKINVDCx20_ASAP7_75t_R g1915 ( 
.A(n_1227),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1322),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1376),
.Y(n_1917)
);

INVxp67_ASAP7_75t_L g1918 ( 
.A(n_1323),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1387),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1407),
.Y(n_1920)
);

CKINVDCx14_ASAP7_75t_R g1921 ( 
.A(n_1203),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1437),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1494),
.Y(n_1923)
);

BUFx2_ASAP7_75t_L g1924 ( 
.A(n_1223),
.Y(n_1924)
);

INVxp33_ASAP7_75t_L g1925 ( 
.A(n_1877),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1581),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1495),
.Y(n_1927)
);

INVxp33_ASAP7_75t_SL g1928 ( 
.A(n_1188),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1516),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1525),
.Y(n_1930)
);

INVxp67_ASAP7_75t_SL g1931 ( 
.A(n_1409),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1557),
.Y(n_1932)
);

INVxp33_ASAP7_75t_SL g1933 ( 
.A(n_1189),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1558),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1569),
.Y(n_1935)
);

CKINVDCx20_ASAP7_75t_R g1936 ( 
.A(n_1227),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1580),
.Y(n_1937)
);

INVxp67_ASAP7_75t_SL g1938 ( 
.A(n_1409),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1616),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1634),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1637),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1654),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_1772),
.Y(n_1943)
);

CKINVDCx20_ASAP7_75t_R g1944 ( 
.A(n_1318),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1660),
.Y(n_1945)
);

INVxp67_ASAP7_75t_SL g1946 ( 
.A(n_1484),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1698),
.Y(n_1947)
);

INVxp67_ASAP7_75t_L g1948 ( 
.A(n_1484),
.Y(n_1948)
);

INVxp33_ASAP7_75t_SL g1949 ( 
.A(n_1197),
.Y(n_1949)
);

INVxp33_ASAP7_75t_SL g1950 ( 
.A(n_1218),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1710),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1772),
.Y(n_1952)
);

BUFx3_ASAP7_75t_L g1953 ( 
.A(n_1640),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1720),
.Y(n_1954)
);

INVxp67_ASAP7_75t_SL g1955 ( 
.A(n_1640),
.Y(n_1955)
);

INVxp33_ASAP7_75t_SL g1956 ( 
.A(n_1222),
.Y(n_1956)
);

INVxp67_ASAP7_75t_L g1957 ( 
.A(n_1681),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1581),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1749),
.Y(n_1959)
);

CKINVDCx20_ASAP7_75t_R g1960 ( 
.A(n_1318),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1750),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1780),
.Y(n_1962)
);

INVxp67_ASAP7_75t_SL g1963 ( 
.A(n_1681),
.Y(n_1963)
);

CKINVDCx14_ASAP7_75t_R g1964 ( 
.A(n_1312),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1581),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1785),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1793),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1845),
.Y(n_1968)
);

INVxp67_ASAP7_75t_L g1969 ( 
.A(n_1705),
.Y(n_1969)
);

INVxp67_ASAP7_75t_SL g1970 ( 
.A(n_1705),
.Y(n_1970)
);

CKINVDCx20_ASAP7_75t_R g1971 ( 
.A(n_1394),
.Y(n_1971)
);

CKINVDCx20_ASAP7_75t_R g1972 ( 
.A(n_1394),
.Y(n_1972)
);

INVxp67_ASAP7_75t_SL g1973 ( 
.A(n_1265),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1856),
.Y(n_1974)
);

CKINVDCx20_ASAP7_75t_R g1975 ( 
.A(n_1424),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1868),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1581),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1550),
.Y(n_1978)
);

INVxp67_ASAP7_75t_SL g1979 ( 
.A(n_1265),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1872),
.Y(n_1980)
);

BUFx3_ASAP7_75t_L g1981 ( 
.A(n_1265),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1874),
.Y(n_1982)
);

BUFx2_ASAP7_75t_L g1983 ( 
.A(n_1236),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1885),
.Y(n_1984)
);

NOR2xp67_ASAP7_75t_L g1985 ( 
.A(n_1452),
.B(n_0),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1309),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1314),
.Y(n_1987)
);

CKINVDCx20_ASAP7_75t_R g1988 ( 
.A(n_1424),
.Y(n_1988)
);

NOR2xp67_ASAP7_75t_L g1989 ( 
.A(n_1452),
.B(n_0),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1697),
.Y(n_1990)
);

INVxp67_ASAP7_75t_SL g1991 ( 
.A(n_1245),
.Y(n_1991)
);

HB1xp67_ASAP7_75t_L g1992 ( 
.A(n_1619),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1602),
.Y(n_1993)
);

CKINVDCx16_ASAP7_75t_R g1994 ( 
.A(n_1767),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_1550),
.Y(n_1995)
);

INVx2_ASAP7_75t_SL g1996 ( 
.A(n_1312),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1602),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1695),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1695),
.Y(n_1999)
);

NOR2xp67_ASAP7_75t_L g2000 ( 
.A(n_1702),
.B(n_0),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1702),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1363),
.Y(n_2002)
);

INVxp33_ASAP7_75t_L g2003 ( 
.A(n_1799),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1581),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1799),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1363),
.Y(n_2006)
);

HB1xp67_ASAP7_75t_L g2007 ( 
.A(n_1867),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1849),
.Y(n_2008)
);

CKINVDCx16_ASAP7_75t_R g2009 ( 
.A(n_1234),
.Y(n_2009)
);

CKINVDCx5p33_ASAP7_75t_R g2010 ( 
.A(n_1870),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1849),
.Y(n_2011)
);

INVxp67_ASAP7_75t_SL g2012 ( 
.A(n_1276),
.Y(n_2012)
);

INVxp67_ASAP7_75t_L g2013 ( 
.A(n_1198),
.Y(n_2013)
);

CKINVDCx20_ASAP7_75t_R g2014 ( 
.A(n_1454),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1171),
.Y(n_2015)
);

INVxp67_ASAP7_75t_L g2016 ( 
.A(n_1198),
.Y(n_2016)
);

INVxp67_ASAP7_75t_L g2017 ( 
.A(n_1212),
.Y(n_2017)
);

HB1xp67_ASAP7_75t_L g2018 ( 
.A(n_1225),
.Y(n_2018)
);

CKINVDCx5p33_ASAP7_75t_R g2019 ( 
.A(n_1884),
.Y(n_2019)
);

CKINVDCx20_ASAP7_75t_R g2020 ( 
.A(n_1454),
.Y(n_2020)
);

CKINVDCx20_ASAP7_75t_R g2021 ( 
.A(n_1455),
.Y(n_2021)
);

HB1xp67_ASAP7_75t_L g2022 ( 
.A(n_1233),
.Y(n_2022)
);

INVxp67_ASAP7_75t_SL g2023 ( 
.A(n_1226),
.Y(n_2023)
);

CKINVDCx20_ASAP7_75t_R g2024 ( 
.A(n_1455),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_1261),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_1273),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_1278),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1182),
.Y(n_2028)
);

INVxp67_ASAP7_75t_SL g2029 ( 
.A(n_1226),
.Y(n_2029)
);

INVxp33_ASAP7_75t_L g2030 ( 
.A(n_1174),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1183),
.Y(n_2031)
);

CKINVDCx20_ASAP7_75t_R g2032 ( 
.A(n_1458),
.Y(n_2032)
);

CKINVDCx20_ASAP7_75t_R g2033 ( 
.A(n_1458),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1184),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1185),
.Y(n_2035)
);

CKINVDCx14_ASAP7_75t_R g2036 ( 
.A(n_1312),
.Y(n_2036)
);

INVxp33_ASAP7_75t_SL g2037 ( 
.A(n_1282),
.Y(n_2037)
);

BUFx6f_ASAP7_75t_L g2038 ( 
.A(n_1953),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1981),
.Y(n_2039)
);

BUFx6f_ASAP7_75t_L g2040 ( 
.A(n_1911),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_L g2041 ( 
.A(n_1996),
.B(n_1887),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_L g2042 ( 
.A(n_1890),
.B(n_1790),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1924),
.B(n_1288),
.Y(n_2043)
);

BUFx6f_ASAP7_75t_L g2044 ( 
.A(n_1907),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1888),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1892),
.B(n_1426),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1991),
.B(n_1303),
.Y(n_2047)
);

HB1xp67_ASAP7_75t_L g2048 ( 
.A(n_1983),
.Y(n_2048)
);

BUFx6f_ASAP7_75t_L g2049 ( 
.A(n_1908),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1938),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1938),
.Y(n_2051)
);

CKINVDCx6p67_ASAP7_75t_R g2052 ( 
.A(n_1994),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1898),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1926),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1901),
.B(n_1523),
.Y(n_2055)
);

HB1xp67_ASAP7_75t_L g2056 ( 
.A(n_1992),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1898),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1918),
.Y(n_2058)
);

OAI22x1_ASAP7_75t_L g2059 ( 
.A1(n_2007),
.A2(n_1577),
.B1(n_1708),
.B2(n_1474),
.Y(n_2059)
);

BUFx6f_ASAP7_75t_L g2060 ( 
.A(n_1909),
.Y(n_2060)
);

OA21x2_ASAP7_75t_L g2061 ( 
.A1(n_1912),
.A2(n_1382),
.B(n_1271),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_2012),
.B(n_1311),
.Y(n_2062)
);

AND2x4_ASAP7_75t_L g2063 ( 
.A(n_1986),
.B(n_1212),
.Y(n_2063)
);

BUFx6f_ASAP7_75t_L g2064 ( 
.A(n_1913),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1918),
.B(n_1315),
.Y(n_2065)
);

HB1xp67_ASAP7_75t_L g2066 ( 
.A(n_1964),
.Y(n_2066)
);

OA21x2_ASAP7_75t_L g2067 ( 
.A1(n_1914),
.A2(n_1382),
.B(n_1271),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1948),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_1987),
.B(n_1253),
.Y(n_2069)
);

INVx6_ASAP7_75t_L g2070 ( 
.A(n_2009),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_1893),
.B(n_1790),
.Y(n_2071)
);

AOI22xp5_ASAP7_75t_L g2072 ( 
.A1(n_1889),
.A2(n_1577),
.B1(n_1708),
.B2(n_1474),
.Y(n_2072)
);

BUFx2_ASAP7_75t_L g2073 ( 
.A(n_2010),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1948),
.Y(n_2074)
);

AND2x4_ASAP7_75t_L g2075 ( 
.A(n_1990),
.B(n_1253),
.Y(n_2075)
);

BUFx6f_ASAP7_75t_L g2076 ( 
.A(n_1916),
.Y(n_2076)
);

AND2x4_ASAP7_75t_L g2077 ( 
.A(n_2018),
.B(n_1337),
.Y(n_2077)
);

INVxp67_ASAP7_75t_L g2078 ( 
.A(n_2022),
.Y(n_2078)
);

BUFx8_ASAP7_75t_SL g2079 ( 
.A(n_1915),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1957),
.Y(n_2080)
);

CKINVDCx6p67_ASAP7_75t_R g2081 ( 
.A(n_1906),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1957),
.B(n_1320),
.Y(n_2082)
);

INVx2_ASAP7_75t_SL g2083 ( 
.A(n_2019),
.Y(n_2083)
);

AND2x4_ASAP7_75t_L g2084 ( 
.A(n_1894),
.B(n_1337),
.Y(n_2084)
);

BUFx6f_ASAP7_75t_L g2085 ( 
.A(n_1917),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1969),
.Y(n_2086)
);

AND2x4_ASAP7_75t_L g2087 ( 
.A(n_1895),
.B(n_1469),
.Y(n_2087)
);

NOR2x1_ASAP7_75t_L g2088 ( 
.A(n_1899),
.B(n_1469),
.Y(n_2088)
);

BUFx8_ASAP7_75t_SL g2089 ( 
.A(n_1936),
.Y(n_2089)
);

BUFx2_ASAP7_75t_L g2090 ( 
.A(n_2025),
.Y(n_2090)
);

NOR2xp33_ASAP7_75t_L g2091 ( 
.A(n_1900),
.B(n_1638),
.Y(n_2091)
);

AND2x4_ASAP7_75t_L g2092 ( 
.A(n_1902),
.B(n_1506),
.Y(n_2092)
);

AND2x4_ASAP7_75t_L g2093 ( 
.A(n_1905),
.B(n_1506),
.Y(n_2093)
);

AND2x4_ASAP7_75t_L g2094 ( 
.A(n_1896),
.B(n_1897),
.Y(n_2094)
);

AND2x4_ASAP7_75t_L g2095 ( 
.A(n_1904),
.B(n_1536),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1969),
.Y(n_2096)
);

OAI22x1_ASAP7_75t_R g2097 ( 
.A1(n_1944),
.A2(n_1232),
.B1(n_1250),
.B2(n_1228),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1931),
.Y(n_2098)
);

BUFx6f_ASAP7_75t_L g2099 ( 
.A(n_1919),
.Y(n_2099)
);

BUFx6f_ASAP7_75t_L g2100 ( 
.A(n_1920),
.Y(n_2100)
);

INVx4_ASAP7_75t_L g2101 ( 
.A(n_2026),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_1925),
.B(n_1693),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1946),
.Y(n_2103)
);

BUFx6f_ASAP7_75t_L g2104 ( 
.A(n_1922),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1955),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1958),
.Y(n_2106)
);

BUFx6f_ASAP7_75t_L g2107 ( 
.A(n_1923),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2036),
.B(n_1334),
.Y(n_2108)
);

BUFx6f_ASAP7_75t_L g2109 ( 
.A(n_1927),
.Y(n_2109)
);

INVx3_ASAP7_75t_L g2110 ( 
.A(n_1993),
.Y(n_2110)
);

INVx6_ASAP7_75t_L g2111 ( 
.A(n_1903),
.Y(n_2111)
);

OA21x2_ASAP7_75t_L g2112 ( 
.A1(n_1929),
.A2(n_1603),
.B(n_1514),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1965),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1977),
.Y(n_2114)
);

BUFx6f_ASAP7_75t_L g2115 ( 
.A(n_1930),
.Y(n_2115)
);

INVxp33_ASAP7_75t_SL g2116 ( 
.A(n_2027),
.Y(n_2116)
);

CKINVDCx5p33_ASAP7_75t_R g2117 ( 
.A(n_1928),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1963),
.Y(n_2118)
);

BUFx12f_ASAP7_75t_L g2119 ( 
.A(n_1891),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1970),
.Y(n_2120)
);

INVx4_ASAP7_75t_L g2121 ( 
.A(n_1943),
.Y(n_2121)
);

NAND2x1_ASAP7_75t_L g2122 ( 
.A(n_1932),
.B(n_1514),
.Y(n_2122)
);

BUFx6f_ASAP7_75t_L g2123 ( 
.A(n_1934),
.Y(n_2123)
);

CKINVDCx20_ASAP7_75t_R g2124 ( 
.A(n_1960),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2004),
.Y(n_2125)
);

OA21x2_ASAP7_75t_L g2126 ( 
.A1(n_1935),
.A2(n_1679),
.B(n_1603),
.Y(n_2126)
);

NOR2xp33_ASAP7_75t_L g2127 ( 
.A(n_1933),
.B(n_1666),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2013),
.B(n_1347),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1973),
.Y(n_2129)
);

HB1xp67_ASAP7_75t_L g2130 ( 
.A(n_1949),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_2002),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_2006),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_2008),
.Y(n_2133)
);

BUFx6f_ASAP7_75t_L g2134 ( 
.A(n_1937),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_2011),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_1910),
.B(n_1921),
.Y(n_2136)
);

INVx6_ASAP7_75t_L g2137 ( 
.A(n_1886),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1979),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2013),
.B(n_1357),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1997),
.Y(n_2140)
);

INVx3_ASAP7_75t_L g2141 ( 
.A(n_1998),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1999),
.Y(n_2142)
);

NOR2xp33_ASAP7_75t_L g2143 ( 
.A(n_1950),
.B(n_1694),
.Y(n_2143)
);

INVx3_ASAP7_75t_L g2144 ( 
.A(n_2001),
.Y(n_2144)
);

AND2x4_ASAP7_75t_L g2145 ( 
.A(n_1952),
.B(n_2016),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2016),
.Y(n_2146)
);

BUFx2_ASAP7_75t_L g2147 ( 
.A(n_1971),
.Y(n_2147)
);

NOR2xp33_ASAP7_75t_L g2148 ( 
.A(n_1956),
.B(n_1361),
.Y(n_2148)
);

OAI22xp5_ASAP7_75t_SL g2149 ( 
.A1(n_1972),
.A2(n_1232),
.B1(n_1250),
.B2(n_1228),
.Y(n_2149)
);

BUFx6f_ASAP7_75t_L g2150 ( 
.A(n_1939),
.Y(n_2150)
);

BUFx12f_ASAP7_75t_L g2151 ( 
.A(n_1978),
.Y(n_2151)
);

BUFx6f_ASAP7_75t_L g2152 ( 
.A(n_1940),
.Y(n_2152)
);

OAI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_2037),
.A2(n_2003),
.B1(n_1362),
.B2(n_1377),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_2015),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2017),
.Y(n_2155)
);

INVx2_ASAP7_75t_SL g2156 ( 
.A(n_2028),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2017),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_2031),
.Y(n_2158)
);

BUFx12f_ASAP7_75t_L g2159 ( 
.A(n_1995),
.Y(n_2159)
);

INVx3_ASAP7_75t_L g2160 ( 
.A(n_1941),
.Y(n_2160)
);

BUFx3_ASAP7_75t_L g2161 ( 
.A(n_1942),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2023),
.Y(n_2162)
);

BUFx6f_ASAP7_75t_L g2163 ( 
.A(n_1945),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2034),
.Y(n_2164)
);

AND2x4_ASAP7_75t_L g2165 ( 
.A(n_2035),
.B(n_2029),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1947),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1951),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1954),
.Y(n_2168)
);

BUFx8_ASAP7_75t_L g2169 ( 
.A(n_2005),
.Y(n_2169)
);

CKINVDCx6p67_ASAP7_75t_R g2170 ( 
.A(n_1975),
.Y(n_2170)
);

AND2x6_ASAP7_75t_L g2171 ( 
.A(n_1959),
.B(n_1536),
.Y(n_2171)
);

BUFx8_ASAP7_75t_L g2172 ( 
.A(n_1988),
.Y(n_2172)
);

OA21x2_ASAP7_75t_L g2173 ( 
.A1(n_1961),
.A2(n_1692),
.B(n_1679),
.Y(n_2173)
);

INVx2_ASAP7_75t_SL g2174 ( 
.A(n_1962),
.Y(n_2174)
);

BUFx3_ASAP7_75t_L g2175 ( 
.A(n_1966),
.Y(n_2175)
);

INVx3_ASAP7_75t_L g2176 ( 
.A(n_1967),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_1968),
.B(n_1374),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1974),
.Y(n_2178)
);

OAI22x1_ASAP7_75t_SL g2179 ( 
.A1(n_2014),
.A2(n_1275),
.B1(n_1279),
.B2(n_1267),
.Y(n_2179)
);

BUFx8_ASAP7_75t_L g2180 ( 
.A(n_2020),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1976),
.Y(n_2181)
);

INVx3_ASAP7_75t_L g2182 ( 
.A(n_1980),
.Y(n_2182)
);

INVxp33_ASAP7_75t_L g2183 ( 
.A(n_2021),
.Y(n_2183)
);

BUFx12f_ASAP7_75t_L g2184 ( 
.A(n_2024),
.Y(n_2184)
);

AND2x4_ASAP7_75t_L g2185 ( 
.A(n_1985),
.B(n_1555),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1982),
.Y(n_2186)
);

INVx3_ASAP7_75t_L g2187 ( 
.A(n_1984),
.Y(n_2187)
);

NOR2x1_ASAP7_75t_L g2188 ( 
.A(n_1989),
.B(n_2000),
.Y(n_2188)
);

INVx3_ASAP7_75t_L g2189 ( 
.A(n_2030),
.Y(n_2189)
);

BUFx6f_ASAP7_75t_L g2190 ( 
.A(n_2032),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2033),
.B(n_1372),
.Y(n_2191)
);

HB1xp67_ASAP7_75t_L g2192 ( 
.A(n_1911),
.Y(n_2192)
);

BUFx8_ASAP7_75t_SL g2193 ( 
.A(n_1915),
.Y(n_2193)
);

BUFx6f_ASAP7_75t_L g2194 ( 
.A(n_1953),
.Y(n_2194)
);

BUFx6f_ASAP7_75t_L g2195 ( 
.A(n_1953),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_1911),
.B(n_1378),
.Y(n_2196)
);

OAI22xp5_ASAP7_75t_SL g2197 ( 
.A1(n_1915),
.A2(n_1275),
.B1(n_1279),
.B2(n_1267),
.Y(n_2197)
);

AOI22xp5_ASAP7_75t_L g2198 ( 
.A1(n_1889),
.A2(n_1753),
.B1(n_1420),
.B2(n_1430),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1953),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1911),
.B(n_1400),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1953),
.Y(n_2201)
);

BUFx6f_ASAP7_75t_L g2202 ( 
.A(n_1953),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1981),
.Y(n_2203)
);

AND2x4_ASAP7_75t_L g2204 ( 
.A(n_1911),
.B(n_1555),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1981),
.Y(n_2205)
);

BUFx6f_ASAP7_75t_L g2206 ( 
.A(n_1953),
.Y(n_2206)
);

INVx5_ASAP7_75t_L g2207 ( 
.A(n_1996),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_1892),
.B(n_1374),
.Y(n_2208)
);

HB1xp67_ASAP7_75t_L g2209 ( 
.A(n_1911),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_1953),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1981),
.Y(n_2211)
);

BUFx6f_ASAP7_75t_L g2212 ( 
.A(n_1953),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_1911),
.B(n_1432),
.Y(n_2213)
);

NOR2xp33_ASAP7_75t_L g2214 ( 
.A(n_1996),
.B(n_1435),
.Y(n_2214)
);

AND2x4_ASAP7_75t_L g2215 ( 
.A(n_1911),
.B(n_1700),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1981),
.Y(n_2216)
);

BUFx6f_ASAP7_75t_L g2217 ( 
.A(n_1953),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1981),
.Y(n_2218)
);

OR2x2_ASAP7_75t_L g2219 ( 
.A(n_1983),
.B(n_1384),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1981),
.Y(n_2220)
);

CKINVDCx16_ASAP7_75t_R g2221 ( 
.A(n_1994),
.Y(n_2221)
);

AOI22xp5_ASAP7_75t_L g2222 ( 
.A1(n_1889),
.A2(n_1753),
.B1(n_1466),
.B2(n_1480),
.Y(n_2222)
);

INVx6_ASAP7_75t_L g2223 ( 
.A(n_1994),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1953),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_1953),
.Y(n_2225)
);

INVx6_ASAP7_75t_L g2226 ( 
.A(n_1994),
.Y(n_2226)
);

BUFx6f_ASAP7_75t_L g2227 ( 
.A(n_1953),
.Y(n_2227)
);

INVx4_ASAP7_75t_L g2228 ( 
.A(n_1911),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1981),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_1953),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1981),
.Y(n_2231)
);

OAI22xp5_ASAP7_75t_L g2232 ( 
.A1(n_1994),
.A2(n_1438),
.B1(n_1486),
.B2(n_1482),
.Y(n_2232)
);

INVxp33_ASAP7_75t_SL g2233 ( 
.A(n_1992),
.Y(n_2233)
);

INVxp67_ASAP7_75t_L g2234 ( 
.A(n_1992),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1911),
.B(n_1504),
.Y(n_2235)
);

INVx5_ASAP7_75t_L g2236 ( 
.A(n_1996),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_1892),
.B(n_1374),
.Y(n_2237)
);

OAI22xp5_ASAP7_75t_L g2238 ( 
.A1(n_1994),
.A2(n_1509),
.B1(n_1521),
.B2(n_1518),
.Y(n_2238)
);

BUFx6f_ASAP7_75t_L g2239 ( 
.A(n_1953),
.Y(n_2239)
);

BUFx8_ASAP7_75t_L g2240 ( 
.A(n_1983),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_1953),
.Y(n_2241)
);

BUFx6f_ASAP7_75t_L g2242 ( 
.A(n_1953),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_1892),
.B(n_1433),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1981),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1981),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_1953),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_1892),
.B(n_1433),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1953),
.Y(n_2248)
);

OAI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_1994),
.A2(n_1522),
.B1(n_1564),
.B2(n_1542),
.Y(n_2249)
);

BUFx6f_ASAP7_75t_L g2250 ( 
.A(n_1953),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_1892),
.B(n_1433),
.Y(n_2251)
);

BUFx2_ASAP7_75t_L g2252 ( 
.A(n_1983),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_1953),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_1892),
.B(n_1507),
.Y(n_2254)
);

NOR2xp33_ASAP7_75t_SL g2255 ( 
.A(n_1889),
.B(n_1598),
.Y(n_2255)
);

HB1xp67_ASAP7_75t_L g2256 ( 
.A(n_1911),
.Y(n_2256)
);

BUFx6f_ASAP7_75t_L g2257 ( 
.A(n_1953),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_1892),
.B(n_1507),
.Y(n_2258)
);

AND2x6_ASAP7_75t_L g2259 ( 
.A(n_1887),
.B(n_1700),
.Y(n_2259)
);

INVx3_ASAP7_75t_L g2260 ( 
.A(n_1981),
.Y(n_2260)
);

AND2x4_ASAP7_75t_L g2261 ( 
.A(n_1911),
.B(n_1703),
.Y(n_2261)
);

INVx3_ASAP7_75t_L g2262 ( 
.A(n_1981),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_1953),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1981),
.Y(n_2264)
);

BUFx6f_ASAP7_75t_L g2265 ( 
.A(n_1953),
.Y(n_2265)
);

INVx6_ASAP7_75t_L g2266 ( 
.A(n_1994),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1953),
.Y(n_2267)
);

HB1xp67_ASAP7_75t_L g2268 ( 
.A(n_1911),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_1996),
.B(n_1600),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1981),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_1953),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_1911),
.B(n_1605),
.Y(n_2272)
);

BUFx8_ASAP7_75t_L g2273 ( 
.A(n_1983),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1981),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1981),
.Y(n_2275)
);

OAI22xp5_ASAP7_75t_SL g2276 ( 
.A1(n_1915),
.A2(n_1306),
.B1(n_1351),
.B2(n_1292),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1981),
.Y(n_2277)
);

INVx4_ASAP7_75t_L g2278 ( 
.A(n_1911),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_1911),
.B(n_1608),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1981),
.Y(n_2280)
);

AND2x4_ASAP7_75t_L g2281 ( 
.A(n_1911),
.B(n_1703),
.Y(n_2281)
);

HB1xp67_ASAP7_75t_L g2282 ( 
.A(n_1911),
.Y(n_2282)
);

NOR2xp33_ASAP7_75t_L g2283 ( 
.A(n_1996),
.B(n_1651),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_1953),
.Y(n_2284)
);

CKINVDCx20_ASAP7_75t_R g2285 ( 
.A(n_2079),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2131),
.Y(n_2286)
);

CKINVDCx5p33_ASAP7_75t_R g2287 ( 
.A(n_2089),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2132),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2133),
.Y(n_2289)
);

CKINVDCx5p33_ASAP7_75t_R g2290 ( 
.A(n_2193),
.Y(n_2290)
);

CKINVDCx16_ASAP7_75t_R g2291 ( 
.A(n_2255),
.Y(n_2291)
);

HB1xp67_ASAP7_75t_L g2292 ( 
.A(n_2056),
.Y(n_2292)
);

CKINVDCx5p33_ASAP7_75t_R g2293 ( 
.A(n_2184),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_2061),
.Y(n_2294)
);

CKINVDCx20_ASAP7_75t_R g2295 ( 
.A(n_2240),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_2052),
.Y(n_2296)
);

AND2x4_ASAP7_75t_L g2297 ( 
.A(n_2177),
.B(n_1802),
.Y(n_2297)
);

CKINVDCx5p33_ASAP7_75t_R g2298 ( 
.A(n_2052),
.Y(n_2298)
);

AND2x2_ASAP7_75t_L g2299 ( 
.A(n_2046),
.B(n_1507),
.Y(n_2299)
);

NOR2xp33_ASAP7_75t_R g2300 ( 
.A(n_2117),
.B(n_1292),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2135),
.Y(n_2301)
);

CKINVDCx5p33_ASAP7_75t_R g2302 ( 
.A(n_2273),
.Y(n_2302)
);

NOR2xp33_ASAP7_75t_R g2303 ( 
.A(n_2221),
.B(n_1306),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2140),
.Y(n_2304)
);

OR2x2_ASAP7_75t_L g2305 ( 
.A(n_2252),
.B(n_1172),
.Y(n_2305)
);

BUFx6f_ASAP7_75t_SL g2306 ( 
.A(n_2101),
.Y(n_2306)
);

CKINVDCx20_ASAP7_75t_R g2307 ( 
.A(n_2124),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2067),
.Y(n_2308)
);

CKINVDCx5p33_ASAP7_75t_R g2309 ( 
.A(n_2116),
.Y(n_2309)
);

CKINVDCx20_ASAP7_75t_R g2310 ( 
.A(n_2170),
.Y(n_2310)
);

CKINVDCx20_ASAP7_75t_R g2311 ( 
.A(n_2170),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2112),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2126),
.Y(n_2313)
);

CKINVDCx5p33_ASAP7_75t_R g2314 ( 
.A(n_2172),
.Y(n_2314)
);

CKINVDCx5p33_ASAP7_75t_R g2315 ( 
.A(n_2180),
.Y(n_2315)
);

BUFx2_ASAP7_75t_L g2316 ( 
.A(n_2048),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2173),
.Y(n_2317)
);

CKINVDCx20_ASAP7_75t_R g2318 ( 
.A(n_2130),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2142),
.Y(n_2319)
);

CKINVDCx5p33_ASAP7_75t_R g2320 ( 
.A(n_2233),
.Y(n_2320)
);

CKINVDCx5p33_ASAP7_75t_R g2321 ( 
.A(n_2081),
.Y(n_2321)
);

BUFx6f_ASAP7_75t_L g2322 ( 
.A(n_2161),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2044),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_2175),
.B(n_1658),
.Y(n_2324)
);

INVx4_ASAP7_75t_L g2325 ( 
.A(n_2171),
.Y(n_2325)
);

CKINVDCx5p33_ASAP7_75t_R g2326 ( 
.A(n_2081),
.Y(n_2326)
);

HB1xp67_ASAP7_75t_L g2327 ( 
.A(n_2234),
.Y(n_2327)
);

CKINVDCx5p33_ASAP7_75t_R g2328 ( 
.A(n_2119),
.Y(n_2328)
);

CKINVDCx5p33_ASAP7_75t_R g2329 ( 
.A(n_2066),
.Y(n_2329)
);

CKINVDCx5p33_ASAP7_75t_R g2330 ( 
.A(n_2151),
.Y(n_2330)
);

CKINVDCx20_ASAP7_75t_R g2331 ( 
.A(n_2073),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2110),
.Y(n_2332)
);

CKINVDCx5p33_ASAP7_75t_R g2333 ( 
.A(n_2159),
.Y(n_2333)
);

CKINVDCx5p33_ASAP7_75t_R g2334 ( 
.A(n_2111),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_2090),
.Y(n_2335)
);

CKINVDCx5p33_ASAP7_75t_R g2336 ( 
.A(n_2147),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2141),
.Y(n_2337)
);

NOR2xp33_ASAP7_75t_R g2338 ( 
.A(n_2223),
.B(n_1351),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2044),
.Y(n_2339)
);

NOR2xp67_ASAP7_75t_L g2340 ( 
.A(n_2078),
.B(n_1),
.Y(n_2340)
);

NOR2xp33_ASAP7_75t_L g2341 ( 
.A(n_2041),
.B(n_1677),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2055),
.B(n_1532),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2144),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2160),
.Y(n_2344)
);

CKINVDCx5p33_ASAP7_75t_R g2345 ( 
.A(n_2169),
.Y(n_2345)
);

HB1xp67_ASAP7_75t_L g2346 ( 
.A(n_2192),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2176),
.Y(n_2347)
);

CKINVDCx20_ASAP7_75t_R g2348 ( 
.A(n_2097),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2182),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2187),
.Y(n_2350)
);

CKINVDCx5p33_ASAP7_75t_R g2351 ( 
.A(n_2226),
.Y(n_2351)
);

AOI22xp5_ASAP7_75t_L g2352 ( 
.A1(n_2091),
.A2(n_1689),
.B1(n_1706),
.B2(n_1683),
.Y(n_2352)
);

NOR2xp33_ASAP7_75t_R g2353 ( 
.A(n_2266),
.B(n_1373),
.Y(n_2353)
);

INVx3_ASAP7_75t_L g2354 ( 
.A(n_2038),
.Y(n_2354)
);

CKINVDCx5p33_ASAP7_75t_R g2355 ( 
.A(n_2070),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_R g2356 ( 
.A(n_2137),
.B(n_1373),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2162),
.Y(n_2357)
);

AND2x4_ASAP7_75t_L g2358 ( 
.A(n_2207),
.B(n_1802),
.Y(n_2358)
);

CKINVDCx5p33_ASAP7_75t_R g2359 ( 
.A(n_2179),
.Y(n_2359)
);

CKINVDCx5p33_ASAP7_75t_R g2360 ( 
.A(n_2072),
.Y(n_2360)
);

CKINVDCx20_ASAP7_75t_R g2361 ( 
.A(n_2149),
.Y(n_2361)
);

CKINVDCx5p33_ASAP7_75t_R g2362 ( 
.A(n_2190),
.Y(n_2362)
);

CKINVDCx5p33_ASAP7_75t_R g2363 ( 
.A(n_2190),
.Y(n_2363)
);

NOR2xp33_ASAP7_75t_R g2364 ( 
.A(n_2083),
.B(n_1385),
.Y(n_2364)
);

CKINVDCx5p33_ASAP7_75t_R g2365 ( 
.A(n_2198),
.Y(n_2365)
);

CKINVDCx5p33_ASAP7_75t_R g2366 ( 
.A(n_2222),
.Y(n_2366)
);

CKINVDCx20_ASAP7_75t_R g2367 ( 
.A(n_2197),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2065),
.B(n_1709),
.Y(n_2368)
);

CKINVDCx5p33_ASAP7_75t_R g2369 ( 
.A(n_2276),
.Y(n_2369)
);

HB1xp67_ASAP7_75t_L g2370 ( 
.A(n_2209),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2050),
.Y(n_2371)
);

NOR2xp33_ASAP7_75t_R g2372 ( 
.A(n_2136),
.B(n_1385),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2082),
.B(n_1715),
.Y(n_2373)
);

CKINVDCx5p33_ASAP7_75t_R g2374 ( 
.A(n_2232),
.Y(n_2374)
);

CKINVDCx5p33_ASAP7_75t_R g2375 ( 
.A(n_2238),
.Y(n_2375)
);

NOR2xp33_ASAP7_75t_R g2376 ( 
.A(n_2102),
.B(n_1396),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2051),
.Y(n_2377)
);

INVx3_ASAP7_75t_L g2378 ( 
.A(n_2038),
.Y(n_2378)
);

CKINVDCx5p33_ASAP7_75t_R g2379 ( 
.A(n_2249),
.Y(n_2379)
);

AOI21x1_ASAP7_75t_L g2380 ( 
.A1(n_2122),
.A2(n_1692),
.B(n_1187),
.Y(n_2380)
);

BUFx6f_ASAP7_75t_L g2381 ( 
.A(n_2171),
.Y(n_2381)
);

CKINVDCx5p33_ASAP7_75t_R g2382 ( 
.A(n_2256),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2084),
.Y(n_2383)
);

CKINVDCx20_ASAP7_75t_R g2384 ( 
.A(n_2268),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2087),
.Y(n_2385)
);

CKINVDCx5p33_ASAP7_75t_R g2386 ( 
.A(n_2282),
.Y(n_2386)
);

NAND2xp33_ASAP7_75t_L g2387 ( 
.A(n_2171),
.B(n_1581),
.Y(n_2387)
);

CKINVDCx5p33_ASAP7_75t_R g2388 ( 
.A(n_2228),
.Y(n_2388)
);

CKINVDCx5p33_ASAP7_75t_R g2389 ( 
.A(n_2278),
.Y(n_2389)
);

CKINVDCx5p33_ASAP7_75t_R g2390 ( 
.A(n_2148),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2049),
.Y(n_2391)
);

CKINVDCx5p33_ASAP7_75t_R g2392 ( 
.A(n_2208),
.Y(n_2392)
);

BUFx2_ASAP7_75t_L g2393 ( 
.A(n_2237),
.Y(n_2393)
);

BUFx3_ASAP7_75t_L g2394 ( 
.A(n_2194),
.Y(n_2394)
);

AND2x4_ASAP7_75t_L g2395 ( 
.A(n_2207),
.B(n_1817),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_R g2396 ( 
.A(n_2243),
.B(n_1396),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2092),
.Y(n_2397)
);

CKINVDCx14_ASAP7_75t_R g2398 ( 
.A(n_2247),
.Y(n_2398)
);

CKINVDCx5p33_ASAP7_75t_R g2399 ( 
.A(n_2251),
.Y(n_2399)
);

NOR2xp33_ASAP7_75t_R g2400 ( 
.A(n_2254),
.B(n_1441),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2093),
.Y(n_2401)
);

CKINVDCx20_ASAP7_75t_R g2402 ( 
.A(n_2258),
.Y(n_2402)
);

OAI21x1_ASAP7_75t_L g2403 ( 
.A1(n_2188),
.A2(n_1281),
.B(n_1220),
.Y(n_2403)
);

INVx2_ASAP7_75t_SL g2404 ( 
.A(n_2204),
.Y(n_2404)
);

CKINVDCx5p33_ASAP7_75t_R g2405 ( 
.A(n_2153),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_SL g2406 ( 
.A(n_2174),
.B(n_1736),
.Y(n_2406)
);

CKINVDCx20_ASAP7_75t_R g2407 ( 
.A(n_2191),
.Y(n_2407)
);

NAND2xp33_ASAP7_75t_R g2408 ( 
.A(n_2094),
.B(n_1745),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2129),
.Y(n_2409)
);

CKINVDCx5p33_ASAP7_75t_R g2410 ( 
.A(n_2040),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2138),
.Y(n_2411)
);

BUFx3_ASAP7_75t_L g2412 ( 
.A(n_2194),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2049),
.Y(n_2413)
);

CKINVDCx5p33_ASAP7_75t_R g2414 ( 
.A(n_2040),
.Y(n_2414)
);

AOI21x1_ASAP7_75t_L g2415 ( 
.A1(n_2045),
.A2(n_1192),
.B(n_1186),
.Y(n_2415)
);

CKINVDCx5p33_ASAP7_75t_R g2416 ( 
.A(n_2059),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2060),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2060),
.Y(n_2418)
);

CKINVDCx20_ASAP7_75t_R g2419 ( 
.A(n_2108),
.Y(n_2419)
);

CKINVDCx20_ASAP7_75t_R g2420 ( 
.A(n_2043),
.Y(n_2420)
);

CKINVDCx20_ASAP7_75t_R g2421 ( 
.A(n_2196),
.Y(n_2421)
);

CKINVDCx5p33_ASAP7_75t_R g2422 ( 
.A(n_2121),
.Y(n_2422)
);

CKINVDCx20_ASAP7_75t_R g2423 ( 
.A(n_2200),
.Y(n_2423)
);

CKINVDCx5p33_ASAP7_75t_R g2424 ( 
.A(n_2127),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2064),
.Y(n_2425)
);

CKINVDCx5p33_ASAP7_75t_R g2426 ( 
.A(n_2143),
.Y(n_2426)
);

NOR2xp33_ASAP7_75t_L g2427 ( 
.A(n_2214),
.B(n_1746),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2064),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2076),
.Y(n_2429)
);

AOI21x1_ASAP7_75t_L g2430 ( 
.A1(n_2054),
.A2(n_2113),
.B(n_2106),
.Y(n_2430)
);

NOR2xp67_ASAP7_75t_L g2431 ( 
.A(n_2236),
.B(n_1),
.Y(n_2431)
);

NOR2x1p5_ASAP7_75t_L g2432 ( 
.A(n_2219),
.B(n_1754),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2076),
.Y(n_2433)
);

BUFx3_ASAP7_75t_L g2434 ( 
.A(n_2195),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2085),
.Y(n_2435)
);

CKINVDCx5p33_ASAP7_75t_R g2436 ( 
.A(n_2145),
.Y(n_2436)
);

CKINVDCx5p33_ASAP7_75t_R g2437 ( 
.A(n_2213),
.Y(n_2437)
);

CKINVDCx5p33_ASAP7_75t_R g2438 ( 
.A(n_2235),
.Y(n_2438)
);

CKINVDCx5p33_ASAP7_75t_R g2439 ( 
.A(n_2272),
.Y(n_2439)
);

HB1xp67_ASAP7_75t_L g2440 ( 
.A(n_2215),
.Y(n_2440)
);

CKINVDCx5p33_ASAP7_75t_R g2441 ( 
.A(n_2279),
.Y(n_2441)
);

CKINVDCx20_ASAP7_75t_R g2442 ( 
.A(n_2047),
.Y(n_2442)
);

BUFx2_ASAP7_75t_L g2443 ( 
.A(n_2189),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2085),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2128),
.B(n_1762),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_2099),
.Y(n_2446)
);

INVx2_ASAP7_75t_SL g2447 ( 
.A(n_2261),
.Y(n_2447)
);

CKINVDCx5p33_ASAP7_75t_R g2448 ( 
.A(n_2062),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2099),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2100),
.Y(n_2450)
);

NOR2xp33_ASAP7_75t_R g2451 ( 
.A(n_2259),
.B(n_1441),
.Y(n_2451)
);

BUFx10_ASAP7_75t_L g2452 ( 
.A(n_2269),
.Y(n_2452)
);

INVx5_ASAP7_75t_L g2453 ( 
.A(n_2195),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2100),
.Y(n_2454)
);

BUFx6f_ASAP7_75t_L g2455 ( 
.A(n_2202),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_SL g2456 ( 
.A(n_2156),
.B(n_1766),
.Y(n_2456)
);

CKINVDCx5p33_ASAP7_75t_R g2457 ( 
.A(n_2281),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2104),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2104),
.Y(n_2459)
);

CKINVDCx20_ASAP7_75t_R g2460 ( 
.A(n_2139),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2077),
.B(n_1532),
.Y(n_2461)
);

CKINVDCx5p33_ASAP7_75t_R g2462 ( 
.A(n_2042),
.Y(n_2462)
);

CKINVDCx5p33_ASAP7_75t_R g2463 ( 
.A(n_2071),
.Y(n_2463)
);

CKINVDCx5p33_ASAP7_75t_R g2464 ( 
.A(n_2236),
.Y(n_2464)
);

CKINVDCx5p33_ASAP7_75t_R g2465 ( 
.A(n_2095),
.Y(n_2465)
);

CKINVDCx5p33_ASAP7_75t_R g2466 ( 
.A(n_2283),
.Y(n_2466)
);

CKINVDCx20_ASAP7_75t_R g2467 ( 
.A(n_2260),
.Y(n_2467)
);

CKINVDCx5p33_ASAP7_75t_R g2468 ( 
.A(n_2262),
.Y(n_2468)
);

CKINVDCx5p33_ASAP7_75t_R g2469 ( 
.A(n_2202),
.Y(n_2469)
);

CKINVDCx5p33_ASAP7_75t_R g2470 ( 
.A(n_2206),
.Y(n_2470)
);

NOR2xp33_ASAP7_75t_R g2471 ( 
.A(n_2259),
.B(n_1451),
.Y(n_2471)
);

CKINVDCx5p33_ASAP7_75t_R g2472 ( 
.A(n_2206),
.Y(n_2472)
);

CKINVDCx5p33_ASAP7_75t_R g2473 ( 
.A(n_2212),
.Y(n_2473)
);

CKINVDCx5p33_ASAP7_75t_R g2474 ( 
.A(n_2212),
.Y(n_2474)
);

CKINVDCx5p33_ASAP7_75t_R g2475 ( 
.A(n_2217),
.Y(n_2475)
);

AND3x2_ASAP7_75t_L g2476 ( 
.A(n_2183),
.B(n_1459),
.C(n_1451),
.Y(n_2476)
);

INVx2_ASAP7_75t_L g2477 ( 
.A(n_2107),
.Y(n_2477)
);

NOR2xp33_ASAP7_75t_R g2478 ( 
.A(n_2259),
.B(n_1459),
.Y(n_2478)
);

CKINVDCx20_ASAP7_75t_R g2479 ( 
.A(n_2217),
.Y(n_2479)
);

BUFx2_ASAP7_75t_L g2480 ( 
.A(n_2185),
.Y(n_2480)
);

HB1xp67_ASAP7_75t_L g2481 ( 
.A(n_2165),
.Y(n_2481)
);

CKINVDCx20_ASAP7_75t_R g2482 ( 
.A(n_2227),
.Y(n_2482)
);

NAND2xp33_ASAP7_75t_R g2483 ( 
.A(n_2063),
.B(n_1807),
.Y(n_2483)
);

CKINVDCx5p33_ASAP7_75t_R g2484 ( 
.A(n_2227),
.Y(n_2484)
);

CKINVDCx5p33_ASAP7_75t_R g2485 ( 
.A(n_2239),
.Y(n_2485)
);

CKINVDCx5p33_ASAP7_75t_R g2486 ( 
.A(n_2239),
.Y(n_2486)
);

CKINVDCx5p33_ASAP7_75t_R g2487 ( 
.A(n_2242),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2107),
.Y(n_2488)
);

NOR2xp67_ASAP7_75t_L g2489 ( 
.A(n_2199),
.B(n_1),
.Y(n_2489)
);

CKINVDCx5p33_ASAP7_75t_R g2490 ( 
.A(n_2242),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2109),
.Y(n_2491)
);

INVx2_ASAP7_75t_SL g2492 ( 
.A(n_2069),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2109),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2115),
.Y(n_2494)
);

CKINVDCx5p33_ASAP7_75t_R g2495 ( 
.A(n_2250),
.Y(n_2495)
);

CKINVDCx5p33_ASAP7_75t_R g2496 ( 
.A(n_2250),
.Y(n_2496)
);

CKINVDCx5p33_ASAP7_75t_R g2497 ( 
.A(n_2257),
.Y(n_2497)
);

CKINVDCx20_ASAP7_75t_R g2498 ( 
.A(n_2257),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2115),
.Y(n_2499)
);

CKINVDCx20_ASAP7_75t_R g2500 ( 
.A(n_2263),
.Y(n_2500)
);

CKINVDCx5p33_ASAP7_75t_R g2501 ( 
.A(n_2263),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2123),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_2265),
.Y(n_2503)
);

CKINVDCx5p33_ASAP7_75t_R g2504 ( 
.A(n_2265),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2123),
.Y(n_2505)
);

CKINVDCx5p33_ASAP7_75t_R g2506 ( 
.A(n_2098),
.Y(n_2506)
);

CKINVDCx5p33_ASAP7_75t_R g2507 ( 
.A(n_2103),
.Y(n_2507)
);

CKINVDCx16_ASAP7_75t_R g2508 ( 
.A(n_2075),
.Y(n_2508)
);

AOI22xp5_ASAP7_75t_L g2509 ( 
.A1(n_2105),
.A2(n_1818),
.B1(n_1823),
.B2(n_1814),
.Y(n_2509)
);

CKINVDCx5p33_ASAP7_75t_R g2510 ( 
.A(n_2118),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2134),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2134),
.Y(n_2512)
);

CKINVDCx5p33_ASAP7_75t_R g2513 ( 
.A(n_2120),
.Y(n_2513)
);

INVxp67_ASAP7_75t_L g2514 ( 
.A(n_2150),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2150),
.Y(n_2515)
);

BUFx2_ASAP7_75t_L g2516 ( 
.A(n_2053),
.Y(n_2516)
);

CKINVDCx5p33_ASAP7_75t_R g2517 ( 
.A(n_2146),
.Y(n_2517)
);

NOR2xp33_ASAP7_75t_R g2518 ( 
.A(n_2057),
.B(n_1473),
.Y(n_2518)
);

CKINVDCx5p33_ASAP7_75t_R g2519 ( 
.A(n_2155),
.Y(n_2519)
);

INVx3_ASAP7_75t_L g2520 ( 
.A(n_2152),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2152),
.Y(n_2521)
);

CKINVDCx5p33_ASAP7_75t_R g2522 ( 
.A(n_2157),
.Y(n_2522)
);

CKINVDCx5p33_ASAP7_75t_R g2523 ( 
.A(n_2058),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2068),
.B(n_1836),
.Y(n_2524)
);

BUFx6f_ASAP7_75t_SL g2525 ( 
.A(n_2074),
.Y(n_2525)
);

CKINVDCx5p33_ASAP7_75t_R g2526 ( 
.A(n_2080),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2163),
.Y(n_2527)
);

CKINVDCx5p33_ASAP7_75t_R g2528 ( 
.A(n_2086),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2163),
.Y(n_2529)
);

CKINVDCx5p33_ASAP7_75t_R g2530 ( 
.A(n_2096),
.Y(n_2530)
);

NOR2xp33_ASAP7_75t_R g2531 ( 
.A(n_2203),
.B(n_1473),
.Y(n_2531)
);

CKINVDCx5p33_ASAP7_75t_R g2532 ( 
.A(n_2201),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2210),
.Y(n_2533)
);

CKINVDCx20_ASAP7_75t_R g2534 ( 
.A(n_2205),
.Y(n_2534)
);

CKINVDCx5p33_ASAP7_75t_R g2535 ( 
.A(n_2224),
.Y(n_2535)
);

CKINVDCx5p33_ASAP7_75t_R g2536 ( 
.A(n_2225),
.Y(n_2536)
);

CKINVDCx20_ASAP7_75t_R g2537 ( 
.A(n_2211),
.Y(n_2537)
);

CKINVDCx5p33_ASAP7_75t_R g2538 ( 
.A(n_2230),
.Y(n_2538)
);

HB1xp67_ASAP7_75t_L g2539 ( 
.A(n_2039),
.Y(n_2539)
);

INVxp67_ASAP7_75t_L g2540 ( 
.A(n_2181),
.Y(n_2540)
);

CKINVDCx5p33_ASAP7_75t_R g2541 ( 
.A(n_2241),
.Y(n_2541)
);

CKINVDCx5p33_ASAP7_75t_R g2542 ( 
.A(n_2246),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2154),
.Y(n_2543)
);

BUFx2_ASAP7_75t_L g2544 ( 
.A(n_2216),
.Y(n_2544)
);

INVx3_ASAP7_75t_L g2545 ( 
.A(n_2248),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2158),
.Y(n_2546)
);

CKINVDCx5p33_ASAP7_75t_R g2547 ( 
.A(n_2253),
.Y(n_2547)
);

INVx3_ASAP7_75t_L g2548 ( 
.A(n_2267),
.Y(n_2548)
);

HB1xp67_ASAP7_75t_L g2549 ( 
.A(n_2218),
.Y(n_2549)
);

CKINVDCx5p33_ASAP7_75t_R g2550 ( 
.A(n_2271),
.Y(n_2550)
);

CKINVDCx5p33_ASAP7_75t_R g2551 ( 
.A(n_2284),
.Y(n_2551)
);

BUFx6f_ASAP7_75t_L g2552 ( 
.A(n_2166),
.Y(n_2552)
);

CKINVDCx5p33_ASAP7_75t_R g2553 ( 
.A(n_2220),
.Y(n_2553)
);

CKINVDCx5p33_ASAP7_75t_R g2554 ( 
.A(n_2229),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2164),
.Y(n_2555)
);

CKINVDCx5p33_ASAP7_75t_R g2556 ( 
.A(n_2231),
.Y(n_2556)
);

NOR2xp67_ASAP7_75t_L g2557 ( 
.A(n_2280),
.B(n_1),
.Y(n_2557)
);

CKINVDCx5p33_ASAP7_75t_R g2558 ( 
.A(n_2244),
.Y(n_2558)
);

CKINVDCx5p33_ASAP7_75t_R g2559 ( 
.A(n_2245),
.Y(n_2559)
);

CKINVDCx5p33_ASAP7_75t_R g2560 ( 
.A(n_2264),
.Y(n_2560)
);

CKINVDCx5p33_ASAP7_75t_R g2561 ( 
.A(n_2270),
.Y(n_2561)
);

INVxp67_ASAP7_75t_SL g2562 ( 
.A(n_2186),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2167),
.Y(n_2563)
);

CKINVDCx5p33_ASAP7_75t_R g2564 ( 
.A(n_2274),
.Y(n_2564)
);

CKINVDCx5p33_ASAP7_75t_R g2565 ( 
.A(n_2275),
.Y(n_2565)
);

BUFx6f_ASAP7_75t_L g2566 ( 
.A(n_2168),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2178),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2277),
.B(n_1855),
.Y(n_2568)
);

NOR2xp33_ASAP7_75t_R g2569 ( 
.A(n_2114),
.B(n_1547),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2088),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2125),
.Y(n_2571)
);

CKINVDCx5p33_ASAP7_75t_R g2572 ( 
.A(n_2079),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2061),
.Y(n_2573)
);

CKINVDCx5p33_ASAP7_75t_R g2574 ( 
.A(n_2079),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2131),
.Y(n_2575)
);

CKINVDCx5p33_ASAP7_75t_R g2576 ( 
.A(n_2079),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2131),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2131),
.Y(n_2578)
);

CKINVDCx5p33_ASAP7_75t_R g2579 ( 
.A(n_2079),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2131),
.Y(n_2580)
);

NOR2xp33_ASAP7_75t_L g2581 ( 
.A(n_2041),
.B(n_1864),
.Y(n_2581)
);

CKINVDCx5p33_ASAP7_75t_R g2582 ( 
.A(n_2079),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2131),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2131),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2131),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2061),
.Y(n_2586)
);

CKINVDCx5p33_ASAP7_75t_R g2587 ( 
.A(n_2079),
.Y(n_2587)
);

NOR2xp67_ASAP7_75t_L g2588 ( 
.A(n_2234),
.B(n_2),
.Y(n_2588)
);

CKINVDCx20_ASAP7_75t_R g2589 ( 
.A(n_2079),
.Y(n_2589)
);

OAI22xp5_ASAP7_75t_SL g2590 ( 
.A1(n_2124),
.A2(n_1561),
.B1(n_1633),
.B2(n_1547),
.Y(n_2590)
);

CKINVDCx20_ASAP7_75t_R g2591 ( 
.A(n_2079),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_SL g2592 ( 
.A(n_2161),
.B(n_1866),
.Y(n_2592)
);

BUFx10_ASAP7_75t_L g2593 ( 
.A(n_2066),
.Y(n_2593)
);

CKINVDCx20_ASAP7_75t_R g2594 ( 
.A(n_2079),
.Y(n_2594)
);

CKINVDCx5p33_ASAP7_75t_R g2595 ( 
.A(n_2079),
.Y(n_2595)
);

CKINVDCx5p33_ASAP7_75t_R g2596 ( 
.A(n_2079),
.Y(n_2596)
);

CKINVDCx5p33_ASAP7_75t_R g2597 ( 
.A(n_2079),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_SL g2598 ( 
.A(n_2161),
.B(n_1873),
.Y(n_2598)
);

CKINVDCx5p33_ASAP7_75t_R g2599 ( 
.A(n_2079),
.Y(n_2599)
);

CKINVDCx20_ASAP7_75t_R g2600 ( 
.A(n_2079),
.Y(n_2600)
);

CKINVDCx5p33_ASAP7_75t_R g2601 ( 
.A(n_2079),
.Y(n_2601)
);

NOR2xp33_ASAP7_75t_R g2602 ( 
.A(n_2117),
.B(n_1561),
.Y(n_2602)
);

HB1xp67_ASAP7_75t_L g2603 ( 
.A(n_2056),
.Y(n_2603)
);

CKINVDCx20_ASAP7_75t_R g2604 ( 
.A(n_2079),
.Y(n_2604)
);

INVx3_ASAP7_75t_L g2605 ( 
.A(n_2110),
.Y(n_2605)
);

CKINVDCx5p33_ASAP7_75t_R g2606 ( 
.A(n_2079),
.Y(n_2606)
);

HB1xp67_ASAP7_75t_L g2607 ( 
.A(n_2056),
.Y(n_2607)
);

CKINVDCx5p33_ASAP7_75t_R g2608 ( 
.A(n_2079),
.Y(n_2608)
);

CKINVDCx5p33_ASAP7_75t_R g2609 ( 
.A(n_2079),
.Y(n_2609)
);

CKINVDCx5p33_ASAP7_75t_R g2610 ( 
.A(n_2079),
.Y(n_2610)
);

CKINVDCx5p33_ASAP7_75t_R g2611 ( 
.A(n_2079),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2131),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2131),
.Y(n_2613)
);

NAND2xp33_ASAP7_75t_R g2614 ( 
.A(n_2116),
.B(n_1166),
.Y(n_2614)
);

CKINVDCx5p33_ASAP7_75t_R g2615 ( 
.A(n_2079),
.Y(n_2615)
);

CKINVDCx5p33_ASAP7_75t_R g2616 ( 
.A(n_2079),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2131),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2357),
.Y(n_2618)
);

INVxp67_ASAP7_75t_L g2619 ( 
.A(n_2292),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_2562),
.B(n_1335),
.Y(n_2620)
);

INVx4_ASAP7_75t_L g2621 ( 
.A(n_2302),
.Y(n_2621)
);

INVxp67_ASAP7_75t_SL g2622 ( 
.A(n_2603),
.Y(n_2622)
);

OR2x2_ASAP7_75t_L g2623 ( 
.A(n_2305),
.B(n_1211),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2552),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_2540),
.B(n_1718),
.Y(n_2625)
);

INVx2_ASAP7_75t_SL g2626 ( 
.A(n_2593),
.Y(n_2626)
);

BUFx2_ASAP7_75t_L g2627 ( 
.A(n_2384),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_2327),
.B(n_1633),
.Y(n_2628)
);

OR2x6_ASAP7_75t_L g2629 ( 
.A(n_2590),
.B(n_1817),
.Y(n_2629)
);

AND2x2_ASAP7_75t_L g2630 ( 
.A(n_2316),
.B(n_1653),
.Y(n_2630)
);

INVx3_ASAP7_75t_L g2631 ( 
.A(n_2593),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2552),
.Y(n_2632)
);

AND2x4_ASAP7_75t_L g2633 ( 
.A(n_2331),
.B(n_1653),
.Y(n_2633)
);

BUFx6f_ASAP7_75t_L g2634 ( 
.A(n_2322),
.Y(n_2634)
);

INVx3_ASAP7_75t_L g2635 ( 
.A(n_2322),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2427),
.B(n_1167),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2352),
.B(n_2297),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2409),
.Y(n_2638)
);

BUFx2_ASAP7_75t_L g2639 ( 
.A(n_2364),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2411),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2297),
.B(n_1168),
.Y(n_2641)
);

NOR2xp33_ASAP7_75t_L g2642 ( 
.A(n_2437),
.B(n_1665),
.Y(n_2642)
);

BUFx6f_ASAP7_75t_L g2643 ( 
.A(n_2322),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2371),
.Y(n_2644)
);

INVx3_ASAP7_75t_L g2645 ( 
.A(n_2306),
.Y(n_2645)
);

CKINVDCx5p33_ASAP7_75t_R g2646 ( 
.A(n_2338),
.Y(n_2646)
);

INVx3_ASAP7_75t_L g2647 ( 
.A(n_2306),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_L g2648 ( 
.A(n_2448),
.B(n_1169),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2377),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2368),
.B(n_1170),
.Y(n_2650)
);

BUFx6f_ASAP7_75t_L g2651 ( 
.A(n_2381),
.Y(n_2651)
);

BUFx6f_ASAP7_75t_L g2652 ( 
.A(n_2381),
.Y(n_2652)
);

CKINVDCx20_ASAP7_75t_R g2653 ( 
.A(n_2295),
.Y(n_2653)
);

AND2x4_ASAP7_75t_L g2654 ( 
.A(n_2607),
.B(n_1665),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2373),
.B(n_1176),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2552),
.Y(n_2656)
);

BUFx6f_ASAP7_75t_L g2657 ( 
.A(n_2381),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2445),
.B(n_1177),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2286),
.Y(n_2659)
);

INVx5_ASAP7_75t_L g2660 ( 
.A(n_2291),
.Y(n_2660)
);

CKINVDCx5p33_ASAP7_75t_R g2661 ( 
.A(n_2353),
.Y(n_2661)
);

NOR2xp33_ASAP7_75t_L g2662 ( 
.A(n_2438),
.B(n_1668),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2288),
.Y(n_2663)
);

BUFx3_ASAP7_75t_L g2664 ( 
.A(n_2479),
.Y(n_2664)
);

HB1xp67_ASAP7_75t_L g2665 ( 
.A(n_2569),
.Y(n_2665)
);

AND2x2_ASAP7_75t_L g2666 ( 
.A(n_2346),
.B(n_1668),
.Y(n_2666)
);

INVx3_ASAP7_75t_L g2667 ( 
.A(n_2394),
.Y(n_2667)
);

NOR2xp33_ASAP7_75t_L g2668 ( 
.A(n_2439),
.B(n_1704),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2289),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2341),
.B(n_1179),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2301),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2566),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_SL g2673 ( 
.A(n_2325),
.B(n_1330),
.Y(n_2673)
);

BUFx2_ASAP7_75t_L g2674 ( 
.A(n_2300),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2304),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2319),
.Y(n_2676)
);

NAND2x1p5_ASAP7_75t_L g2677 ( 
.A(n_2443),
.B(n_1215),
.Y(n_2677)
);

NOR2xp33_ASAP7_75t_L g2678 ( 
.A(n_2441),
.B(n_1704),
.Y(n_2678)
);

NOR2xp33_ASAP7_75t_L g2679 ( 
.A(n_2398),
.B(n_1729),
.Y(n_2679)
);

NOR2xp33_ASAP7_75t_L g2680 ( 
.A(n_2393),
.B(n_1729),
.Y(n_2680)
);

INVx2_ASAP7_75t_SL g2681 ( 
.A(n_2358),
.Y(n_2681)
);

NOR2xp33_ASAP7_75t_L g2682 ( 
.A(n_2462),
.B(n_2463),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_SL g2683 ( 
.A(n_2325),
.B(n_1443),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2581),
.B(n_1180),
.Y(n_2684)
);

INVx4_ASAP7_75t_L g2685 ( 
.A(n_2334),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2575),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2577),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2578),
.Y(n_2688)
);

HB1xp67_ASAP7_75t_L g2689 ( 
.A(n_2370),
.Y(n_2689)
);

NAND2x1p5_ASAP7_75t_L g2690 ( 
.A(n_2605),
.B(n_1286),
.Y(n_2690)
);

AND2x6_ASAP7_75t_L g2691 ( 
.A(n_2299),
.B(n_1406),
.Y(n_2691)
);

INVx2_ASAP7_75t_L g2692 ( 
.A(n_2566),
.Y(n_2692)
);

INVx5_ASAP7_75t_L g2693 ( 
.A(n_2455),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2580),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2342),
.B(n_1743),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2509),
.B(n_1181),
.Y(n_2696)
);

INVx4_ASAP7_75t_L g2697 ( 
.A(n_2422),
.Y(n_2697)
);

AND2x4_ASAP7_75t_L g2698 ( 
.A(n_2351),
.B(n_1743),
.Y(n_2698)
);

BUFx3_ASAP7_75t_L g2699 ( 
.A(n_2482),
.Y(n_2699)
);

OR2x2_ASAP7_75t_L g2700 ( 
.A(n_2320),
.B(n_1293),
.Y(n_2700)
);

AND2x2_ASAP7_75t_L g2701 ( 
.A(n_2518),
.B(n_1813),
.Y(n_2701)
);

AND2x4_ASAP7_75t_L g2702 ( 
.A(n_2355),
.B(n_1813),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2583),
.Y(n_2703)
);

INVxp67_ASAP7_75t_L g2704 ( 
.A(n_2614),
.Y(n_2704)
);

NOR2xp33_ASAP7_75t_L g2705 ( 
.A(n_2424),
.B(n_1816),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2566),
.Y(n_2706)
);

AND2x6_ASAP7_75t_L g2707 ( 
.A(n_2294),
.B(n_1406),
.Y(n_2707)
);

AOI22xp5_ASAP7_75t_L g2708 ( 
.A1(n_2442),
.A2(n_1822),
.B1(n_1832),
.B2(n_1816),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2584),
.Y(n_2709)
);

INVx2_ASAP7_75t_L g2710 ( 
.A(n_2308),
.Y(n_2710)
);

AND3x2_ASAP7_75t_L g2711 ( 
.A(n_2348),
.B(n_1832),
.C(n_1822),
.Y(n_2711)
);

CKINVDCx5p33_ASAP7_75t_R g2712 ( 
.A(n_2356),
.Y(n_2712)
);

AND2x2_ASAP7_75t_L g2713 ( 
.A(n_2382),
.B(n_1840),
.Y(n_2713)
);

BUFx10_ASAP7_75t_L g2714 ( 
.A(n_2314),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2312),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2313),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2585),
.Y(n_2717)
);

AND2x6_ASAP7_75t_L g2718 ( 
.A(n_2317),
.B(n_1406),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2524),
.B(n_1190),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2612),
.Y(n_2720)
);

AND2x6_ASAP7_75t_L g2721 ( 
.A(n_2573),
.B(n_1406),
.Y(n_2721)
);

AND2x4_ASAP7_75t_L g2722 ( 
.A(n_2318),
.B(n_1840),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2613),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2617),
.Y(n_2724)
);

AOI22xp33_ASAP7_75t_L g2725 ( 
.A1(n_2516),
.A2(n_1879),
.B1(n_1567),
.B2(n_1657),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2543),
.Y(n_2726)
);

CKINVDCx16_ASAP7_75t_R g2727 ( 
.A(n_2303),
.Y(n_2727)
);

INVx2_ASAP7_75t_SL g2728 ( 
.A(n_2358),
.Y(n_2728)
);

NAND2x1p5_ASAP7_75t_L g2729 ( 
.A(n_2605),
.B(n_1308),
.Y(n_2729)
);

INVx1_ASAP7_75t_SL g2730 ( 
.A(n_2602),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_SL g2731 ( 
.A(n_2340),
.B(n_1497),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2586),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_SL g2733 ( 
.A(n_2588),
.B(n_2388),
.Y(n_2733)
);

AND2x4_ASAP7_75t_L g2734 ( 
.A(n_2461),
.B(n_1879),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2546),
.Y(n_2735)
);

INVx5_ASAP7_75t_L g2736 ( 
.A(n_2455),
.Y(n_2736)
);

AND2x2_ASAP7_75t_L g2737 ( 
.A(n_2386),
.B(n_1532),
.Y(n_2737)
);

INVx4_ASAP7_75t_L g2738 ( 
.A(n_2389),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2555),
.Y(n_2739)
);

INVx2_ASAP7_75t_SL g2740 ( 
.A(n_2395),
.Y(n_2740)
);

OR2x6_ASAP7_75t_L g2741 ( 
.A(n_2404),
.B(n_1220),
.Y(n_2741)
);

NOR2xp33_ASAP7_75t_L g2742 ( 
.A(n_2426),
.B(n_1191),
.Y(n_2742)
);

INVx3_ASAP7_75t_L g2743 ( 
.A(n_2412),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2430),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_SL g2745 ( 
.A(n_2506),
.B(n_1194),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2563),
.B(n_1202),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2335),
.B(n_1567),
.Y(n_2747)
);

INVxp67_ASAP7_75t_SL g2748 ( 
.A(n_2467),
.Y(n_2748)
);

AOI22xp33_ASAP7_75t_L g2749 ( 
.A1(n_2507),
.A2(n_1657),
.B1(n_1659),
.B2(n_1567),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2567),
.Y(n_2750)
);

BUFx2_ASAP7_75t_L g2751 ( 
.A(n_2531),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2415),
.Y(n_2752)
);

BUFx6f_ASAP7_75t_L g2753 ( 
.A(n_2455),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2380),
.Y(n_2754)
);

AND2x6_ASAP7_75t_L g2755 ( 
.A(n_2344),
.B(n_1527),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2539),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2403),
.Y(n_2757)
);

AND2x4_ASAP7_75t_L g2758 ( 
.A(n_2309),
.B(n_1317),
.Y(n_2758)
);

BUFx3_ASAP7_75t_L g2759 ( 
.A(n_2498),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2510),
.B(n_1204),
.Y(n_2760)
);

BUFx6f_ASAP7_75t_L g2761 ( 
.A(n_2434),
.Y(n_2761)
);

OR2x2_ASAP7_75t_L g2762 ( 
.A(n_2360),
.B(n_1366),
.Y(n_2762)
);

BUFx6f_ASAP7_75t_L g2763 ( 
.A(n_2453),
.Y(n_2763)
);

INVx2_ASAP7_75t_SL g2764 ( 
.A(n_2395),
.Y(n_2764)
);

INVx3_ASAP7_75t_L g2765 ( 
.A(n_2315),
.Y(n_2765)
);

OAI22xp33_ASAP7_75t_SL g2766 ( 
.A1(n_2416),
.A2(n_1207),
.B1(n_1208),
.B2(n_1205),
.Y(n_2766)
);

AND2x6_ASAP7_75t_L g2767 ( 
.A(n_2347),
.B(n_1527),
.Y(n_2767)
);

INVx2_ASAP7_75t_L g2768 ( 
.A(n_2533),
.Y(n_2768)
);

AND2x6_ASAP7_75t_L g2769 ( 
.A(n_2349),
.B(n_1527),
.Y(n_2769)
);

INVx2_ASAP7_75t_SL g2770 ( 
.A(n_2451),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2513),
.B(n_1209),
.Y(n_2771)
);

BUFx6f_ASAP7_75t_L g2772 ( 
.A(n_2453),
.Y(n_2772)
);

INVx3_ASAP7_75t_L g2773 ( 
.A(n_2354),
.Y(n_2773)
);

AND2x6_ASAP7_75t_L g2774 ( 
.A(n_2350),
.B(n_1527),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2571),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2568),
.B(n_1214),
.Y(n_2776)
);

HB1xp67_ASAP7_75t_L g2777 ( 
.A(n_2376),
.Y(n_2777)
);

AND2x2_ASAP7_75t_L g2778 ( 
.A(n_2396),
.B(n_1657),
.Y(n_2778)
);

INVx4_ASAP7_75t_L g2779 ( 
.A(n_2296),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2549),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2332),
.Y(n_2781)
);

NOR2xp33_ASAP7_75t_L g2782 ( 
.A(n_2392),
.B(n_1217),
.Y(n_2782)
);

NOR2xp33_ASAP7_75t_L g2783 ( 
.A(n_2399),
.B(n_1219),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2337),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_SL g2785 ( 
.A(n_2471),
.B(n_2478),
.Y(n_2785)
);

HB1xp67_ASAP7_75t_L g2786 ( 
.A(n_2410),
.Y(n_2786)
);

OR2x6_ASAP7_75t_L g2787 ( 
.A(n_2447),
.B(n_1281),
.Y(n_2787)
);

INVx3_ASAP7_75t_L g2788 ( 
.A(n_2354),
.Y(n_2788)
);

INVxp67_ASAP7_75t_L g2789 ( 
.A(n_2483),
.Y(n_2789)
);

AND2x4_ASAP7_75t_L g2790 ( 
.A(n_2432),
.B(n_1392),
.Y(n_2790)
);

AND2x4_ASAP7_75t_L g2791 ( 
.A(n_2298),
.B(n_1398),
.Y(n_2791)
);

NOR2xp33_ASAP7_75t_L g2792 ( 
.A(n_2466),
.B(n_1221),
.Y(n_2792)
);

INVx4_ASAP7_75t_L g2793 ( 
.A(n_2329),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2343),
.Y(n_2794)
);

CKINVDCx8_ASAP7_75t_R g2795 ( 
.A(n_2345),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2383),
.Y(n_2796)
);

NOR2xp33_ASAP7_75t_L g2797 ( 
.A(n_2460),
.B(n_1224),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2385),
.Y(n_2798)
);

INVx4_ASAP7_75t_SL g2799 ( 
.A(n_2525),
.Y(n_2799)
);

AND2x4_ASAP7_75t_L g2800 ( 
.A(n_2492),
.B(n_1402),
.Y(n_2800)
);

INVx3_ASAP7_75t_L g2801 ( 
.A(n_2378),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2397),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2406),
.B(n_2456),
.Y(n_2803)
);

AND2x6_ASAP7_75t_L g2804 ( 
.A(n_2570),
.B(n_1596),
.Y(n_2804)
);

BUFx2_ASAP7_75t_L g2805 ( 
.A(n_2400),
.Y(n_2805)
);

BUFx6f_ASAP7_75t_L g2806 ( 
.A(n_2453),
.Y(n_2806)
);

AND2x2_ASAP7_75t_SL g2807 ( 
.A(n_2508),
.B(n_1313),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2517),
.B(n_1229),
.Y(n_2808)
);

OR2x2_ASAP7_75t_L g2809 ( 
.A(n_2365),
.B(n_1422),
.Y(n_2809)
);

INVx3_ASAP7_75t_L g2810 ( 
.A(n_2378),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2545),
.Y(n_2811)
);

INVx2_ASAP7_75t_L g2812 ( 
.A(n_2545),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_SL g2813 ( 
.A(n_2519),
.B(n_1231),
.Y(n_2813)
);

AND2x4_ASAP7_75t_L g2814 ( 
.A(n_2310),
.B(n_1444),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2548),
.Y(n_2815)
);

AND2x4_ASAP7_75t_L g2816 ( 
.A(n_2311),
.B(n_1543),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2401),
.Y(n_2817)
);

NOR2xp33_ASAP7_75t_L g2818 ( 
.A(n_2522),
.B(n_1237),
.Y(n_2818)
);

AND2x6_ASAP7_75t_L g2819 ( 
.A(n_2548),
.B(n_1596),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2489),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2520),
.Y(n_2821)
);

INVx4_ASAP7_75t_L g2822 ( 
.A(n_2469),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2544),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2523),
.B(n_1238),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2520),
.Y(n_2825)
);

BUFx3_ASAP7_75t_L g2826 ( 
.A(n_2500),
.Y(n_2826)
);

AND2x6_ASAP7_75t_L g2827 ( 
.A(n_2425),
.B(n_1596),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2481),
.Y(n_2828)
);

BUFx3_ASAP7_75t_L g2829 ( 
.A(n_2293),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2557),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2431),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2323),
.Y(n_2832)
);

NAND3xp33_ASAP7_75t_L g2833 ( 
.A(n_2390),
.B(n_1242),
.C(n_1240),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_SL g2834 ( 
.A(n_2526),
.B(n_1243),
.Y(n_2834)
);

BUFx3_ASAP7_75t_L g2835 ( 
.A(n_2285),
.Y(n_2835)
);

BUFx3_ASAP7_75t_L g2836 ( 
.A(n_2589),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2339),
.Y(n_2837)
);

NAND2xp33_ASAP7_75t_L g2838 ( 
.A(n_2464),
.B(n_2528),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2324),
.Y(n_2839)
);

CKINVDCx5p33_ASAP7_75t_R g2840 ( 
.A(n_2287),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2530),
.B(n_1244),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2592),
.Y(n_2842)
);

INVx5_ASAP7_75t_L g2843 ( 
.A(n_2480),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2366),
.B(n_1659),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_SL g2845 ( 
.A(n_2452),
.B(n_1247),
.Y(n_2845)
);

OR2x2_ASAP7_75t_L g2846 ( 
.A(n_2336),
.B(n_1551),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2598),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2391),
.Y(n_2848)
);

OR2x2_ASAP7_75t_SL g2849 ( 
.A(n_2591),
.B(n_1193),
.Y(n_2849)
);

BUFx3_ASAP7_75t_L g2850 ( 
.A(n_2594),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2452),
.B(n_1248),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2514),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2553),
.B(n_1251),
.Y(n_2853)
);

AND2x2_ASAP7_75t_L g2854 ( 
.A(n_2420),
.B(n_1659),
.Y(n_2854)
);

INVx2_ASAP7_75t_SL g2855 ( 
.A(n_2414),
.Y(n_2855)
);

OR2x2_ASAP7_75t_L g2856 ( 
.A(n_2436),
.B(n_1556),
.Y(n_2856)
);

BUFx3_ASAP7_75t_L g2857 ( 
.A(n_2600),
.Y(n_2857)
);

INVx3_ASAP7_75t_SL g2858 ( 
.A(n_2290),
.Y(n_2858)
);

CKINVDCx5p33_ASAP7_75t_R g2859 ( 
.A(n_2572),
.Y(n_2859)
);

INVx3_ASAP7_75t_L g2860 ( 
.A(n_2453),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2413),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2532),
.Y(n_2862)
);

INVx1_ASAP7_75t_SL g2863 ( 
.A(n_2372),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2535),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2536),
.Y(n_2865)
);

INVx4_ASAP7_75t_L g2866 ( 
.A(n_2470),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2538),
.Y(n_2867)
);

INVx3_ASAP7_75t_L g2868 ( 
.A(n_2472),
.Y(n_2868)
);

NOR2xp33_ASAP7_75t_L g2869 ( 
.A(n_2405),
.B(n_1255),
.Y(n_2869)
);

AND2x4_ASAP7_75t_L g2870 ( 
.A(n_2321),
.B(n_1628),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_SL g2871 ( 
.A(n_2554),
.B(n_1256),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2541),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2421),
.B(n_1788),
.Y(n_2873)
);

AND2x2_ASAP7_75t_L g2874 ( 
.A(n_2423),
.B(n_1788),
.Y(n_2874)
);

NOR2xp33_ASAP7_75t_L g2875 ( 
.A(n_2402),
.B(n_1258),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2556),
.B(n_1260),
.Y(n_2876)
);

OAI21xp33_ASAP7_75t_SL g2877 ( 
.A1(n_2428),
.A2(n_1734),
.B(n_1642),
.Y(n_2877)
);

INVx3_ASAP7_75t_L g2878 ( 
.A(n_2473),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2542),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2547),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_SL g2881 ( 
.A(n_2558),
.B(n_1262),
.Y(n_2881)
);

NOR2xp33_ASAP7_75t_L g2882 ( 
.A(n_2440),
.B(n_1263),
.Y(n_2882)
);

BUFx2_ASAP7_75t_L g2883 ( 
.A(n_2307),
.Y(n_2883)
);

NOR2xp33_ASAP7_75t_L g2884 ( 
.A(n_2457),
.B(n_1264),
.Y(n_2884)
);

NOR2xp33_ASAP7_75t_L g2885 ( 
.A(n_2559),
.B(n_2560),
.Y(n_2885)
);

AND2x2_ASAP7_75t_SL g2886 ( 
.A(n_2387),
.B(n_1313),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2550),
.Y(n_2887)
);

INVx4_ASAP7_75t_L g2888 ( 
.A(n_2474),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2551),
.Y(n_2889)
);

INVx4_ASAP7_75t_SL g2890 ( 
.A(n_2525),
.Y(n_2890)
);

AND2x2_ASAP7_75t_L g2891 ( 
.A(n_2374),
.B(n_1788),
.Y(n_2891)
);

NOR2xp33_ASAP7_75t_L g2892 ( 
.A(n_2561),
.B(n_2564),
.Y(n_2892)
);

INVx4_ASAP7_75t_L g2893 ( 
.A(n_2475),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2565),
.B(n_1266),
.Y(n_2894)
);

AND2x2_ASAP7_75t_L g2895 ( 
.A(n_2375),
.B(n_1268),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2468),
.B(n_1272),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2435),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2417),
.Y(n_2898)
);

NOR2xp33_ASAP7_75t_L g2899 ( 
.A(n_2465),
.B(n_1274),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2418),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2444),
.Y(n_2901)
);

BUFx6f_ASAP7_75t_L g2902 ( 
.A(n_2484),
.Y(n_2902)
);

INVx4_ASAP7_75t_L g2903 ( 
.A(n_2485),
.Y(n_2903)
);

BUFx6f_ASAP7_75t_L g2904 ( 
.A(n_2486),
.Y(n_2904)
);

INVx2_ASAP7_75t_SL g2905 ( 
.A(n_2362),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2429),
.Y(n_2906)
);

INVx8_ASAP7_75t_L g2907 ( 
.A(n_2487),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_SL g2908 ( 
.A(n_2379),
.B(n_1280),
.Y(n_2908)
);

BUFx3_ASAP7_75t_L g2909 ( 
.A(n_2604),
.Y(n_2909)
);

INVx4_ASAP7_75t_L g2910 ( 
.A(n_2490),
.Y(n_2910)
);

INVxp33_ASAP7_75t_SL g2911 ( 
.A(n_2326),
.Y(n_2911)
);

AND2x6_ASAP7_75t_L g2912 ( 
.A(n_2449),
.B(n_1596),
.Y(n_2912)
);

BUFx6f_ASAP7_75t_L g2913 ( 
.A(n_2495),
.Y(n_2913)
);

OR2x6_ASAP7_75t_L g2914 ( 
.A(n_2574),
.B(n_1341),
.Y(n_2914)
);

BUFx3_ASAP7_75t_L g2915 ( 
.A(n_2496),
.Y(n_2915)
);

AND2x2_ASAP7_75t_L g2916 ( 
.A(n_2407),
.B(n_1283),
.Y(n_2916)
);

BUFx10_ASAP7_75t_L g2917 ( 
.A(n_2576),
.Y(n_2917)
);

INVxp67_ASAP7_75t_SL g2918 ( 
.A(n_2408),
.Y(n_2918)
);

BUFx3_ASAP7_75t_L g2919 ( 
.A(n_2497),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2454),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2433),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2459),
.Y(n_2922)
);

BUFx4f_ASAP7_75t_L g2923 ( 
.A(n_2328),
.Y(n_2923)
);

OAI22xp33_ASAP7_75t_L g2924 ( 
.A1(n_2369),
.A2(n_1289),
.B1(n_1294),
.B2(n_1285),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2494),
.Y(n_2925)
);

NOR2xp33_ASAP7_75t_L g2926 ( 
.A(n_2419),
.B(n_1296),
.Y(n_2926)
);

INVx6_ASAP7_75t_L g2927 ( 
.A(n_2501),
.Y(n_2927)
);

BUFx2_ASAP7_75t_L g2928 ( 
.A(n_2476),
.Y(n_2928)
);

INVxp67_ASAP7_75t_SL g2929 ( 
.A(n_2534),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2499),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2502),
.Y(n_2931)
);

HB1xp67_ASAP7_75t_L g2932 ( 
.A(n_2363),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_SL g2933 ( 
.A(n_2446),
.B(n_2450),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_SL g2934 ( 
.A(n_2458),
.B(n_1298),
.Y(n_2934)
);

CKINVDCx5p33_ASAP7_75t_R g2935 ( 
.A(n_2579),
.Y(n_2935)
);

INVxp67_ASAP7_75t_L g2936 ( 
.A(n_2503),
.Y(n_2936)
);

INVxp33_ASAP7_75t_L g2937 ( 
.A(n_2477),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_SL g2938 ( 
.A(n_2488),
.B(n_1299),
.Y(n_2938)
);

XOR2x2_ASAP7_75t_L g2939 ( 
.A(n_2361),
.B(n_2367),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2505),
.Y(n_2940)
);

INVx4_ASAP7_75t_L g2941 ( 
.A(n_2504),
.Y(n_2941)
);

BUFx6f_ASAP7_75t_L g2942 ( 
.A(n_2491),
.Y(n_2942)
);

AOI22xp5_ASAP7_75t_L g2943 ( 
.A1(n_2537),
.A2(n_1301),
.B1(n_1302),
.B2(n_1300),
.Y(n_2943)
);

BUFx4f_ASAP7_75t_L g2944 ( 
.A(n_2330),
.Y(n_2944)
);

INVx3_ASAP7_75t_L g2945 ( 
.A(n_2333),
.Y(n_2945)
);

BUFx3_ASAP7_75t_L g2946 ( 
.A(n_2582),
.Y(n_2946)
);

BUFx3_ASAP7_75t_L g2947 ( 
.A(n_2587),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_SL g2948 ( 
.A(n_2493),
.B(n_1304),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2511),
.Y(n_2949)
);

AND2x6_ASAP7_75t_L g2950 ( 
.A(n_2512),
.B(n_1606),
.Y(n_2950)
);

INVx2_ASAP7_75t_SL g2951 ( 
.A(n_2515),
.Y(n_2951)
);

NOR2xp33_ASAP7_75t_L g2952 ( 
.A(n_2521),
.B(n_2527),
.Y(n_2952)
);

NOR2x1p5_ASAP7_75t_L g2953 ( 
.A(n_2595),
.B(n_1307),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2529),
.B(n_1310),
.Y(n_2954)
);

AND2x2_ASAP7_75t_SL g2955 ( 
.A(n_2596),
.B(n_1341),
.Y(n_2955)
);

NAND3x1_ASAP7_75t_L g2956 ( 
.A(n_2359),
.B(n_1196),
.C(n_1195),
.Y(n_2956)
);

BUFx6f_ASAP7_75t_L g2957 ( 
.A(n_2597),
.Y(n_2957)
);

NOR2xp33_ASAP7_75t_L g2958 ( 
.A(n_2599),
.B(n_1316),
.Y(n_2958)
);

AND2x2_ASAP7_75t_L g2959 ( 
.A(n_2601),
.B(n_1319),
.Y(n_2959)
);

BUFx3_ASAP7_75t_L g2960 ( 
.A(n_2606),
.Y(n_2960)
);

INVx2_ASAP7_75t_SL g2961 ( 
.A(n_2608),
.Y(n_2961)
);

INVx2_ASAP7_75t_L g2962 ( 
.A(n_2609),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2610),
.Y(n_2963)
);

BUFx3_ASAP7_75t_L g2964 ( 
.A(n_2611),
.Y(n_2964)
);

INVx3_ASAP7_75t_L g2965 ( 
.A(n_2615),
.Y(n_2965)
);

INVx4_ASAP7_75t_L g2966 ( 
.A(n_2616),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_SL g2967 ( 
.A(n_2381),
.B(n_1324),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_L g2968 ( 
.A(n_2437),
.B(n_1325),
.Y(n_2968)
);

INVx3_ASAP7_75t_L g2969 ( 
.A(n_2593),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2552),
.Y(n_2970)
);

INVx5_ASAP7_75t_L g2971 ( 
.A(n_2593),
.Y(n_2971)
);

INVx4_ASAP7_75t_L g2972 ( 
.A(n_2302),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2562),
.B(n_1327),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2552),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2552),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2357),
.Y(n_2976)
);

CKINVDCx8_ASAP7_75t_R g2977 ( 
.A(n_2302),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_SL g2978 ( 
.A(n_2381),
.B(n_1329),
.Y(n_2978)
);

NOR2xp33_ASAP7_75t_L g2979 ( 
.A(n_2437),
.B(n_1332),
.Y(n_2979)
);

AND2x6_ASAP7_75t_L g2980 ( 
.A(n_2381),
.B(n_1606),
.Y(n_2980)
);

AND2x2_ASAP7_75t_SL g2981 ( 
.A(n_2291),
.B(n_1359),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2357),
.Y(n_2982)
);

CKINVDCx5p33_ASAP7_75t_R g2983 ( 
.A(n_2364),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2357),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_SL g2985 ( 
.A(n_2381),
.B(n_1333),
.Y(n_2985)
);

INVx2_ASAP7_75t_SL g2986 ( 
.A(n_2593),
.Y(n_2986)
);

OAI21xp33_ASAP7_75t_SL g2987 ( 
.A1(n_2562),
.A2(n_1841),
.B(n_1200),
.Y(n_2987)
);

BUFx6f_ASAP7_75t_L g2988 ( 
.A(n_2593),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2357),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2357),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2562),
.B(n_1336),
.Y(n_2991)
);

OAI22xp5_ASAP7_75t_L g2992 ( 
.A1(n_2562),
.A2(n_1340),
.B1(n_1345),
.B2(n_1338),
.Y(n_2992)
);

INVxp67_ASAP7_75t_L g2993 ( 
.A(n_2292),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2552),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2357),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2357),
.Y(n_2996)
);

INVx3_ASAP7_75t_L g2997 ( 
.A(n_2593),
.Y(n_2997)
);

BUFx3_ASAP7_75t_L g2998 ( 
.A(n_2479),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2562),
.B(n_1346),
.Y(n_2999)
);

INVx3_ASAP7_75t_L g3000 ( 
.A(n_2593),
.Y(n_3000)
);

NOR2xp33_ASAP7_75t_L g3001 ( 
.A(n_2437),
.B(n_1348),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2562),
.B(n_1349),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2562),
.B(n_1352),
.Y(n_3003)
);

BUFx6f_ASAP7_75t_L g3004 ( 
.A(n_2593),
.Y(n_3004)
);

INVx3_ASAP7_75t_L g3005 ( 
.A(n_2593),
.Y(n_3005)
);

OR2x2_ASAP7_75t_L g3006 ( 
.A(n_2305),
.B(n_1353),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2357),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_L g3008 ( 
.A(n_2562),
.B(n_1354),
.Y(n_3008)
);

HB1xp67_ASAP7_75t_L g3009 ( 
.A(n_2316),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2562),
.B(n_1358),
.Y(n_3010)
);

HB1xp67_ASAP7_75t_L g3011 ( 
.A(n_2316),
.Y(n_3011)
);

NOR2xp33_ASAP7_75t_SL g3012 ( 
.A(n_2309),
.B(n_1360),
.Y(n_3012)
);

INVx2_ASAP7_75t_L g3013 ( 
.A(n_2552),
.Y(n_3013)
);

NOR2xp33_ASAP7_75t_L g3014 ( 
.A(n_2437),
.B(n_1364),
.Y(n_3014)
);

NOR2xp33_ASAP7_75t_L g3015 ( 
.A(n_2437),
.B(n_1368),
.Y(n_3015)
);

INVx4_ASAP7_75t_L g3016 ( 
.A(n_2302),
.Y(n_3016)
);

INVx3_ASAP7_75t_L g3017 ( 
.A(n_2593),
.Y(n_3017)
);

NAND2x1p5_ASAP7_75t_L g3018 ( 
.A(n_2316),
.B(n_1199),
.Y(n_3018)
);

NOR2xp33_ASAP7_75t_L g3019 ( 
.A(n_2437),
.B(n_1369),
.Y(n_3019)
);

AND2x2_ASAP7_75t_SL g3020 ( 
.A(n_2291),
.B(n_1359),
.Y(n_3020)
);

AND2x2_ASAP7_75t_L g3021 ( 
.A(n_2327),
.B(n_1371),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2562),
.B(n_1379),
.Y(n_3022)
);

INVx2_ASAP7_75t_SL g3023 ( 
.A(n_2593),
.Y(n_3023)
);

INVx2_ASAP7_75t_L g3024 ( 
.A(n_2552),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2357),
.Y(n_3025)
);

OR2x2_ASAP7_75t_L g3026 ( 
.A(n_2305),
.B(n_1380),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2552),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_2552),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2357),
.Y(n_3029)
);

OAI22xp33_ASAP7_75t_L g3030 ( 
.A1(n_2291),
.A2(n_1383),
.B1(n_1386),
.B2(n_1381),
.Y(n_3030)
);

NOR2xp33_ASAP7_75t_R g3031 ( 
.A(n_2309),
.B(n_1391),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2562),
.B(n_1393),
.Y(n_3032)
);

NOR2xp33_ASAP7_75t_L g3033 ( 
.A(n_2437),
.B(n_1403),
.Y(n_3033)
);

OAI22xp5_ASAP7_75t_L g3034 ( 
.A1(n_2741),
.A2(n_1408),
.B1(n_1411),
.B2(n_1405),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2623),
.B(n_1414),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_SL g3036 ( 
.A(n_3018),
.B(n_1415),
.Y(n_3036)
);

NOR2xp33_ASAP7_75t_L g3037 ( 
.A(n_2705),
.B(n_1416),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2623),
.B(n_1417),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2620),
.B(n_3006),
.Y(n_3039)
);

INVxp67_ASAP7_75t_L g3040 ( 
.A(n_3009),
.Y(n_3040)
);

NOR3xp33_ASAP7_75t_L g3041 ( 
.A(n_2682),
.B(n_1206),
.C(n_1201),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_SL g3042 ( 
.A(n_2988),
.B(n_1425),
.Y(n_3042)
);

NOR2xp33_ASAP7_75t_L g3043 ( 
.A(n_2642),
.B(n_2662),
.Y(n_3043)
);

AOI22xp5_ASAP7_75t_L g3044 ( 
.A1(n_2987),
.A2(n_1431),
.B1(n_1434),
.B2(n_1429),
.Y(n_3044)
);

NOR2xp33_ASAP7_75t_L g3045 ( 
.A(n_2668),
.B(n_1440),
.Y(n_3045)
);

NOR2xp33_ASAP7_75t_L g3046 ( 
.A(n_2678),
.B(n_3006),
.Y(n_3046)
);

A2O1A1Ixp33_ASAP7_75t_L g3047 ( 
.A1(n_2650),
.A2(n_1439),
.B(n_1485),
.C(n_1412),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2618),
.B(n_1445),
.Y(n_3048)
);

AND2x2_ASAP7_75t_L g3049 ( 
.A(n_2695),
.B(n_1447),
.Y(n_3049)
);

NAND2x1_ASAP7_75t_L g3050 ( 
.A(n_2980),
.B(n_1606),
.Y(n_3050)
);

AOI22xp5_ASAP7_75t_L g3051 ( 
.A1(n_2637),
.A2(n_1450),
.B1(n_1453),
.B2(n_1449),
.Y(n_3051)
);

NOR2xp33_ASAP7_75t_L g3052 ( 
.A(n_2734),
.B(n_1456),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2638),
.B(n_1457),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_2710),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2715),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2640),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_L g3057 ( 
.A(n_2976),
.B(n_1460),
.Y(n_3057)
);

BUFx2_ASAP7_75t_L g3058 ( 
.A(n_3011),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_2982),
.B(n_1461),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_SL g3060 ( 
.A(n_2988),
.B(n_3004),
.Y(n_3060)
);

INVx2_ASAP7_75t_L g3061 ( 
.A(n_2716),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2984),
.B(n_1464),
.Y(n_3062)
);

INVx2_ASAP7_75t_L g3063 ( 
.A(n_2732),
.Y(n_3063)
);

AOI22xp33_ASAP7_75t_L g3064 ( 
.A1(n_2762),
.A2(n_1468),
.B1(n_1470),
.B2(n_1467),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_2989),
.B(n_1471),
.Y(n_3065)
);

NAND2xp33_ASAP7_75t_L g3066 ( 
.A(n_2707),
.B(n_2718),
.Y(n_3066)
);

NOR2xp33_ASAP7_75t_L g3067 ( 
.A(n_2680),
.B(n_1472),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2990),
.B(n_1478),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2995),
.B(n_1479),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_2996),
.B(n_1481),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_3007),
.B(n_3025),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_3029),
.Y(n_3072)
);

BUFx3_ASAP7_75t_L g3073 ( 
.A(n_3004),
.Y(n_3073)
);

INVx2_ASAP7_75t_SL g3074 ( 
.A(n_2971),
.Y(n_3074)
);

INVx1_ASAP7_75t_SL g3075 ( 
.A(n_2689),
.Y(n_3075)
);

OR2x2_ASAP7_75t_L g3076 ( 
.A(n_2708),
.B(n_1483),
.Y(n_3076)
);

NAND3xp33_ASAP7_75t_L g3077 ( 
.A(n_2877),
.B(n_1688),
.C(n_1606),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_2625),
.B(n_1488),
.Y(n_3078)
);

NOR2xp33_ASAP7_75t_L g3079 ( 
.A(n_2619),
.B(n_1490),
.Y(n_3079)
);

AND2x2_ASAP7_75t_L g3080 ( 
.A(n_2628),
.B(n_1491),
.Y(n_3080)
);

BUFx3_ASAP7_75t_L g3081 ( 
.A(n_2971),
.Y(n_3081)
);

NOR2xp33_ASAP7_75t_L g3082 ( 
.A(n_2993),
.B(n_1498),
.Y(n_3082)
);

BUFx8_ASAP7_75t_SL g3083 ( 
.A(n_2653),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2644),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_2649),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2775),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2622),
.B(n_1501),
.Y(n_3087)
);

INVx8_ASAP7_75t_L g3088 ( 
.A(n_2907),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_3021),
.B(n_1502),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2756),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_2781),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_3026),
.B(n_1503),
.Y(n_3092)
);

NOR2xp33_ASAP7_75t_L g3093 ( 
.A(n_2762),
.B(n_1505),
.Y(n_3093)
);

AOI22xp33_ASAP7_75t_L g3094 ( 
.A1(n_2629),
.A2(n_1513),
.B1(n_1517),
.B2(n_1511),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2973),
.B(n_1519),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_2991),
.B(n_1524),
.Y(n_3096)
);

BUFx5_ASAP7_75t_L g3097 ( 
.A(n_2980),
.Y(n_3097)
);

AND2x2_ASAP7_75t_L g3098 ( 
.A(n_2630),
.B(n_1526),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_2999),
.B(n_1528),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_3002),
.B(n_1534),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2780),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_3003),
.B(n_1535),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_2784),
.Y(n_3103)
);

INVx2_ASAP7_75t_SL g3104 ( 
.A(n_2907),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_SL g3105 ( 
.A(n_3012),
.B(n_1539),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_3008),
.B(n_1544),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_SL g3107 ( 
.A(n_2690),
.B(n_1545),
.Y(n_3107)
);

AOI22xp33_ASAP7_75t_L g3108 ( 
.A1(n_2629),
.A2(n_2666),
.B1(n_2809),
.B2(n_2895),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_3010),
.B(n_1546),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_2659),
.Y(n_3110)
);

INVx2_ASAP7_75t_SL g3111 ( 
.A(n_2927),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_3022),
.B(n_1548),
.Y(n_3112)
);

INVx3_ASAP7_75t_L g3113 ( 
.A(n_2634),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_SL g3114 ( 
.A(n_2729),
.B(n_1552),
.Y(n_3114)
);

NOR2xp33_ASAP7_75t_L g3115 ( 
.A(n_2869),
.B(n_1553),
.Y(n_3115)
);

NOR2xp33_ASAP7_75t_L g3116 ( 
.A(n_2809),
.B(n_1560),
.Y(n_3116)
);

AOI22xp5_ASAP7_75t_L g3117 ( 
.A1(n_2691),
.A2(n_1563),
.B1(n_1565),
.B2(n_1562),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_3032),
.B(n_1566),
.Y(n_3118)
);

AOI22xp33_ASAP7_75t_L g3119 ( 
.A1(n_2844),
.A2(n_1572),
.B1(n_1575),
.B2(n_1570),
.Y(n_3119)
);

NAND2xp33_ASAP7_75t_L g3120 ( 
.A(n_2707),
.B(n_1578),
.Y(n_3120)
);

NOR2xp67_ASAP7_75t_SL g3121 ( 
.A(n_2977),
.B(n_1586),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2655),
.B(n_1588),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_2663),
.Y(n_3123)
);

AOI22xp5_ASAP7_75t_L g3124 ( 
.A1(n_2691),
.A2(n_1593),
.B1(n_1595),
.B2(n_1590),
.Y(n_3124)
);

INVx8_ASAP7_75t_L g3125 ( 
.A(n_2741),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2658),
.B(n_1597),
.Y(n_3126)
);

INVx2_ASAP7_75t_SL g3127 ( 
.A(n_2927),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2669),
.Y(n_3128)
);

INVx8_ASAP7_75t_L g3129 ( 
.A(n_2787),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2671),
.Y(n_3130)
);

INVx2_ASAP7_75t_SL g3131 ( 
.A(n_2664),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_2719),
.B(n_1599),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2675),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2670),
.B(n_1609),
.Y(n_3134)
);

BUFx8_ASAP7_75t_SL g3135 ( 
.A(n_2627),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_2676),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_SL g3137 ( 
.A(n_2626),
.B(n_1610),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_2684),
.B(n_1612),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_2968),
.B(n_1613),
.Y(n_3139)
);

NOR2xp33_ASAP7_75t_SL g3140 ( 
.A(n_2980),
.B(n_1614),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2979),
.B(n_1615),
.Y(n_3141)
);

BUFx8_ASAP7_75t_L g3142 ( 
.A(n_2957),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2686),
.Y(n_3143)
);

INVxp67_ASAP7_75t_SL g3144 ( 
.A(n_2677),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2687),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_SL g3146 ( 
.A(n_2986),
.B(n_1621),
.Y(n_3146)
);

AND2x6_ASAP7_75t_SL g3147 ( 
.A(n_2722),
.B(n_2633),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_SL g3148 ( 
.A(n_3023),
.B(n_1622),
.Y(n_3148)
);

NOR2xp33_ASAP7_75t_L g3149 ( 
.A(n_2654),
.B(n_1623),
.Y(n_3149)
);

OR2x2_ASAP7_75t_L g3150 ( 
.A(n_2700),
.B(n_1624),
.Y(n_3150)
);

NOR2xp33_ASAP7_75t_L g3151 ( 
.A(n_2875),
.B(n_1625),
.Y(n_3151)
);

OR2x6_ASAP7_75t_L g3152 ( 
.A(n_2787),
.B(n_2685),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2688),
.Y(n_3153)
);

INVx2_ASAP7_75t_L g3154 ( 
.A(n_2694),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_3001),
.B(n_1626),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_2703),
.Y(n_3156)
);

NOR2xp33_ASAP7_75t_L g3157 ( 
.A(n_2891),
.B(n_1630),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2709),
.Y(n_3158)
);

AOI221xp5_ASAP7_75t_L g3159 ( 
.A1(n_2766),
.A2(n_1639),
.B1(n_1643),
.B2(n_1632),
.C(n_1631),
.Y(n_3159)
);

O2A1O1Ixp33_ASAP7_75t_L g3160 ( 
.A1(n_2731),
.A2(n_1216),
.B(n_1230),
.C(n_1213),
.Y(n_3160)
);

INVx2_ASAP7_75t_L g3161 ( 
.A(n_2717),
.Y(n_3161)
);

INVx2_ASAP7_75t_SL g3162 ( 
.A(n_2699),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_3014),
.B(n_1648),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_SL g3164 ( 
.A(n_2885),
.B(n_1649),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_3015),
.B(n_1652),
.Y(n_3165)
);

CKINVDCx5p33_ASAP7_75t_R g3166 ( 
.A(n_2795),
.Y(n_3166)
);

BUFx3_ASAP7_75t_L g3167 ( 
.A(n_2902),
.Y(n_3167)
);

OAI22x1_ASAP7_75t_R g3168 ( 
.A1(n_2727),
.A2(n_1656),
.B1(n_1661),
.B2(n_1655),
.Y(n_3168)
);

INVx8_ASAP7_75t_L g3169 ( 
.A(n_2691),
.Y(n_3169)
);

INVx8_ASAP7_75t_L g3170 ( 
.A(n_2902),
.Y(n_3170)
);

AND2x2_ASAP7_75t_L g3171 ( 
.A(n_2713),
.B(n_1662),
.Y(n_3171)
);

AND2x4_ASAP7_75t_L g3172 ( 
.A(n_2631),
.B(n_2969),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2720),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_3019),
.B(n_1669),
.Y(n_3174)
);

AOI22xp5_ASAP7_75t_L g3175 ( 
.A1(n_2790),
.A2(n_1674),
.B1(n_1676),
.B2(n_1672),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_3033),
.B(n_1680),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_2723),
.Y(n_3177)
);

INVx2_ASAP7_75t_SL g3178 ( 
.A(n_2759),
.Y(n_3178)
);

INVx2_ASAP7_75t_SL g3179 ( 
.A(n_2826),
.Y(n_3179)
);

NOR2xp33_ASAP7_75t_L g3180 ( 
.A(n_2856),
.B(n_1685),
.Y(n_3180)
);

INVx8_ASAP7_75t_L g3181 ( 
.A(n_2904),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_SL g3182 ( 
.A(n_2892),
.B(n_1686),
.Y(n_3182)
);

INVx2_ASAP7_75t_SL g3183 ( 
.A(n_2998),
.Y(n_3183)
);

AND2x4_ASAP7_75t_L g3184 ( 
.A(n_2997),
.B(n_1235),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_SL g3185 ( 
.A(n_3030),
.B(n_1690),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2724),
.Y(n_3186)
);

AOI22xp33_ASAP7_75t_SL g3187 ( 
.A1(n_2807),
.A2(n_1691),
.B1(n_1707),
.B2(n_1696),
.Y(n_3187)
);

INVx2_ASAP7_75t_L g3188 ( 
.A(n_2726),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_2992),
.B(n_1711),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_2636),
.B(n_2776),
.Y(n_3190)
);

NOR2xp33_ASAP7_75t_L g3191 ( 
.A(n_2856),
.B(n_1712),
.Y(n_3191)
);

NOR2xp33_ASAP7_75t_L g3192 ( 
.A(n_2700),
.B(n_1714),
.Y(n_3192)
);

BUFx6f_ASAP7_75t_L g3193 ( 
.A(n_2753),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2735),
.Y(n_3194)
);

NOR2xp33_ASAP7_75t_L g3195 ( 
.A(n_2701),
.B(n_1717),
.Y(n_3195)
);

BUFx3_ASAP7_75t_L g3196 ( 
.A(n_2904),
.Y(n_3196)
);

NOR2xp33_ASAP7_75t_L g3197 ( 
.A(n_2778),
.B(n_1723),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_2725),
.B(n_1724),
.Y(n_3198)
);

INVx2_ASAP7_75t_L g3199 ( 
.A(n_2739),
.Y(n_3199)
);

NOR3xp33_ASAP7_75t_L g3200 ( 
.A(n_2792),
.B(n_1241),
.C(n_1239),
.Y(n_3200)
);

O2A1O1Ixp33_ASAP7_75t_L g3201 ( 
.A1(n_2665),
.A2(n_1249),
.B(n_1257),
.C(n_1246),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_SL g3202 ( 
.A(n_2639),
.B(n_1727),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2750),
.Y(n_3203)
);

O2A1O1Ixp33_ASAP7_75t_L g3204 ( 
.A1(n_2696),
.A2(n_2641),
.B(n_2846),
.C(n_2824),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_2648),
.B(n_1730),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_2796),
.Y(n_3206)
);

AND2x6_ASAP7_75t_SL g3207 ( 
.A(n_2914),
.B(n_1259),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_2737),
.B(n_1731),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_L g3209 ( 
.A(n_2846),
.B(n_1733),
.Y(n_3209)
);

BUFx12f_ASAP7_75t_L g3210 ( 
.A(n_2714),
.Y(n_3210)
);

NAND3xp33_ASAP7_75t_L g3211 ( 
.A(n_2830),
.B(n_1716),
.C(n_1688),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_SL g3212 ( 
.A(n_2758),
.B(n_1737),
.Y(n_3212)
);

NOR2xp33_ASAP7_75t_L g3213 ( 
.A(n_2742),
.B(n_1738),
.Y(n_3213)
);

OAI22xp5_ASAP7_75t_L g3214 ( 
.A1(n_2886),
.A2(n_1740),
.B1(n_1741),
.B2(n_1739),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_L g3215 ( 
.A(n_2823),
.B(n_1744),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_SL g3216 ( 
.A(n_3000),
.B(n_1748),
.Y(n_3216)
);

NOR2xp33_ASAP7_75t_L g3217 ( 
.A(n_2818),
.B(n_1751),
.Y(n_3217)
);

NOR2xp33_ASAP7_75t_L g3218 ( 
.A(n_2777),
.B(n_1752),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_2746),
.B(n_1755),
.Y(n_3219)
);

AOI21xp5_ASAP7_75t_L g3220 ( 
.A1(n_2744),
.A2(n_1270),
.B(n_1269),
.Y(n_3220)
);

NOR2xp33_ASAP7_75t_L g3221 ( 
.A(n_2854),
.B(n_1757),
.Y(n_3221)
);

NOR2xp33_ASAP7_75t_L g3222 ( 
.A(n_2873),
.B(n_1760),
.Y(n_3222)
);

NOR2xp33_ASAP7_75t_L g3223 ( 
.A(n_2874),
.B(n_2908),
.Y(n_3223)
);

NOR2xp33_ASAP7_75t_L g3224 ( 
.A(n_2782),
.B(n_1763),
.Y(n_3224)
);

INVx2_ASAP7_75t_L g3225 ( 
.A(n_2794),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2798),
.Y(n_3226)
);

NAND2x1p5_ASAP7_75t_L g3227 ( 
.A(n_2693),
.B(n_2736),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_L g3228 ( 
.A(n_2747),
.B(n_1764),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2802),
.Y(n_3229)
);

NOR3x1_ASAP7_75t_L g3230 ( 
.A(n_2928),
.B(n_1284),
.C(n_1277),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_2760),
.B(n_1771),
.Y(n_3231)
);

A2O1A1Ixp33_ASAP7_75t_L g3232 ( 
.A1(n_2757),
.A2(n_1439),
.B(n_1485),
.C(n_1412),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_2754),
.Y(n_3233)
);

OAI21xp5_ASAP7_75t_L g3234 ( 
.A1(n_2752),
.A2(n_1290),
.B(n_1287),
.Y(n_3234)
);

NOR3xp33_ASAP7_75t_L g3235 ( 
.A(n_2797),
.B(n_1295),
.C(n_1291),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_L g3236 ( 
.A(n_2771),
.B(n_1775),
.Y(n_3236)
);

O2A1O1Ixp5_ASAP7_75t_L g3237 ( 
.A1(n_2831),
.A2(n_1500),
.B(n_1540),
.C(n_1499),
.Y(n_3237)
);

AOI22xp33_ASAP7_75t_L g3238 ( 
.A1(n_2981),
.A2(n_1776),
.B1(n_1781),
.B2(n_1777),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_2768),
.Y(n_3239)
);

NOR2xp33_ASAP7_75t_L g3240 ( 
.A(n_2783),
.B(n_1782),
.Y(n_3240)
);

AOI22xp5_ASAP7_75t_L g3241 ( 
.A1(n_3020),
.A2(n_1784),
.B1(n_1786),
.B2(n_1783),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_2817),
.B(n_1787),
.Y(n_3242)
);

AOI21xp5_ASAP7_75t_L g3243 ( 
.A1(n_2803),
.A2(n_1305),
.B(n_1297),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_SL g3244 ( 
.A(n_3005),
.B(n_1791),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_2828),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_2839),
.B(n_2842),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2852),
.Y(n_3247)
);

INVx2_ASAP7_75t_SL g3248 ( 
.A(n_2913),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_2753),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_2954),
.Y(n_3250)
);

OAI22xp5_ASAP7_75t_SL g3251 ( 
.A1(n_2849),
.A2(n_1795),
.B1(n_1796),
.B2(n_1794),
.Y(n_3251)
);

AND2x2_ASAP7_75t_L g3252 ( 
.A(n_2916),
.B(n_1797),
.Y(n_3252)
);

INVx2_ASAP7_75t_L g3253 ( 
.A(n_2897),
.Y(n_3253)
);

AND2x2_ASAP7_75t_L g3254 ( 
.A(n_2800),
.B(n_1800),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_2847),
.B(n_1801),
.Y(n_3255)
);

AOI22xp5_ASAP7_75t_L g3256 ( 
.A1(n_2918),
.A2(n_1806),
.B1(n_1809),
.B2(n_1804),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_2943),
.B(n_1810),
.Y(n_3257)
);

AND2x2_ASAP7_75t_L g3258 ( 
.A(n_2926),
.B(n_2955),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_2820),
.Y(n_3259)
);

INVx2_ASAP7_75t_L g3260 ( 
.A(n_2901),
.Y(n_3260)
);

NOR2xp33_ASAP7_75t_L g3261 ( 
.A(n_2805),
.B(n_1812),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_SL g3262 ( 
.A(n_3017),
.B(n_1815),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_2808),
.B(n_1820),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_2920),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_L g3265 ( 
.A(n_2841),
.B(n_1827),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_2922),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_SL g3267 ( 
.A(n_2738),
.B(n_1830),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_2853),
.B(n_1835),
.Y(n_3268)
);

AOI22xp5_ASAP7_75t_L g3269 ( 
.A1(n_2862),
.A2(n_1838),
.B1(n_1842),
.B2(n_1837),
.Y(n_3269)
);

AOI21xp5_ASAP7_75t_L g3270 ( 
.A1(n_2933),
.A2(n_1328),
.B(n_1326),
.Y(n_3270)
);

AOI22xp33_ASAP7_75t_L g3271 ( 
.A1(n_2882),
.A2(n_1843),
.B1(n_1847),
.B2(n_1846),
.Y(n_3271)
);

OR2x2_ASAP7_75t_L g3272 ( 
.A(n_2929),
.B(n_1850),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_L g3273 ( 
.A(n_2876),
.B(n_1852),
.Y(n_3273)
);

BUFx8_ASAP7_75t_L g3274 ( 
.A(n_2957),
.Y(n_3274)
);

HB1xp67_ASAP7_75t_L g3275 ( 
.A(n_2786),
.Y(n_3275)
);

NOR2xp33_ASAP7_75t_L g3276 ( 
.A(n_2789),
.B(n_1853),
.Y(n_3276)
);

INVxp67_ASAP7_75t_L g3277 ( 
.A(n_2814),
.Y(n_3277)
);

OR2x2_ASAP7_75t_L g3278 ( 
.A(n_2698),
.B(n_2702),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_2894),
.B(n_1854),
.Y(n_3279)
);

INVxp67_ASAP7_75t_L g3280 ( 
.A(n_2816),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2749),
.B(n_1859),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_SL g3282 ( 
.A(n_3031),
.B(n_1860),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_SL g3283 ( 
.A(n_2791),
.B(n_1861),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_2925),
.Y(n_3284)
);

NOR2xp33_ASAP7_75t_L g3285 ( 
.A(n_2864),
.B(n_1869),
.Y(n_3285)
);

AOI21xp5_ASAP7_75t_L g3286 ( 
.A1(n_2624),
.A2(n_1339),
.B(n_1331),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_2930),
.Y(n_3287)
);

INVx2_ASAP7_75t_L g3288 ( 
.A(n_2931),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_SL g3289 ( 
.A(n_2697),
.B(n_1871),
.Y(n_3289)
);

INVxp33_ASAP7_75t_L g3290 ( 
.A(n_2870),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_2940),
.Y(n_3291)
);

AND2x4_ASAP7_75t_L g3292 ( 
.A(n_2799),
.B(n_1342),
.Y(n_3292)
);

BUFx8_ASAP7_75t_L g3293 ( 
.A(n_2883),
.Y(n_3293)
);

INVx2_ASAP7_75t_L g3294 ( 
.A(n_2811),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_2812),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_2865),
.B(n_1876),
.Y(n_3296)
);

NOR2xp67_ASAP7_75t_L g3297 ( 
.A(n_2621),
.B(n_245),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_2867),
.B(n_1878),
.Y(n_3298)
);

INVx8_ASAP7_75t_L g3299 ( 
.A(n_2913),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_2815),
.Y(n_3300)
);

INVx2_ASAP7_75t_L g3301 ( 
.A(n_2634),
.Y(n_3301)
);

INVxp67_ASAP7_75t_L g3302 ( 
.A(n_2751),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_2872),
.B(n_1880),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_2681),
.Y(n_3304)
);

OR2x2_ASAP7_75t_L g3305 ( 
.A(n_2730),
.B(n_2793),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_SL g3306 ( 
.A(n_2983),
.B(n_1881),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_2879),
.B(n_1883),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_SL g3308 ( 
.A(n_2643),
.B(n_1174),
.Y(n_3308)
);

OR2x6_ASAP7_75t_L g3309 ( 
.A(n_2972),
.B(n_1499),
.Y(n_3309)
);

AOI22xp5_ASAP7_75t_L g3310 ( 
.A1(n_2880),
.A2(n_1343),
.B1(n_1350),
.B2(n_1344),
.Y(n_3310)
);

O2A1O1Ixp5_ASAP7_75t_L g3311 ( 
.A1(n_2967),
.A2(n_1540),
.B(n_1636),
.C(n_1500),
.Y(n_3311)
);

OR2x2_ASAP7_75t_L g3312 ( 
.A(n_2679),
.B(n_1356),
.Y(n_3312)
);

NOR2xp33_ASAP7_75t_L g3313 ( 
.A(n_2887),
.B(n_1365),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_2889),
.B(n_1370),
.Y(n_3314)
);

OR2x2_ASAP7_75t_L g3315 ( 
.A(n_2863),
.B(n_1375),
.Y(n_3315)
);

INVx2_ASAP7_75t_L g3316 ( 
.A(n_2643),
.Y(n_3316)
);

INVx4_ASAP7_75t_L g3317 ( 
.A(n_2693),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_2728),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_2832),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_L g3320 ( 
.A(n_2851),
.B(n_1388),
.Y(n_3320)
);

INVx2_ASAP7_75t_SL g3321 ( 
.A(n_2915),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_SL g3322 ( 
.A(n_2896),
.B(n_1174),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_2740),
.B(n_1389),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_2764),
.Y(n_3324)
);

NOR2xp33_ASAP7_75t_L g3325 ( 
.A(n_2745),
.B(n_1390),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_2934),
.Y(n_3326)
);

AOI21xp5_ASAP7_75t_L g3327 ( 
.A1(n_2632),
.A2(n_1399),
.B(n_1395),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_2924),
.B(n_2884),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_SL g3329 ( 
.A(n_2736),
.B(n_1174),
.Y(n_3329)
);

AOI22xp5_ASAP7_75t_L g3330 ( 
.A1(n_2673),
.A2(n_1401),
.B1(n_1410),
.B2(n_1404),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_2938),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_2899),
.B(n_1413),
.Y(n_3332)
);

NOR3x1_ASAP7_75t_L g3333 ( 
.A(n_2674),
.B(n_1833),
.C(n_1829),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_SL g3334 ( 
.A(n_2651),
.B(n_1355),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_2683),
.B(n_1418),
.Y(n_3335)
);

AND2x4_ASAP7_75t_L g3336 ( 
.A(n_2799),
.B(n_1419),
.Y(n_3336)
);

NOR2xp33_ASAP7_75t_SL g3337 ( 
.A(n_2707),
.B(n_1584),
.Y(n_3337)
);

AOI22xp33_ASAP7_75t_L g3338 ( 
.A1(n_2833),
.A2(n_1584),
.B1(n_1421),
.B2(n_1427),
.Y(n_3338)
);

NOR2xp33_ASAP7_75t_L g3339 ( 
.A(n_2813),
.B(n_1423),
.Y(n_3339)
);

INVx2_ASAP7_75t_L g3340 ( 
.A(n_2837),
.Y(n_3340)
);

INVx2_ASAP7_75t_L g3341 ( 
.A(n_2848),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_2948),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_L g3343 ( 
.A(n_2834),
.B(n_1428),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_2871),
.B(n_1436),
.Y(n_3344)
);

INVx2_ASAP7_75t_L g3345 ( 
.A(n_2861),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_SL g3346 ( 
.A(n_2651),
.B(n_1355),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_2978),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_2898),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_2881),
.B(n_2845),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_2985),
.Y(n_3350)
);

INVx2_ASAP7_75t_SL g3351 ( 
.A(n_2919),
.Y(n_3351)
);

OR2x2_ASAP7_75t_L g3352 ( 
.A(n_2748),
.B(n_1442),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_SL g3353 ( 
.A(n_2652),
.B(n_1355),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_SL g3354 ( 
.A(n_2652),
.B(n_1355),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_SL g3355 ( 
.A(n_2657),
.B(n_1508),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_SL g3356 ( 
.A(n_2657),
.B(n_1508),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_L g3357 ( 
.A(n_2733),
.B(n_1446),
.Y(n_3357)
);

INVx2_ASAP7_75t_L g3358 ( 
.A(n_2900),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_SL g3359 ( 
.A(n_2646),
.B(n_1508),
.Y(n_3359)
);

AND2x2_ASAP7_75t_L g3360 ( 
.A(n_2959),
.B(n_1448),
.Y(n_3360)
);

INVx2_ASAP7_75t_SL g3361 ( 
.A(n_2835),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_SL g3362 ( 
.A(n_2661),
.B(n_2770),
.Y(n_3362)
);

O2A1O1Ixp33_ASAP7_75t_L g3363 ( 
.A1(n_2785),
.A2(n_1463),
.B(n_1465),
.C(n_1462),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_2704),
.B(n_1475),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_SL g3365 ( 
.A(n_2712),
.B(n_1508),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_2761),
.B(n_1476),
.Y(n_3366)
);

INVx2_ASAP7_75t_L g3367 ( 
.A(n_2906),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_SL g3368 ( 
.A(n_2855),
.B(n_1617),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_2761),
.B(n_1477),
.Y(n_3369)
);

BUFx6f_ASAP7_75t_L g3370 ( 
.A(n_2763),
.Y(n_3370)
);

AOI22xp5_ASAP7_75t_L g3371 ( 
.A1(n_2838),
.A2(n_1489),
.B1(n_1492),
.B2(n_1487),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_L g3372 ( 
.A(n_2843),
.B(n_2868),
.Y(n_3372)
);

INVxp67_ASAP7_75t_L g3373 ( 
.A(n_2932),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_2773),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_SL g3375 ( 
.A(n_2660),
.B(n_1617),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_2843),
.B(n_1493),
.Y(n_3376)
);

INVx2_ASAP7_75t_L g3377 ( 
.A(n_2921),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_SL g3378 ( 
.A(n_2660),
.B(n_1617),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_2949),
.Y(n_3379)
);

INVx2_ASAP7_75t_L g3380 ( 
.A(n_2656),
.Y(n_3380)
);

NOR2xp33_ASAP7_75t_L g3381 ( 
.A(n_2911),
.B(n_1496),
.Y(n_3381)
);

AOI22xp33_ASAP7_75t_L g3382 ( 
.A1(n_2958),
.A2(n_1584),
.B1(n_1512),
.B2(n_1520),
.Y(n_3382)
);

INVxp67_ASAP7_75t_L g3383 ( 
.A(n_2914),
.Y(n_3383)
);

NOR2xp67_ASAP7_75t_L g3384 ( 
.A(n_3016),
.B(n_245),
.Y(n_3384)
);

INVx5_ASAP7_75t_L g3385 ( 
.A(n_2819),
.Y(n_3385)
);

NOR2xp33_ASAP7_75t_L g3386 ( 
.A(n_2936),
.B(n_1510),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_2672),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_2878),
.B(n_1529),
.Y(n_3388)
);

NOR3xp33_ASAP7_75t_L g3389 ( 
.A(n_2963),
.B(n_1882),
.C(n_1875),
.Y(n_3389)
);

NOR2xp33_ASAP7_75t_L g3390 ( 
.A(n_2779),
.B(n_1530),
.Y(n_3390)
);

OAI22x1_ASAP7_75t_L g3391 ( 
.A1(n_2953),
.A2(n_1533),
.B1(n_1537),
.B2(n_1531),
.Y(n_3391)
);

INVx2_ASAP7_75t_L g3392 ( 
.A(n_2692),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_2706),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_2788),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_2801),
.Y(n_3395)
);

AOI21xp5_ASAP7_75t_L g3396 ( 
.A1(n_2970),
.A2(n_1549),
.B(n_1541),
.Y(n_3396)
);

INVxp67_ASAP7_75t_SL g3397 ( 
.A(n_2905),
.Y(n_3397)
);

AND2x4_ASAP7_75t_L g3398 ( 
.A(n_2890),
.B(n_1554),
.Y(n_3398)
);

OAI221xp5_ASAP7_75t_L g3399 ( 
.A1(n_2961),
.A2(n_1684),
.B1(n_1721),
.B2(n_1607),
.C(n_1568),
.Y(n_3399)
);

INVx2_ASAP7_75t_L g3400 ( 
.A(n_2974),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_2667),
.B(n_1559),
.Y(n_3401)
);

OR2x2_ASAP7_75t_L g3402 ( 
.A(n_2822),
.B(n_1571),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_SL g3403 ( 
.A(n_2763),
.B(n_1617),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_2743),
.B(n_1573),
.Y(n_3404)
);

O2A1O1Ixp33_ASAP7_75t_L g3405 ( 
.A1(n_2962),
.A2(n_1576),
.B(n_1579),
.C(n_1574),
.Y(n_3405)
);

NAND2x1_ASAP7_75t_L g3406 ( 
.A(n_2819),
.B(n_1688),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_2635),
.B(n_1582),
.Y(n_3407)
);

AND2x6_ASAP7_75t_SL g3408 ( 
.A(n_2711),
.B(n_1825),
.Y(n_3408)
);

OAI22xp5_ASAP7_75t_L g3409 ( 
.A1(n_2951),
.A2(n_1645),
.B1(n_1664),
.B2(n_1636),
.Y(n_3409)
);

BUFx2_ASAP7_75t_L g3410 ( 
.A(n_2866),
.Y(n_3410)
);

AND2x2_ASAP7_75t_L g3411 ( 
.A(n_2890),
.B(n_2888),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_SL g3412 ( 
.A(n_2772),
.B(n_2806),
.Y(n_3412)
);

AOI21xp5_ASAP7_75t_L g3413 ( 
.A1(n_2975),
.A2(n_1585),
.B(n_1583),
.Y(n_3413)
);

NOR2x1p5_ASAP7_75t_L g3414 ( 
.A(n_2836),
.B(n_1839),
.Y(n_3414)
);

NAND3xp33_ASAP7_75t_SL g3415 ( 
.A(n_2840),
.B(n_1589),
.C(n_1587),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_2893),
.B(n_1591),
.Y(n_3416)
);

NAND3xp33_ASAP7_75t_L g3417 ( 
.A(n_2952),
.B(n_1716),
.C(n_1688),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_L g3418 ( 
.A(n_2903),
.B(n_1592),
.Y(n_3418)
);

AND2x2_ASAP7_75t_L g3419 ( 
.A(n_2910),
.B(n_1594),
.Y(n_3419)
);

O2A1O1Ixp5_ASAP7_75t_L g3420 ( 
.A1(n_2994),
.A2(n_1664),
.B(n_1671),
.C(n_1645),
.Y(n_3420)
);

INVx2_ASAP7_75t_L g3421 ( 
.A(n_3013),
.Y(n_3421)
);

INVx2_ASAP7_75t_L g3422 ( 
.A(n_3024),
.Y(n_3422)
);

BUFx6f_ASAP7_75t_L g3423 ( 
.A(n_2772),
.Y(n_3423)
);

INVx2_ASAP7_75t_L g3424 ( 
.A(n_3027),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_2941),
.B(n_1604),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_2810),
.B(n_1611),
.Y(n_3426)
);

INVx2_ASAP7_75t_L g3427 ( 
.A(n_3028),
.Y(n_3427)
);

INVx3_ASAP7_75t_L g3428 ( 
.A(n_2806),
.Y(n_3428)
);

OR2x2_ASAP7_75t_L g3429 ( 
.A(n_2829),
.B(n_1618),
.Y(n_3429)
);

BUFx3_ASAP7_75t_L g3430 ( 
.A(n_2850),
.Y(n_3430)
);

O2A1O1Ixp33_ASAP7_75t_L g3431 ( 
.A1(n_2765),
.A2(n_1620),
.B(n_1629),
.C(n_1627),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_L g3432 ( 
.A(n_2645),
.B(n_1635),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_SL g3433 ( 
.A(n_2923),
.B(n_1584),
.Y(n_3433)
);

OAI22xp33_ASAP7_75t_L g3434 ( 
.A1(n_2944),
.A2(n_1644),
.B1(n_1646),
.B2(n_1641),
.Y(n_3434)
);

AND2x4_ASAP7_75t_L g3435 ( 
.A(n_2647),
.B(n_1647),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_2819),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_SL g3437 ( 
.A(n_2945),
.B(n_1584),
.Y(n_3437)
);

BUFx6f_ASAP7_75t_L g3438 ( 
.A(n_2718),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_2860),
.B(n_1650),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_2718),
.B(n_1663),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_2721),
.B(n_1667),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_L g3442 ( 
.A(n_2721),
.B(n_1670),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_2721),
.B(n_1673),
.Y(n_3443)
);

OR2x2_ASAP7_75t_L g3444 ( 
.A(n_2857),
.B(n_1675),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_2937),
.B(n_1713),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_SL g3446 ( 
.A(n_2942),
.B(n_1584),
.Y(n_3446)
);

AND2x2_ASAP7_75t_SL g3447 ( 
.A(n_2966),
.B(n_1671),
.Y(n_3447)
);

AOI21xp5_ASAP7_75t_L g3448 ( 
.A1(n_2821),
.A2(n_1725),
.B(n_1722),
.Y(n_3448)
);

AO22x1_ASAP7_75t_L g3449 ( 
.A1(n_2859),
.A2(n_1834),
.B1(n_1844),
.B2(n_1826),
.Y(n_3449)
);

AOI22xp5_ASAP7_75t_L g3450 ( 
.A1(n_2956),
.A2(n_1726),
.B1(n_1735),
.B2(n_1728),
.Y(n_3450)
);

NOR3xp33_ASAP7_75t_L g3451 ( 
.A(n_2965),
.B(n_1858),
.C(n_1857),
.Y(n_3451)
);

OAI22xp33_ASAP7_75t_L g3452 ( 
.A1(n_2858),
.A2(n_1747),
.B1(n_1756),
.B2(n_1742),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_2825),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_L g3454 ( 
.A(n_2755),
.B(n_1758),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_SL g3455 ( 
.A(n_2942),
.B(n_1584),
.Y(n_3455)
);

BUFx6f_ASAP7_75t_SL g3456 ( 
.A(n_2909),
.Y(n_3456)
);

INVx2_ASAP7_75t_L g3457 ( 
.A(n_2755),
.Y(n_3457)
);

INVxp67_ASAP7_75t_L g3458 ( 
.A(n_2964),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_2755),
.B(n_1759),
.Y(n_3459)
);

NAND2xp5_ASAP7_75t_L g3460 ( 
.A(n_2767),
.B(n_1768),
.Y(n_3460)
);

BUFx3_ASAP7_75t_L g3461 ( 
.A(n_2946),
.Y(n_3461)
);

HB1xp67_ASAP7_75t_L g3462 ( 
.A(n_2947),
.Y(n_3462)
);

AND2x2_ASAP7_75t_L g3463 ( 
.A(n_2939),
.B(n_1769),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_2804),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_2804),
.Y(n_3465)
);

NOR2xp67_ASAP7_75t_SL g3466 ( 
.A(n_2960),
.B(n_1716),
.Y(n_3466)
);

INVx1_ASAP7_75t_L g3467 ( 
.A(n_2804),
.Y(n_3467)
);

AND2x2_ASAP7_75t_L g3468 ( 
.A(n_2935),
.B(n_1774),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_2767),
.Y(n_3469)
);

AOI22xp33_ASAP7_75t_L g3470 ( 
.A1(n_2767),
.A2(n_1779),
.B1(n_1789),
.B2(n_1778),
.Y(n_3470)
);

O2A1O1Ixp33_ASAP7_75t_L g3471 ( 
.A1(n_2917),
.A2(n_1798),
.B(n_1803),
.C(n_1792),
.Y(n_3471)
);

AOI22xp33_ASAP7_75t_L g3472 ( 
.A1(n_2769),
.A2(n_1808),
.B1(n_1811),
.B2(n_1805),
.Y(n_3472)
);

INVxp67_ASAP7_75t_L g3473 ( 
.A(n_2769),
.Y(n_3473)
);

NOR2xp33_ASAP7_75t_L g3474 ( 
.A(n_2769),
.B(n_1821),
.Y(n_3474)
);

INVx3_ASAP7_75t_L g3475 ( 
.A(n_2774),
.Y(n_3475)
);

OAI22xp5_ASAP7_75t_L g3476 ( 
.A1(n_2774),
.A2(n_1682),
.B1(n_1687),
.B2(n_1678),
.Y(n_3476)
);

NOR2xp33_ASAP7_75t_L g3477 ( 
.A(n_2774),
.B(n_1824),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_2950),
.Y(n_3478)
);

NAND3xp33_ASAP7_75t_L g3479 ( 
.A(n_2827),
.B(n_1732),
.C(n_1716),
.Y(n_3479)
);

INVx4_ASAP7_75t_L g3480 ( 
.A(n_2827),
.Y(n_3480)
);

AND2x2_ASAP7_75t_L g3481 ( 
.A(n_2950),
.B(n_1851),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_2950),
.Y(n_3482)
);

O2A1O1Ixp33_ASAP7_75t_L g3483 ( 
.A1(n_2827),
.A2(n_1862),
.B(n_1865),
.C(n_1863),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_2912),
.B(n_1678),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_2912),
.B(n_1682),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_2912),
.Y(n_3486)
);

AOI21xp5_ASAP7_75t_L g3487 ( 
.A1(n_2744),
.A2(n_1699),
.B(n_1687),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_2623),
.B(n_1699),
.Y(n_3488)
);

NOR2x1p5_ASAP7_75t_L g3489 ( 
.A(n_2835),
.B(n_1701),
.Y(n_3489)
);

NOR2xp33_ASAP7_75t_L g3490 ( 
.A(n_2705),
.B(n_1701),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_SL g3491 ( 
.A(n_3018),
.B(n_1765),
.Y(n_3491)
);

NOR2x1p5_ASAP7_75t_L g3492 ( 
.A(n_2835),
.B(n_1719),
.Y(n_3492)
);

OR2x2_ASAP7_75t_L g3493 ( 
.A(n_2708),
.B(n_1765),
.Y(n_3493)
);

CKINVDCx20_ASAP7_75t_R g3494 ( 
.A(n_2653),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_2618),
.Y(n_3495)
);

A2O1A1Ixp33_ASAP7_75t_L g3496 ( 
.A1(n_2987),
.A2(n_1719),
.B(n_1819),
.C(n_1732),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_2623),
.B(n_2),
.Y(n_3497)
);

NOR2xp33_ASAP7_75t_R g3498 ( 
.A(n_2653),
.B(n_2),
.Y(n_3498)
);

BUFx6f_ASAP7_75t_L g3499 ( 
.A(n_2753),
.Y(n_3499)
);

NOR2xp33_ASAP7_75t_L g3500 ( 
.A(n_2705),
.B(n_240),
.Y(n_3500)
);

NOR2xp33_ASAP7_75t_L g3501 ( 
.A(n_2705),
.B(n_240),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_2618),
.Y(n_3502)
);

NOR2xp33_ASAP7_75t_L g3503 ( 
.A(n_2705),
.B(n_240),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_2623),
.B(n_2),
.Y(n_3504)
);

AOI22xp33_ASAP7_75t_SL g3505 ( 
.A1(n_2807),
.A2(n_1819),
.B1(n_1831),
.B2(n_1732),
.Y(n_3505)
);

BUFx6f_ASAP7_75t_L g3506 ( 
.A(n_2753),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_SL g3507 ( 
.A(n_3018),
.B(n_1732),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_2618),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_2623),
.B(n_3),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_2618),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_2623),
.B(n_3),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_2618),
.Y(n_3512)
);

AND2x2_ASAP7_75t_L g3513 ( 
.A(n_2623),
.B(n_241),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_2623),
.B(n_3),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_SL g3515 ( 
.A(n_3018),
.B(n_1819),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_L g3516 ( 
.A(n_2623),
.B(n_4),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_2710),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_L g3518 ( 
.A(n_2623),
.B(n_4),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_2623),
.B(n_4),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_2623),
.B(n_4),
.Y(n_3520)
);

INVx2_ASAP7_75t_L g3521 ( 
.A(n_2710),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_2623),
.B(n_5),
.Y(n_3522)
);

INVx3_ASAP7_75t_L g3523 ( 
.A(n_2634),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_2618),
.Y(n_3524)
);

NOR3x1_ASAP7_75t_L g3525 ( 
.A(n_2627),
.B(n_242),
.C(n_241),
.Y(n_3525)
);

NAND2xp33_ASAP7_75t_L g3526 ( 
.A(n_2707),
.B(n_1819),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_2623),
.B(n_5),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_2623),
.B(n_5),
.Y(n_3528)
);

AOI22xp5_ASAP7_75t_L g3529 ( 
.A1(n_2987),
.A2(n_1848),
.B1(n_1831),
.B2(n_242),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_2710),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_2623),
.B(n_6),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_2623),
.B(n_6),
.Y(n_3532)
);

NOR2xp67_ASAP7_75t_L g3533 ( 
.A(n_2971),
.B(n_242),
.Y(n_3533)
);

AOI22xp5_ASAP7_75t_L g3534 ( 
.A1(n_2987),
.A2(n_1848),
.B1(n_1831),
.B2(n_243),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_L g3535 ( 
.A(n_2623),
.B(n_6),
.Y(n_3535)
);

INVx2_ASAP7_75t_L g3536 ( 
.A(n_2710),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_2623),
.B(n_6),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_2618),
.Y(n_3538)
);

INVx2_ASAP7_75t_SL g3539 ( 
.A(n_2971),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_2710),
.Y(n_3540)
);

INVx5_ASAP7_75t_L g3541 ( 
.A(n_2988),
.Y(n_3541)
);

AOI22xp5_ASAP7_75t_L g3542 ( 
.A1(n_2987),
.A2(n_1848),
.B1(n_1831),
.B2(n_243),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_2618),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_SL g3544 ( 
.A(n_3018),
.B(n_1848),
.Y(n_3544)
);

OR2x6_ASAP7_75t_L g3545 ( 
.A(n_2907),
.B(n_241),
.Y(n_3545)
);

INVx2_ASAP7_75t_L g3546 ( 
.A(n_2710),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_2623),
.B(n_7),
.Y(n_3547)
);

A2O1A1Ixp33_ASAP7_75t_L g3548 ( 
.A1(n_2987),
.A2(n_244),
.B(n_245),
.C(n_243),
.Y(n_3548)
);

INVx2_ASAP7_75t_L g3549 ( 
.A(n_2710),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_SL g3550 ( 
.A(n_3018),
.B(n_244),
.Y(n_3550)
);

O2A1O1Ixp33_ASAP7_75t_L g3551 ( 
.A1(n_2987),
.A2(n_246),
.B(n_247),
.C(n_244),
.Y(n_3551)
);

NOR2xp33_ASAP7_75t_L g3552 ( 
.A(n_2705),
.B(n_246),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_2623),
.B(n_7),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_2623),
.B(n_7),
.Y(n_3554)
);

INVx2_ASAP7_75t_L g3555 ( 
.A(n_2710),
.Y(n_3555)
);

INVx3_ASAP7_75t_L g3556 ( 
.A(n_2634),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_SL g3557 ( 
.A(n_3018),
.B(n_247),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_SL g3558 ( 
.A(n_3018),
.B(n_247),
.Y(n_3558)
);

NOR2xp33_ASAP7_75t_L g3559 ( 
.A(n_2705),
.B(n_248),
.Y(n_3559)
);

INVx2_ASAP7_75t_L g3560 ( 
.A(n_2710),
.Y(n_3560)
);

NOR2xp33_ASAP7_75t_L g3561 ( 
.A(n_2705),
.B(n_248),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_2623),
.B(n_7),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_2618),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_2623),
.B(n_8),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_2618),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_2623),
.B(n_8),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_2623),
.B(n_8),
.Y(n_3567)
);

BUFx3_ASAP7_75t_L g3568 ( 
.A(n_2988),
.Y(n_3568)
);

INVx2_ASAP7_75t_SL g3569 ( 
.A(n_2971),
.Y(n_3569)
);

AOI22xp5_ASAP7_75t_L g3570 ( 
.A1(n_2987),
.A2(n_249),
.B1(n_250),
.B2(n_248),
.Y(n_3570)
);

NOR2xp33_ASAP7_75t_L g3571 ( 
.A(n_2705),
.B(n_249),
.Y(n_3571)
);

A2O1A1Ixp33_ASAP7_75t_L g3572 ( 
.A1(n_2987),
.A2(n_251),
.B(n_252),
.C(n_250),
.Y(n_3572)
);

OAI221xp5_ASAP7_75t_L g3573 ( 
.A1(n_2725),
.A2(n_252),
.B1(n_253),
.B2(n_251),
.C(n_250),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_2618),
.Y(n_3574)
);

NOR2xp67_ASAP7_75t_L g3575 ( 
.A(n_2971),
.B(n_256),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_2623),
.B(n_9),
.Y(n_3576)
);

AND2x2_ASAP7_75t_L g3577 ( 
.A(n_2623),
.B(n_1154),
.Y(n_3577)
);

AND2x2_ASAP7_75t_L g3578 ( 
.A(n_2623),
.B(n_1154),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_2623),
.B(n_9),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_SL g3580 ( 
.A(n_3018),
.B(n_251),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_2618),
.Y(n_3581)
);

INVx2_ASAP7_75t_L g3582 ( 
.A(n_2710),
.Y(n_3582)
);

INVx4_ASAP7_75t_L g3583 ( 
.A(n_2971),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_SL g3584 ( 
.A(n_3018),
.B(n_252),
.Y(n_3584)
);

AND2x2_ASAP7_75t_L g3585 ( 
.A(n_2623),
.B(n_1158),
.Y(n_3585)
);

AOI22xp5_ASAP7_75t_L g3586 ( 
.A1(n_2987),
.A2(n_255),
.B1(n_256),
.B2(n_254),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_SL g3587 ( 
.A(n_3018),
.B(n_254),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_2618),
.Y(n_3588)
);

OAI22xp5_ASAP7_75t_L g3589 ( 
.A1(n_2741),
.A2(n_255),
.B1(n_256),
.B2(n_254),
.Y(n_3589)
);

INVx3_ASAP7_75t_L g3590 ( 
.A(n_2634),
.Y(n_3590)
);

NAND2xp5_ASAP7_75t_SL g3591 ( 
.A(n_3018),
.B(n_257),
.Y(n_3591)
);

OAI22xp5_ASAP7_75t_L g3592 ( 
.A1(n_2741),
.A2(n_258),
.B1(n_259),
.B2(n_257),
.Y(n_3592)
);

CKINVDCx5p33_ASAP7_75t_R g3593 ( 
.A(n_2653),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_2623),
.B(n_10),
.Y(n_3594)
);

NOR2xp33_ASAP7_75t_L g3595 ( 
.A(n_2705),
.B(n_258),
.Y(n_3595)
);

AOI21xp5_ASAP7_75t_L g3596 ( 
.A1(n_2744),
.A2(n_10),
.B(n_11),
.Y(n_3596)
);

INVx2_ASAP7_75t_L g3597 ( 
.A(n_2710),
.Y(n_3597)
);

AND2x2_ASAP7_75t_L g3598 ( 
.A(n_2623),
.B(n_1163),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_2623),
.B(n_11),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_2623),
.B(n_11),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_2623),
.B(n_11),
.Y(n_3601)
);

INVx8_ASAP7_75t_L g3602 ( 
.A(n_2971),
.Y(n_3602)
);

INVx2_ASAP7_75t_L g3603 ( 
.A(n_2710),
.Y(n_3603)
);

NOR2xp33_ASAP7_75t_L g3604 ( 
.A(n_2705),
.B(n_258),
.Y(n_3604)
);

INVx8_ASAP7_75t_L g3605 ( 
.A(n_2971),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_2618),
.Y(n_3606)
);

HB1xp67_ASAP7_75t_L g3607 ( 
.A(n_3009),
.Y(n_3607)
);

BUFx8_ASAP7_75t_L g3608 ( 
.A(n_2988),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_SL g3609 ( 
.A(n_3018),
.B(n_259),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_2623),
.B(n_12),
.Y(n_3610)
);

INVx2_ASAP7_75t_L g3611 ( 
.A(n_2710),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_L g3612 ( 
.A(n_2623),
.B(n_12),
.Y(n_3612)
);

NOR2xp33_ASAP7_75t_L g3613 ( 
.A(n_2705),
.B(n_259),
.Y(n_3613)
);

INVx2_ASAP7_75t_L g3614 ( 
.A(n_2710),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_2618),
.Y(n_3615)
);

OAI22xp5_ASAP7_75t_L g3616 ( 
.A1(n_2741),
.A2(n_261),
.B1(n_262),
.B2(n_260),
.Y(n_3616)
);

INVx2_ASAP7_75t_SL g3617 ( 
.A(n_2971),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_L g3618 ( 
.A(n_2623),
.B(n_12),
.Y(n_3618)
);

INVx4_ASAP7_75t_L g3619 ( 
.A(n_2971),
.Y(n_3619)
);

NOR2xp33_ASAP7_75t_L g3620 ( 
.A(n_2705),
.B(n_260),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_2623),
.B(n_13),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_2623),
.B(n_13),
.Y(n_3622)
);

NOR2xp33_ASAP7_75t_L g3623 ( 
.A(n_2705),
.B(n_260),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_SL g3624 ( 
.A(n_3018),
.B(n_261),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_2623),
.B(n_14),
.Y(n_3625)
);

AO22x1_ASAP7_75t_L g3626 ( 
.A1(n_2983),
.A2(n_263),
.B1(n_264),
.B2(n_261),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_SL g3627 ( 
.A(n_3018),
.B(n_262),
.Y(n_3627)
);

O2A1O1Ixp33_ASAP7_75t_L g3628 ( 
.A1(n_2987),
.A2(n_263),
.B(n_264),
.C(n_262),
.Y(n_3628)
);

AND2x6_ASAP7_75t_SL g3629 ( 
.A(n_2629),
.B(n_263),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_SL g3630 ( 
.A(n_3018),
.B(n_264),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_2618),
.Y(n_3631)
);

OAI221xp5_ASAP7_75t_L g3632 ( 
.A1(n_2725),
.A2(n_267),
.B1(n_268),
.B2(n_266),
.C(n_265),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_2618),
.Y(n_3633)
);

NOR2xp33_ASAP7_75t_L g3634 ( 
.A(n_2705),
.B(n_265),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_SL g3635 ( 
.A(n_3018),
.B(n_265),
.Y(n_3635)
);

OR2x2_ASAP7_75t_L g3636 ( 
.A(n_2708),
.B(n_266),
.Y(n_3636)
);

BUFx5_ASAP7_75t_L g3637 ( 
.A(n_2980),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_2623),
.B(n_14),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_2618),
.Y(n_3639)
);

AND2x2_ASAP7_75t_L g3640 ( 
.A(n_2623),
.B(n_1158),
.Y(n_3640)
);

NOR2xp33_ASAP7_75t_L g3641 ( 
.A(n_2705),
.B(n_266),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_2623),
.B(n_14),
.Y(n_3642)
);

AOI22xp5_ASAP7_75t_L g3643 ( 
.A1(n_2987),
.A2(n_268),
.B1(n_269),
.B2(n_267),
.Y(n_3643)
);

O2A1O1Ixp5_ASAP7_75t_L g3644 ( 
.A1(n_2731),
.A2(n_269),
.B(n_270),
.C(n_267),
.Y(n_3644)
);

BUFx6f_ASAP7_75t_SL g3645 ( 
.A(n_2714),
.Y(n_3645)
);

HB1xp67_ASAP7_75t_L g3646 ( 
.A(n_3009),
.Y(n_3646)
);

AOI22xp5_ASAP7_75t_L g3647 ( 
.A1(n_2987),
.A2(n_271),
.B1(n_272),
.B2(n_270),
.Y(n_3647)
);

CKINVDCx14_ASAP7_75t_R g3648 ( 
.A(n_2653),
.Y(n_3648)
);

INVx2_ASAP7_75t_L g3649 ( 
.A(n_2710),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_L g3650 ( 
.A(n_2623),
.B(n_14),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_2710),
.Y(n_3651)
);

NOR2xp67_ASAP7_75t_L g3652 ( 
.A(n_2971),
.B(n_272),
.Y(n_3652)
);

INVx2_ASAP7_75t_L g3653 ( 
.A(n_2710),
.Y(n_3653)
);

INVx2_ASAP7_75t_L g3654 ( 
.A(n_2710),
.Y(n_3654)
);

AND2x2_ASAP7_75t_L g3655 ( 
.A(n_2623),
.B(n_1163),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_SL g3656 ( 
.A(n_3018),
.B(n_270),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_2623),
.B(n_15),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_2618),
.Y(n_3658)
);

INVx2_ASAP7_75t_L g3659 ( 
.A(n_2710),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_SL g3660 ( 
.A(n_3018),
.B(n_271),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_2623),
.B(n_15),
.Y(n_3661)
);

OR2x2_ASAP7_75t_L g3662 ( 
.A(n_2708),
.B(n_272),
.Y(n_3662)
);

NOR2xp33_ASAP7_75t_L g3663 ( 
.A(n_2705),
.B(n_273),
.Y(n_3663)
);

NOR2x1p5_ASAP7_75t_L g3664 ( 
.A(n_2835),
.B(n_273),
.Y(n_3664)
);

NOR2xp67_ASAP7_75t_L g3665 ( 
.A(n_2971),
.B(n_276),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_SL g3666 ( 
.A(n_3018),
.B(n_273),
.Y(n_3666)
);

OAI22xp33_ASAP7_75t_L g3667 ( 
.A1(n_2708),
.A2(n_275),
.B1(n_276),
.B2(n_274),
.Y(n_3667)
);

AOI22xp33_ASAP7_75t_L g3668 ( 
.A1(n_2695),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_2623),
.B(n_16),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_SL g3670 ( 
.A(n_3018),
.B(n_274),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_2618),
.Y(n_3671)
);

NOR3xp33_ASAP7_75t_L g3672 ( 
.A(n_2682),
.B(n_275),
.C(n_274),
.Y(n_3672)
);

INVxp67_ASAP7_75t_L g3673 ( 
.A(n_3009),
.Y(n_3673)
);

AOI22xp33_ASAP7_75t_L g3674 ( 
.A1(n_2695),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_3674)
);

NAND2xp33_ASAP7_75t_L g3675 ( 
.A(n_2707),
.B(n_16),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_SL g3676 ( 
.A(n_3018),
.B(n_275),
.Y(n_3676)
);

NOR2xp33_ASAP7_75t_L g3677 ( 
.A(n_2705),
.B(n_276),
.Y(n_3677)
);

AOI22xp5_ASAP7_75t_L g3678 ( 
.A1(n_2987),
.A2(n_278),
.B1(n_279),
.B2(n_277),
.Y(n_3678)
);

NOR2xp33_ASAP7_75t_L g3679 ( 
.A(n_2705),
.B(n_277),
.Y(n_3679)
);

INVx2_ASAP7_75t_L g3680 ( 
.A(n_2710),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_2623),
.B(n_17),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_2623),
.B(n_17),
.Y(n_3682)
);

INVx4_ASAP7_75t_L g3683 ( 
.A(n_2971),
.Y(n_3683)
);

NAND2xp33_ASAP7_75t_L g3684 ( 
.A(n_2707),
.B(n_18),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_SL g3685 ( 
.A(n_3018),
.B(n_277),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_SL g3686 ( 
.A(n_3018),
.B(n_278),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_2623),
.B(n_18),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_L g3688 ( 
.A(n_2623),
.B(n_19),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_2618),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_2618),
.Y(n_3690)
);

NAND2xp33_ASAP7_75t_L g3691 ( 
.A(n_2707),
.B(n_19),
.Y(n_3691)
);

AOI22xp5_ASAP7_75t_L g3692 ( 
.A1(n_2987),
.A2(n_280),
.B1(n_281),
.B2(n_278),
.Y(n_3692)
);

INVxp67_ASAP7_75t_L g3693 ( 
.A(n_3009),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_SL g3694 ( 
.A(n_3018),
.B(n_280),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_2623),
.B(n_19),
.Y(n_3695)
);

AOI22xp33_ASAP7_75t_SL g3696 ( 
.A1(n_2807),
.A2(n_281),
.B1(n_282),
.B2(n_280),
.Y(n_3696)
);

BUFx3_ASAP7_75t_L g3697 ( 
.A(n_2988),
.Y(n_3697)
);

NOR2xp33_ASAP7_75t_L g3698 ( 
.A(n_2705),
.B(n_281),
.Y(n_3698)
);

AOI22xp33_ASAP7_75t_L g3699 ( 
.A1(n_2695),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_3699)
);

NOR2xp67_ASAP7_75t_L g3700 ( 
.A(n_2971),
.B(n_289),
.Y(n_3700)
);

INVx2_ASAP7_75t_L g3701 ( 
.A(n_2710),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_2623),
.B(n_20),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_2623),
.B(n_20),
.Y(n_3703)
);

NOR2xp33_ASAP7_75t_L g3704 ( 
.A(n_2705),
.B(n_282),
.Y(n_3704)
);

OAI22xp5_ASAP7_75t_L g3705 ( 
.A1(n_2741),
.A2(n_283),
.B1(n_284),
.B2(n_282),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_SL g3706 ( 
.A(n_3018),
.B(n_284),
.Y(n_3706)
);

INVx2_ASAP7_75t_L g3707 ( 
.A(n_2710),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_2618),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_2623),
.B(n_20),
.Y(n_3709)
);

AND2x6_ASAP7_75t_SL g3710 ( 
.A(n_2629),
.B(n_285),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_3039),
.B(n_284),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3051),
.B(n_285),
.Y(n_3712)
);

A2O1A1Ixp33_ASAP7_75t_L g3713 ( 
.A1(n_3204),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_3713)
);

AOI21xp5_ASAP7_75t_L g3714 ( 
.A1(n_3526),
.A2(n_287),
.B(n_286),
.Y(n_3714)
);

OAI22xp5_ASAP7_75t_L g3715 ( 
.A1(n_3051),
.A2(n_287),
.B1(n_288),
.B2(n_286),
.Y(n_3715)
);

AND2x4_ASAP7_75t_SL g3716 ( 
.A(n_3583),
.B(n_286),
.Y(n_3716)
);

AND2x2_ASAP7_75t_L g3717 ( 
.A(n_3046),
.B(n_3049),
.Y(n_3717)
);

INVx2_ASAP7_75t_L g3718 ( 
.A(n_3085),
.Y(n_3718)
);

A2O1A1Ixp33_ASAP7_75t_L g3719 ( 
.A1(n_3190),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_3719)
);

AND2x4_ASAP7_75t_L g3720 ( 
.A(n_3541),
.B(n_287),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3101),
.Y(n_3721)
);

AOI21xp5_ASAP7_75t_L g3722 ( 
.A1(n_3337),
.A2(n_290),
.B(n_288),
.Y(n_3722)
);

BUFx6f_ASAP7_75t_L g3723 ( 
.A(n_3193),
.Y(n_3723)
);

NOR2xp33_ASAP7_75t_SL g3724 ( 
.A(n_3083),
.B(n_290),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_SL g3725 ( 
.A(n_3447),
.B(n_291),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_SL g3726 ( 
.A(n_3140),
.B(n_291),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_L g3727 ( 
.A(n_3513),
.B(n_292),
.Y(n_3727)
);

OAI21xp5_ASAP7_75t_L g3728 ( 
.A1(n_3420),
.A2(n_3237),
.B(n_3243),
.Y(n_3728)
);

INVx3_ASAP7_75t_L g3729 ( 
.A(n_3602),
.Y(n_3729)
);

AOI21xp5_ASAP7_75t_L g3730 ( 
.A1(n_3337),
.A2(n_293),
.B(n_292),
.Y(n_3730)
);

INVx2_ASAP7_75t_L g3731 ( 
.A(n_3110),
.Y(n_3731)
);

INVx2_ASAP7_75t_L g3732 ( 
.A(n_3123),
.Y(n_3732)
);

INVx3_ASAP7_75t_L g3733 ( 
.A(n_3602),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_L g3734 ( 
.A(n_3577),
.B(n_292),
.Y(n_3734)
);

AND2x2_ASAP7_75t_L g3735 ( 
.A(n_3180),
.B(n_293),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3090),
.Y(n_3736)
);

INVx2_ASAP7_75t_L g3737 ( 
.A(n_3136),
.Y(n_3737)
);

AOI21xp5_ASAP7_75t_L g3738 ( 
.A1(n_3066),
.A2(n_295),
.B(n_294),
.Y(n_3738)
);

INVx3_ASAP7_75t_L g3739 ( 
.A(n_3602),
.Y(n_3739)
);

AND2x6_ASAP7_75t_L g3740 ( 
.A(n_3438),
.B(n_294),
.Y(n_3740)
);

AOI21xp5_ASAP7_75t_L g3741 ( 
.A1(n_3120),
.A2(n_295),
.B(n_294),
.Y(n_3741)
);

NOR2xp33_ASAP7_75t_L g3742 ( 
.A(n_3043),
.B(n_296),
.Y(n_3742)
);

AOI21xp5_ASAP7_75t_L g3743 ( 
.A1(n_3487),
.A2(n_297),
.B(n_296),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3578),
.B(n_296),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3245),
.Y(n_3745)
);

INVxp67_ASAP7_75t_L g3746 ( 
.A(n_3075),
.Y(n_3746)
);

AOI21xp5_ASAP7_75t_L g3747 ( 
.A1(n_3233),
.A2(n_299),
.B(n_298),
.Y(n_3747)
);

INVxp67_ASAP7_75t_L g3748 ( 
.A(n_3075),
.Y(n_3748)
);

AOI21xp5_ASAP7_75t_L g3749 ( 
.A1(n_3675),
.A2(n_299),
.B(n_298),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3056),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3072),
.Y(n_3751)
);

BUFx6f_ASAP7_75t_L g3752 ( 
.A(n_3193),
.Y(n_3752)
);

NOR2xp33_ASAP7_75t_L g3753 ( 
.A(n_3290),
.B(n_298),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_L g3754 ( 
.A(n_3585),
.B(n_300),
.Y(n_3754)
);

BUFx2_ASAP7_75t_L g3755 ( 
.A(n_3494),
.Y(n_3755)
);

NOR2xp33_ASAP7_75t_L g3756 ( 
.A(n_3328),
.B(n_300),
.Y(n_3756)
);

NAND2xp5_ASAP7_75t_L g3757 ( 
.A(n_3598),
.B(n_300),
.Y(n_3757)
);

AOI21xp5_ASAP7_75t_L g3758 ( 
.A1(n_3684),
.A2(n_302),
.B(n_301),
.Y(n_3758)
);

AOI21xp5_ASAP7_75t_L g3759 ( 
.A1(n_3691),
.A2(n_302),
.B(n_301),
.Y(n_3759)
);

OAI21xp5_ASAP7_75t_L g3760 ( 
.A1(n_3122),
.A2(n_3126),
.B(n_3096),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_SL g3761 ( 
.A(n_3140),
.B(n_3117),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_L g3762 ( 
.A(n_3640),
.B(n_301),
.Y(n_3762)
);

AOI21xp5_ASAP7_75t_L g3763 ( 
.A1(n_3234),
.A2(n_303),
.B(n_302),
.Y(n_3763)
);

AOI21xp5_ASAP7_75t_L g3764 ( 
.A1(n_3234),
.A2(n_304),
.B(n_303),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_L g3765 ( 
.A(n_3655),
.B(n_303),
.Y(n_3765)
);

BUFx3_ASAP7_75t_L g3766 ( 
.A(n_3608),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_SL g3767 ( 
.A(n_3117),
.B(n_3124),
.Y(n_3767)
);

BUFx8_ASAP7_75t_L g3768 ( 
.A(n_3645),
.Y(n_3768)
);

A2O1A1Ixp33_ASAP7_75t_L g3769 ( 
.A1(n_3077),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_3769)
);

AOI21xp5_ASAP7_75t_L g3770 ( 
.A1(n_3220),
.A2(n_3322),
.B(n_3071),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3084),
.Y(n_3771)
);

AOI21xp5_ASAP7_75t_L g3772 ( 
.A1(n_3320),
.A2(n_305),
.B(n_304),
.Y(n_3772)
);

NOR2xp33_ASAP7_75t_L g3773 ( 
.A(n_3277),
.B(n_305),
.Y(n_3773)
);

AOI21xp5_ASAP7_75t_L g3774 ( 
.A1(n_3446),
.A2(n_307),
.B(n_306),
.Y(n_3774)
);

A2O1A1Ixp33_ASAP7_75t_L g3775 ( 
.A1(n_3077),
.A2(n_24),
.B(n_22),
.C(n_23),
.Y(n_3775)
);

O2A1O1Ixp33_ASAP7_75t_L g3776 ( 
.A1(n_3471),
.A2(n_307),
.B(n_308),
.C(n_306),
.Y(n_3776)
);

OAI21xp33_ASAP7_75t_L g3777 ( 
.A1(n_3490),
.A2(n_24),
.B(n_25),
.Y(n_3777)
);

AOI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_3455),
.A2(n_3250),
.B(n_3417),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_3192),
.B(n_306),
.Y(n_3779)
);

AOI21xp5_ASAP7_75t_L g3780 ( 
.A1(n_3417),
.A2(n_309),
.B(n_308),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3143),
.Y(n_3781)
);

OAI22xp5_ASAP7_75t_L g3782 ( 
.A1(n_3108),
.A2(n_310),
.B1(n_311),
.B2(n_309),
.Y(n_3782)
);

O2A1O1Ixp33_ASAP7_75t_L g3783 ( 
.A1(n_3415),
.A2(n_311),
.B(n_312),
.C(n_310),
.Y(n_3783)
);

BUFx2_ASAP7_75t_SL g3784 ( 
.A(n_3645),
.Y(n_3784)
);

NOR2xp33_ASAP7_75t_L g3785 ( 
.A(n_3280),
.B(n_310),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_3093),
.B(n_311),
.Y(n_3786)
);

INVx2_ASAP7_75t_L g3787 ( 
.A(n_3154),
.Y(n_3787)
);

OAI22xp5_ASAP7_75t_L g3788 ( 
.A1(n_3545),
.A2(n_313),
.B1(n_314),
.B2(n_312),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_SL g3789 ( 
.A(n_3124),
.B(n_313),
.Y(n_3789)
);

BUFx6f_ASAP7_75t_L g3790 ( 
.A(n_3193),
.Y(n_3790)
);

OAI21xp5_ASAP7_75t_L g3791 ( 
.A1(n_3095),
.A2(n_24),
.B(n_25),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3116),
.B(n_313),
.Y(n_3792)
);

OAI21xp5_ASAP7_75t_L g3793 ( 
.A1(n_3099),
.A2(n_24),
.B(n_25),
.Y(n_3793)
);

INVx4_ASAP7_75t_L g3794 ( 
.A(n_3605),
.Y(n_3794)
);

OAI21xp5_ASAP7_75t_L g3795 ( 
.A1(n_3100),
.A2(n_26),
.B(n_27),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3495),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_SL g3797 ( 
.A(n_3541),
.B(n_3251),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3502),
.Y(n_3798)
);

BUFx6f_ASAP7_75t_L g3799 ( 
.A(n_3499),
.Y(n_3799)
);

AOI21xp5_ASAP7_75t_L g3800 ( 
.A1(n_3707),
.A2(n_316),
.B(n_315),
.Y(n_3800)
);

NAND2x1p5_ASAP7_75t_L g3801 ( 
.A(n_3541),
.B(n_316),
.Y(n_3801)
);

INVx1_ASAP7_75t_SL g3802 ( 
.A(n_3058),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_L g3803 ( 
.A(n_3191),
.B(n_316),
.Y(n_3803)
);

INVx2_ASAP7_75t_L g3804 ( 
.A(n_3156),
.Y(n_3804)
);

AOI21xp5_ASAP7_75t_L g3805 ( 
.A1(n_3054),
.A2(n_319),
.B(n_318),
.Y(n_3805)
);

BUFx8_ASAP7_75t_L g3806 ( 
.A(n_3456),
.Y(n_3806)
);

OR2x2_ASAP7_75t_L g3807 ( 
.A(n_3150),
.B(n_318),
.Y(n_3807)
);

AOI22xp33_ASAP7_75t_L g3808 ( 
.A1(n_3451),
.A2(n_320),
.B1(n_321),
.B2(n_319),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_L g3809 ( 
.A(n_3360),
.B(n_319),
.Y(n_3809)
);

NAND2xp33_ASAP7_75t_L g3810 ( 
.A(n_3097),
.B(n_320),
.Y(n_3810)
);

AND2x2_ASAP7_75t_L g3811 ( 
.A(n_3098),
.B(n_321),
.Y(n_3811)
);

AOI21xp5_ASAP7_75t_L g3812 ( 
.A1(n_3701),
.A2(n_322),
.B(n_321),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3508),
.Y(n_3813)
);

NOR2x1_ASAP7_75t_R g3814 ( 
.A(n_3593),
.B(n_322),
.Y(n_3814)
);

NOR2xp33_ASAP7_75t_L g3815 ( 
.A(n_3076),
.B(n_322),
.Y(n_3815)
);

AOI21xp5_ASAP7_75t_L g3816 ( 
.A1(n_3055),
.A2(n_324),
.B(n_323),
.Y(n_3816)
);

NOR3xp33_ASAP7_75t_L g3817 ( 
.A(n_3449),
.B(n_325),
.C(n_324),
.Y(n_3817)
);

OAI22xp5_ASAP7_75t_L g3818 ( 
.A1(n_3545),
.A2(n_326),
.B1(n_327),
.B2(n_325),
.Y(n_3818)
);

AOI21xp33_ASAP7_75t_L g3819 ( 
.A1(n_3213),
.A2(n_327),
.B(n_326),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3510),
.B(n_327),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_3512),
.B(n_328),
.Y(n_3821)
);

OAI22xp5_ASAP7_75t_L g3822 ( 
.A1(n_3545),
.A2(n_329),
.B1(n_330),
.B2(n_328),
.Y(n_3822)
);

AOI21xp5_ASAP7_75t_L g3823 ( 
.A1(n_3061),
.A2(n_330),
.B(n_329),
.Y(n_3823)
);

NOR2xp33_ASAP7_75t_L g3824 ( 
.A(n_3278),
.B(n_329),
.Y(n_3824)
);

NOR2xp33_ASAP7_75t_L g3825 ( 
.A(n_3223),
.B(n_330),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_L g3826 ( 
.A(n_3524),
.B(n_331),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_L g3827 ( 
.A(n_3538),
.B(n_3543),
.Y(n_3827)
);

NAND2xp5_ASAP7_75t_L g3828 ( 
.A(n_3563),
.B(n_331),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_SL g3829 ( 
.A(n_3251),
.B(n_332),
.Y(n_3829)
);

AOI21xp5_ASAP7_75t_L g3830 ( 
.A1(n_3063),
.A2(n_3521),
.B(n_3517),
.Y(n_3830)
);

INVx2_ASAP7_75t_L g3831 ( 
.A(n_3161),
.Y(n_3831)
);

OAI21xp5_ASAP7_75t_L g3832 ( 
.A1(n_3102),
.A2(n_26),
.B(n_27),
.Y(n_3832)
);

AND2x2_ASAP7_75t_L g3833 ( 
.A(n_3080),
.B(n_332),
.Y(n_3833)
);

NOR2xp33_ASAP7_75t_SL g3834 ( 
.A(n_3088),
.B(n_333),
.Y(n_3834)
);

AOI21xp5_ASAP7_75t_L g3835 ( 
.A1(n_3530),
.A2(n_334),
.B(n_333),
.Y(n_3835)
);

AO21x1_ASAP7_75t_L g3836 ( 
.A1(n_3596),
.A2(n_334),
.B(n_333),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3565),
.B(n_334),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_3574),
.B(n_335),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3581),
.Y(n_3839)
);

AO21x1_ASAP7_75t_L g3840 ( 
.A1(n_3551),
.A2(n_336),
.B(n_335),
.Y(n_3840)
);

AOI21xp5_ASAP7_75t_L g3841 ( 
.A1(n_3536),
.A2(n_336),
.B(n_335),
.Y(n_3841)
);

NOR2xp33_ASAP7_75t_L g3842 ( 
.A(n_3221),
.B(n_336),
.Y(n_3842)
);

HB1xp67_ASAP7_75t_L g3843 ( 
.A(n_3607),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_L g3844 ( 
.A(n_3588),
.B(n_337),
.Y(n_3844)
);

BUFx3_ASAP7_75t_L g3845 ( 
.A(n_3608),
.Y(n_3845)
);

AOI21xp5_ASAP7_75t_L g3846 ( 
.A1(n_3540),
.A2(n_338),
.B(n_337),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_3606),
.B(n_338),
.Y(n_3847)
);

AOI21xp5_ASAP7_75t_L g3848 ( 
.A1(n_3546),
.A2(n_340),
.B(n_339),
.Y(n_3848)
);

AOI21xp5_ASAP7_75t_L g3849 ( 
.A1(n_3549),
.A2(n_3560),
.B(n_3555),
.Y(n_3849)
);

NAND2x1p5_ASAP7_75t_L g3850 ( 
.A(n_3583),
.B(n_339),
.Y(n_3850)
);

O2A1O1Ixp33_ASAP7_75t_L g3851 ( 
.A1(n_3399),
.A2(n_340),
.B(n_341),
.C(n_339),
.Y(n_3851)
);

AND2x2_ASAP7_75t_L g3852 ( 
.A(n_3252),
.B(n_3171),
.Y(n_3852)
);

BUFx6f_ASAP7_75t_L g3853 ( 
.A(n_3499),
.Y(n_3853)
);

NOR2xp33_ASAP7_75t_L g3854 ( 
.A(n_3222),
.B(n_3383),
.Y(n_3854)
);

NOR2xp67_ASAP7_75t_L g3855 ( 
.A(n_3619),
.B(n_340),
.Y(n_3855)
);

INVx2_ASAP7_75t_L g3856 ( 
.A(n_3177),
.Y(n_3856)
);

AO21x1_ASAP7_75t_L g3857 ( 
.A1(n_3628),
.A2(n_342),
.B(n_341),
.Y(n_3857)
);

BUFx12f_ASAP7_75t_L g3858 ( 
.A(n_3210),
.Y(n_3858)
);

AND2x2_ASAP7_75t_L g3859 ( 
.A(n_3044),
.B(n_342),
.Y(n_3859)
);

OAI21xp33_ASAP7_75t_SL g3860 ( 
.A1(n_3570),
.A2(n_343),
.B(n_342),
.Y(n_3860)
);

BUFx6f_ASAP7_75t_L g3861 ( 
.A(n_3499),
.Y(n_3861)
);

A2O1A1Ixp33_ASAP7_75t_L g3862 ( 
.A1(n_3496),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_3862)
);

AOI21xp5_ASAP7_75t_L g3863 ( 
.A1(n_3582),
.A2(n_344),
.B(n_343),
.Y(n_3863)
);

AOI21x1_ASAP7_75t_L g3864 ( 
.A1(n_3368),
.A2(n_344),
.B(n_343),
.Y(n_3864)
);

INVxp67_ASAP7_75t_L g3865 ( 
.A(n_3646),
.Y(n_3865)
);

AOI21xp5_ASAP7_75t_L g3866 ( 
.A1(n_3597),
.A2(n_345),
.B(n_344),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_L g3867 ( 
.A(n_3615),
.B(n_346),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3631),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_SL g3869 ( 
.A(n_3187),
.B(n_346),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_3633),
.B(n_347),
.Y(n_3870)
);

AOI21xp5_ASAP7_75t_L g3871 ( 
.A1(n_3603),
.A2(n_348),
.B(n_347),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_SL g3872 ( 
.A(n_3125),
.B(n_348),
.Y(n_3872)
);

AOI21x1_ASAP7_75t_L g3873 ( 
.A1(n_3412),
.A2(n_350),
.B(n_349),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_SL g3874 ( 
.A(n_3125),
.B(n_349),
.Y(n_3874)
);

INVx2_ASAP7_75t_L g3875 ( 
.A(n_3188),
.Y(n_3875)
);

BUFx6f_ASAP7_75t_L g3876 ( 
.A(n_3506),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_3639),
.B(n_349),
.Y(n_3877)
);

OR2x2_ASAP7_75t_L g3878 ( 
.A(n_3209),
.B(n_350),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_L g3879 ( 
.A(n_3658),
.B(n_350),
.Y(n_3879)
);

OAI21xp5_ASAP7_75t_L g3880 ( 
.A1(n_3106),
.A2(n_27),
.B(n_28),
.Y(n_3880)
);

NOR2x1p5_ASAP7_75t_SL g3881 ( 
.A(n_3097),
.B(n_351),
.Y(n_3881)
);

AOI21xp5_ASAP7_75t_L g3882 ( 
.A1(n_3611),
.A2(n_352),
.B(n_351),
.Y(n_3882)
);

INVx3_ASAP7_75t_L g3883 ( 
.A(n_3605),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_L g3884 ( 
.A(n_3671),
.B(n_351),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_3689),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_L g3886 ( 
.A(n_3690),
.B(n_352),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_SL g3887 ( 
.A(n_3125),
.B(n_352),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_3708),
.B(n_353),
.Y(n_3888)
);

AOI21xp5_ASAP7_75t_L g3889 ( 
.A1(n_3614),
.A2(n_354),
.B(n_353),
.Y(n_3889)
);

AOI22xp5_ASAP7_75t_L g3890 ( 
.A1(n_3067),
.A2(n_355),
.B1(n_356),
.B2(n_354),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_SL g3891 ( 
.A(n_3129),
.B(n_354),
.Y(n_3891)
);

AOI22xp5_ASAP7_75t_L g3892 ( 
.A1(n_3045),
.A2(n_356),
.B1(n_357),
.B2(n_355),
.Y(n_3892)
);

AOI21xp5_ASAP7_75t_L g3893 ( 
.A1(n_3649),
.A2(n_356),
.B(n_355),
.Y(n_3893)
);

NAND2xp5_ASAP7_75t_L g3894 ( 
.A(n_3488),
.B(n_3497),
.Y(n_3894)
);

NOR2xp33_ASAP7_75t_SL g3895 ( 
.A(n_3088),
.B(n_357),
.Y(n_3895)
);

O2A1O1Ixp5_ASAP7_75t_L g3896 ( 
.A1(n_3232),
.A2(n_358),
.B(n_359),
.C(n_357),
.Y(n_3896)
);

O2A1O1Ixp33_ASAP7_75t_L g3897 ( 
.A1(n_3452),
.A2(n_360),
.B(n_361),
.C(n_358),
.Y(n_3897)
);

INVx4_ASAP7_75t_L g3898 ( 
.A(n_3605),
.Y(n_3898)
);

OAI21xp5_ASAP7_75t_L g3899 ( 
.A1(n_3109),
.A2(n_28),
.B(n_29),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_SL g3900 ( 
.A(n_3129),
.B(n_358),
.Y(n_3900)
);

NOR2xp33_ASAP7_75t_L g3901 ( 
.A(n_3212),
.B(n_360),
.Y(n_3901)
);

INVx3_ASAP7_75t_L g3902 ( 
.A(n_3370),
.Y(n_3902)
);

A2O1A1Ixp33_ASAP7_75t_L g3903 ( 
.A1(n_3405),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_3903)
);

NOR2xp33_ASAP7_75t_L g3904 ( 
.A(n_3037),
.B(n_360),
.Y(n_3904)
);

AOI22xp5_ASAP7_75t_L g3905 ( 
.A1(n_3034),
.A2(n_362),
.B1(n_363),
.B2(n_361),
.Y(n_3905)
);

INVxp67_ASAP7_75t_L g3906 ( 
.A(n_3144),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_SL g3907 ( 
.A(n_3129),
.B(n_361),
.Y(n_3907)
);

INVx3_ASAP7_75t_L g3908 ( 
.A(n_3370),
.Y(n_3908)
);

AOI21xp5_ASAP7_75t_L g3909 ( 
.A1(n_3651),
.A2(n_364),
.B(n_363),
.Y(n_3909)
);

NOR2xp33_ASAP7_75t_L g3910 ( 
.A(n_3157),
.B(n_363),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_3504),
.B(n_364),
.Y(n_3911)
);

AND2x4_ASAP7_75t_L g3912 ( 
.A(n_3073),
.B(n_3568),
.Y(n_3912)
);

AND2x4_ASAP7_75t_L g3913 ( 
.A(n_3697),
.B(n_365),
.Y(n_3913)
);

INVx2_ASAP7_75t_L g3914 ( 
.A(n_3199),
.Y(n_3914)
);

OAI22xp5_ASAP7_75t_L g3915 ( 
.A1(n_3044),
.A2(n_3529),
.B1(n_3542),
.B2(n_3534),
.Y(n_3915)
);

AOI21xp5_ASAP7_75t_L g3916 ( 
.A1(n_3653),
.A2(n_366),
.B(n_365),
.Y(n_3916)
);

NOR2xp33_ASAP7_75t_L g3917 ( 
.A(n_3283),
.B(n_365),
.Y(n_3917)
);

CKINVDCx10_ASAP7_75t_R g3918 ( 
.A(n_3456),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_SL g3919 ( 
.A(n_3241),
.B(n_366),
.Y(n_3919)
);

AOI21xp5_ASAP7_75t_L g3920 ( 
.A1(n_3654),
.A2(n_367),
.B(n_366),
.Y(n_3920)
);

AO21x1_ASAP7_75t_L g3921 ( 
.A1(n_3589),
.A2(n_368),
.B(n_367),
.Y(n_3921)
);

INVx3_ASAP7_75t_L g3922 ( 
.A(n_3370),
.Y(n_3922)
);

AOI21xp5_ASAP7_75t_L g3923 ( 
.A1(n_3659),
.A2(n_368),
.B(n_367),
.Y(n_3923)
);

AND2x4_ASAP7_75t_L g3924 ( 
.A(n_3152),
.B(n_368),
.Y(n_3924)
);

INVx3_ASAP7_75t_L g3925 ( 
.A(n_3423),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_SL g3926 ( 
.A(n_3241),
.B(n_369),
.Y(n_3926)
);

BUFx8_ASAP7_75t_L g3927 ( 
.A(n_3430),
.Y(n_3927)
);

AOI21xp5_ASAP7_75t_L g3928 ( 
.A1(n_3680),
.A2(n_370),
.B(n_369),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_3509),
.B(n_369),
.Y(n_3929)
);

NAND2xp33_ASAP7_75t_L g3930 ( 
.A(n_3097),
.B(n_370),
.Y(n_3930)
);

NOR2xp33_ASAP7_75t_L g3931 ( 
.A(n_3258),
.B(n_370),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_SL g3932 ( 
.A(n_3371),
.B(n_371),
.Y(n_3932)
);

BUFx2_ASAP7_75t_L g3933 ( 
.A(n_3152),
.Y(n_3933)
);

NOR2xp33_ASAP7_75t_L g3934 ( 
.A(n_3052),
.B(n_371),
.Y(n_3934)
);

AOI21xp5_ASAP7_75t_L g3935 ( 
.A1(n_3047),
.A2(n_372),
.B(n_371),
.Y(n_3935)
);

AOI21xp5_ASAP7_75t_L g3936 ( 
.A1(n_3255),
.A2(n_373),
.B(n_372),
.Y(n_3936)
);

NAND2xp5_ASAP7_75t_SL g3937 ( 
.A(n_3371),
.B(n_3175),
.Y(n_3937)
);

NAND2xp5_ASAP7_75t_L g3938 ( 
.A(n_3511),
.B(n_3514),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3128),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_L g3940 ( 
.A(n_3516),
.B(n_372),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_3518),
.B(n_373),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3519),
.B(n_374),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3130),
.Y(n_3943)
);

AOI22xp5_ASAP7_75t_L g3944 ( 
.A1(n_3381),
.A2(n_375),
.B1(n_376),
.B2(n_374),
.Y(n_3944)
);

OAI21xp5_ASAP7_75t_L g3945 ( 
.A1(n_3112),
.A2(n_29),
.B(n_30),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_L g3946 ( 
.A(n_3520),
.B(n_374),
.Y(n_3946)
);

NOR2xp33_ASAP7_75t_L g3947 ( 
.A(n_3036),
.B(n_375),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_3522),
.B(n_375),
.Y(n_3948)
);

AOI21xp5_ASAP7_75t_L g3949 ( 
.A1(n_3437),
.A2(n_377),
.B(n_376),
.Y(n_3949)
);

INVx2_ASAP7_75t_SL g3950 ( 
.A(n_3088),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3225),
.Y(n_3951)
);

AND2x2_ASAP7_75t_SL g3952 ( 
.A(n_3230),
.B(n_376),
.Y(n_3952)
);

INVx2_ASAP7_75t_L g3953 ( 
.A(n_3091),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3133),
.Y(n_3954)
);

OAI21xp5_ASAP7_75t_L g3955 ( 
.A1(n_3118),
.A2(n_29),
.B(n_30),
.Y(n_3955)
);

NOR2xp33_ASAP7_75t_SL g3956 ( 
.A(n_3166),
.B(n_377),
.Y(n_3956)
);

INVx2_ASAP7_75t_L g3957 ( 
.A(n_3103),
.Y(n_3957)
);

OR2x2_ASAP7_75t_L g3958 ( 
.A(n_3035),
.B(n_378),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_3527),
.B(n_379),
.Y(n_3959)
);

AND2x2_ASAP7_75t_L g3960 ( 
.A(n_3254),
.B(n_379),
.Y(n_3960)
);

INVx2_ASAP7_75t_L g3961 ( 
.A(n_3145),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_SL g3962 ( 
.A(n_3175),
.B(n_381),
.Y(n_3962)
);

NOR2xp67_ASAP7_75t_L g3963 ( 
.A(n_3619),
.B(n_382),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_L g3964 ( 
.A(n_3528),
.B(n_382),
.Y(n_3964)
);

AOI21xp5_ASAP7_75t_L g3965 ( 
.A1(n_3246),
.A2(n_384),
.B(n_383),
.Y(n_3965)
);

NOR2xp33_ASAP7_75t_L g3966 ( 
.A(n_3115),
.B(n_383),
.Y(n_3966)
);

AOI21xp5_ASAP7_75t_L g3967 ( 
.A1(n_3311),
.A2(n_384),
.B(n_383),
.Y(n_3967)
);

INVx2_ASAP7_75t_L g3968 ( 
.A(n_3153),
.Y(n_3968)
);

AOI21xp5_ASAP7_75t_L g3969 ( 
.A1(n_3219),
.A2(n_385),
.B(n_384),
.Y(n_3969)
);

BUFx6f_ASAP7_75t_L g3970 ( 
.A(n_3506),
.Y(n_3970)
);

INVx2_ASAP7_75t_L g3971 ( 
.A(n_3158),
.Y(n_3971)
);

NOR2x1_ASAP7_75t_L g3972 ( 
.A(n_3683),
.B(n_1165),
.Y(n_3972)
);

AOI21xp5_ASAP7_75t_L g3973 ( 
.A1(n_3380),
.A2(n_386),
.B(n_385),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_3531),
.B(n_386),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3173),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_L g3976 ( 
.A(n_3532),
.B(n_386),
.Y(n_3976)
);

AND2x2_ASAP7_75t_SL g3977 ( 
.A(n_3525),
.B(n_387),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_SL g3978 ( 
.A(n_3505),
.B(n_387),
.Y(n_3978)
);

INVx2_ASAP7_75t_L g3979 ( 
.A(n_3186),
.Y(n_3979)
);

INVx11_ASAP7_75t_L g3980 ( 
.A(n_3142),
.Y(n_3980)
);

NAND2xp5_ASAP7_75t_L g3981 ( 
.A(n_3535),
.B(n_388),
.Y(n_3981)
);

AND2x4_ASAP7_75t_L g3982 ( 
.A(n_3152),
.B(n_388),
.Y(n_3982)
);

INVx2_ASAP7_75t_L g3983 ( 
.A(n_3194),
.Y(n_3983)
);

BUFx3_ASAP7_75t_L g3984 ( 
.A(n_3170),
.Y(n_3984)
);

HB1xp67_ASAP7_75t_L g3985 ( 
.A(n_3040),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_SL g3986 ( 
.A(n_3423),
.B(n_389),
.Y(n_3986)
);

AOI21xp5_ASAP7_75t_L g3987 ( 
.A1(n_3387),
.A2(n_390),
.B(n_389),
.Y(n_3987)
);

AOI21xp5_ASAP7_75t_L g3988 ( 
.A1(n_3392),
.A2(n_390),
.B(n_389),
.Y(n_3988)
);

AOI21x1_ASAP7_75t_L g3989 ( 
.A1(n_3440),
.A2(n_392),
.B(n_391),
.Y(n_3989)
);

INVx2_ASAP7_75t_L g3990 ( 
.A(n_3203),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_SL g3991 ( 
.A(n_3423),
.B(n_391),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_L g3992 ( 
.A(n_3537),
.B(n_392),
.Y(n_3992)
);

AND2x2_ASAP7_75t_L g3993 ( 
.A(n_3038),
.B(n_393),
.Y(n_3993)
);

NOR2xp33_ASAP7_75t_L g3994 ( 
.A(n_3147),
.B(n_3197),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_3547),
.B(n_393),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_3553),
.B(n_393),
.Y(n_3996)
);

NAND2xp5_ASAP7_75t_L g3997 ( 
.A(n_3554),
.B(n_394),
.Y(n_3997)
);

AOI21xp5_ASAP7_75t_L g3998 ( 
.A1(n_3393),
.A2(n_395),
.B(n_394),
.Y(n_3998)
);

AOI21x1_ASAP7_75t_L g3999 ( 
.A1(n_3441),
.A2(n_395),
.B(n_394),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3206),
.Y(n_4000)
);

AOI21xp5_ASAP7_75t_L g4001 ( 
.A1(n_3400),
.A2(n_396),
.B(n_395),
.Y(n_4001)
);

NOR2xp33_ASAP7_75t_L g4002 ( 
.A(n_3147),
.B(n_396),
.Y(n_4002)
);

INVx2_ASAP7_75t_L g4003 ( 
.A(n_3253),
.Y(n_4003)
);

AOI21xp5_ASAP7_75t_L g4004 ( 
.A1(n_3421),
.A2(n_398),
.B(n_397),
.Y(n_4004)
);

AOI21xp5_ASAP7_75t_L g4005 ( 
.A1(n_3422),
.A2(n_399),
.B(n_397),
.Y(n_4005)
);

AOI22xp5_ASAP7_75t_L g4006 ( 
.A1(n_3079),
.A2(n_400),
.B1(n_401),
.B2(n_397),
.Y(n_4006)
);

NAND2xp5_ASAP7_75t_L g4007 ( 
.A(n_3562),
.B(n_3564),
.Y(n_4007)
);

OAI22xp5_ASAP7_75t_L g4008 ( 
.A1(n_3529),
.A2(n_401),
.B1(n_402),
.B2(n_400),
.Y(n_4008)
);

AND2x2_ASAP7_75t_L g4009 ( 
.A(n_3269),
.B(n_401),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_L g4010 ( 
.A(n_3566),
.B(n_402),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_SL g4011 ( 
.A(n_3438),
.B(n_402),
.Y(n_4011)
);

AO21x1_ASAP7_75t_L g4012 ( 
.A1(n_3592),
.A2(n_404),
.B(n_403),
.Y(n_4012)
);

AOI21xp5_ASAP7_75t_L g4013 ( 
.A1(n_3424),
.A2(n_404),
.B(n_403),
.Y(n_4013)
);

HB1xp67_ASAP7_75t_L g4014 ( 
.A(n_3673),
.Y(n_4014)
);

AOI21xp5_ASAP7_75t_L g4015 ( 
.A1(n_3427),
.A2(n_405),
.B(n_404),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_L g4016 ( 
.A(n_3567),
.B(n_3576),
.Y(n_4016)
);

INVx3_ASAP7_75t_L g4017 ( 
.A(n_3227),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_L g4018 ( 
.A(n_3579),
.B(n_405),
.Y(n_4018)
);

O2A1O1Ixp33_ASAP7_75t_SL g4019 ( 
.A1(n_3548),
.A2(n_407),
.B(n_408),
.C(n_406),
.Y(n_4019)
);

OAI21xp33_ASAP7_75t_L g4020 ( 
.A1(n_3500),
.A2(n_31),
.B(n_32),
.Y(n_4020)
);

AOI21xp5_ASAP7_75t_L g4021 ( 
.A1(n_3132),
.A2(n_407),
.B(n_406),
.Y(n_4021)
);

NOR2xp33_ASAP7_75t_SL g4022 ( 
.A(n_3683),
.B(n_406),
.Y(n_4022)
);

AOI21xp5_ASAP7_75t_L g4023 ( 
.A1(n_3086),
.A2(n_408),
.B(n_407),
.Y(n_4023)
);

OAI22xp5_ASAP7_75t_L g4024 ( 
.A1(n_3534),
.A2(n_410),
.B1(n_411),
.B2(n_409),
.Y(n_4024)
);

NOR3xp33_ASAP7_75t_L g4025 ( 
.A(n_3667),
.B(n_410),
.C(n_409),
.Y(n_4025)
);

O2A1O1Ixp33_ASAP7_75t_L g4026 ( 
.A1(n_3572),
.A2(n_410),
.B(n_411),
.C(n_409),
.Y(n_4026)
);

INVx3_ASAP7_75t_L g4027 ( 
.A(n_3227),
.Y(n_4027)
);

NOR2xp33_ASAP7_75t_L g4028 ( 
.A(n_3151),
.B(n_411),
.Y(n_4028)
);

AND2x2_ASAP7_75t_L g4029 ( 
.A(n_3269),
.B(n_413),
.Y(n_4029)
);

AOI21xp5_ASAP7_75t_L g4030 ( 
.A1(n_3239),
.A2(n_3138),
.B(n_3134),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_L g4031 ( 
.A(n_3594),
.B(n_413),
.Y(n_4031)
);

BUFx6f_ASAP7_75t_L g4032 ( 
.A(n_3506),
.Y(n_4032)
);

AOI21xp5_ASAP7_75t_L g4033 ( 
.A1(n_3319),
.A2(n_414),
.B(n_413),
.Y(n_4033)
);

AND2x2_ASAP7_75t_L g4034 ( 
.A(n_3064),
.B(n_414),
.Y(n_4034)
);

O2A1O1Ixp5_ASAP7_75t_L g4035 ( 
.A1(n_3375),
.A2(n_415),
.B(n_416),
.C(n_414),
.Y(n_4035)
);

AND2x2_ASAP7_75t_L g4036 ( 
.A(n_3463),
.B(n_415),
.Y(n_4036)
);

AOI21xp5_ASAP7_75t_L g4037 ( 
.A1(n_3340),
.A2(n_418),
.B(n_417),
.Y(n_4037)
);

NOR2xp33_ASAP7_75t_L g4038 ( 
.A(n_3149),
.B(n_417),
.Y(n_4038)
);

AOI21xp5_ASAP7_75t_L g4039 ( 
.A1(n_3341),
.A2(n_418),
.B(n_417),
.Y(n_4039)
);

OAI22xp5_ASAP7_75t_L g4040 ( 
.A1(n_3542),
.A2(n_419),
.B1(n_420),
.B2(n_418),
.Y(n_4040)
);

INVx3_ASAP7_75t_L g4041 ( 
.A(n_3317),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_L g4042 ( 
.A(n_3599),
.B(n_419),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_3600),
.B(n_420),
.Y(n_4043)
);

O2A1O1Ixp33_ASAP7_75t_L g4044 ( 
.A1(n_3431),
.A2(n_421),
.B(n_422),
.C(n_420),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_SL g4045 ( 
.A(n_3438),
.B(n_421),
.Y(n_4045)
);

AOI21xp5_ASAP7_75t_L g4046 ( 
.A1(n_3345),
.A2(n_3358),
.B(n_3348),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_L g4047 ( 
.A(n_3601),
.B(n_421),
.Y(n_4047)
);

AOI21xp5_ASAP7_75t_L g4048 ( 
.A1(n_3367),
.A2(n_423),
.B(n_422),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_L g4049 ( 
.A(n_3610),
.B(n_3612),
.Y(n_4049)
);

AOI21xp5_ASAP7_75t_L g4050 ( 
.A1(n_3377),
.A2(n_425),
.B(n_424),
.Y(n_4050)
);

BUFx6f_ASAP7_75t_L g4051 ( 
.A(n_3385),
.Y(n_4051)
);

OAI21xp5_ASAP7_75t_L g4052 ( 
.A1(n_3205),
.A2(n_31),
.B(n_32),
.Y(n_4052)
);

AND2x2_ASAP7_75t_L g4053 ( 
.A(n_3041),
.B(n_424),
.Y(n_4053)
);

AOI21x1_ASAP7_75t_L g4054 ( 
.A1(n_3442),
.A2(n_425),
.B(n_424),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_L g4055 ( 
.A(n_3618),
.B(n_425),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_L g4056 ( 
.A(n_3621),
.B(n_426),
.Y(n_4056)
);

O2A1O1Ixp5_ASAP7_75t_L g4057 ( 
.A1(n_3378),
.A2(n_427),
.B(n_428),
.C(n_426),
.Y(n_4057)
);

INVx3_ASAP7_75t_L g4058 ( 
.A(n_3317),
.Y(n_4058)
);

NOR2xp33_ASAP7_75t_SL g4059 ( 
.A(n_3142),
.B(n_426),
.Y(n_4059)
);

OAI21xp5_ASAP7_75t_L g4060 ( 
.A1(n_3330),
.A2(n_31),
.B(n_32),
.Y(n_4060)
);

AOI22xp5_ASAP7_75t_L g4061 ( 
.A1(n_3082),
.A2(n_429),
.B1(n_430),
.B2(n_427),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3226),
.Y(n_4062)
);

OAI21xp5_ASAP7_75t_L g4063 ( 
.A1(n_3330),
.A2(n_33),
.B(n_34),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_3622),
.B(n_427),
.Y(n_4064)
);

A2O1A1Ixp33_ASAP7_75t_L g4065 ( 
.A1(n_3501),
.A2(n_35),
.B(n_33),
.C(n_34),
.Y(n_4065)
);

A2O1A1Ixp33_ASAP7_75t_L g4066 ( 
.A1(n_3503),
.A2(n_35),
.B(n_33),
.C(n_34),
.Y(n_4066)
);

O2A1O1Ixp33_ASAP7_75t_L g4067 ( 
.A1(n_3550),
.A2(n_3558),
.B(n_3580),
.C(n_3557),
.Y(n_4067)
);

A2O1A1Ixp33_ASAP7_75t_L g4068 ( 
.A1(n_3552),
.A2(n_36),
.B(n_33),
.C(n_35),
.Y(n_4068)
);

AOI21xp5_ASAP7_75t_L g4069 ( 
.A1(n_3379),
.A2(n_430),
.B(n_429),
.Y(n_4069)
);

NAND2xp5_ASAP7_75t_SL g4070 ( 
.A(n_3385),
.B(n_429),
.Y(n_4070)
);

A2O1A1Ixp33_ASAP7_75t_L g4071 ( 
.A1(n_3559),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_4071)
);

AOI21xp5_ASAP7_75t_L g4072 ( 
.A1(n_3286),
.A2(n_431),
.B(n_430),
.Y(n_4072)
);

AND2x2_ASAP7_75t_L g4073 ( 
.A(n_3235),
.B(n_3419),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3229),
.Y(n_4074)
);

NAND3xp33_ASAP7_75t_L g4075 ( 
.A(n_3672),
.B(n_432),
.C(n_431),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_L g4076 ( 
.A(n_3625),
.B(n_432),
.Y(n_4076)
);

NOR2xp33_ASAP7_75t_L g4077 ( 
.A(n_3217),
.B(n_433),
.Y(n_4077)
);

OAI21xp33_ASAP7_75t_L g4078 ( 
.A1(n_3561),
.A2(n_36),
.B(n_37),
.Y(n_4078)
);

NAND2xp5_ASAP7_75t_SL g4079 ( 
.A(n_3385),
.B(n_433),
.Y(n_4079)
);

NAND2xp5_ASAP7_75t_L g4080 ( 
.A(n_3638),
.B(n_434),
.Y(n_4080)
);

AND2x2_ASAP7_75t_L g4081 ( 
.A(n_3200),
.B(n_434),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3642),
.B(n_434),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_L g4083 ( 
.A(n_3650),
.B(n_3657),
.Y(n_4083)
);

NOR2xp33_ASAP7_75t_L g4084 ( 
.A(n_3491),
.B(n_435),
.Y(n_4084)
);

O2A1O1Ixp33_ASAP7_75t_L g4085 ( 
.A1(n_3584),
.A2(n_436),
.B(n_437),
.C(n_435),
.Y(n_4085)
);

BUFx3_ASAP7_75t_L g4086 ( 
.A(n_3170),
.Y(n_4086)
);

NAND2xp5_ASAP7_75t_L g4087 ( 
.A(n_3661),
.B(n_435),
.Y(n_4087)
);

NAND2xp5_ASAP7_75t_L g4088 ( 
.A(n_3669),
.B(n_436),
.Y(n_4088)
);

AND2x2_ASAP7_75t_L g4089 ( 
.A(n_3450),
.B(n_436),
.Y(n_4089)
);

INVx2_ASAP7_75t_L g4090 ( 
.A(n_3260),
.Y(n_4090)
);

AND2x2_ASAP7_75t_L g4091 ( 
.A(n_3450),
.B(n_437),
.Y(n_4091)
);

AOI21x1_ASAP7_75t_L g4092 ( 
.A1(n_3443),
.A2(n_438),
.B(n_437),
.Y(n_4092)
);

AOI21xp5_ASAP7_75t_L g4093 ( 
.A1(n_3327),
.A2(n_439),
.B(n_438),
.Y(n_4093)
);

AND2x2_ASAP7_75t_L g4094 ( 
.A(n_3195),
.B(n_438),
.Y(n_4094)
);

NAND2x1p5_ASAP7_75t_L g4095 ( 
.A(n_3081),
.B(n_439),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_L g4096 ( 
.A(n_3681),
.B(n_440),
.Y(n_4096)
);

AOI21xp5_ASAP7_75t_L g4097 ( 
.A1(n_3396),
.A2(n_441),
.B(n_440),
.Y(n_4097)
);

BUFx6f_ASAP7_75t_L g4098 ( 
.A(n_3169),
.Y(n_4098)
);

NOR2xp67_ASAP7_75t_L g4099 ( 
.A(n_3074),
.B(n_441),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_3682),
.B(n_3687),
.Y(n_4100)
);

NAND2xp5_ASAP7_75t_L g4101 ( 
.A(n_3688),
.B(n_441),
.Y(n_4101)
);

HB1xp67_ASAP7_75t_L g4102 ( 
.A(n_3693),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_SL g4103 ( 
.A(n_3256),
.B(n_442),
.Y(n_4103)
);

AND2x2_ASAP7_75t_L g4104 ( 
.A(n_3310),
.B(n_3389),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_3247),
.Y(n_4105)
);

NOR2xp33_ASAP7_75t_L g4106 ( 
.A(n_3224),
.B(n_442),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_L g4107 ( 
.A(n_3695),
.B(n_443),
.Y(n_4107)
);

AOI21xp5_ASAP7_75t_L g4108 ( 
.A1(n_3413),
.A2(n_444),
.B(n_443),
.Y(n_4108)
);

AOI21xp5_ASAP7_75t_L g4109 ( 
.A1(n_3334),
.A2(n_445),
.B(n_444),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_L g4110 ( 
.A(n_3702),
.B(n_444),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_L g4111 ( 
.A(n_3703),
.B(n_445),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_3709),
.B(n_445),
.Y(n_4112)
);

OAI21xp5_ASAP7_75t_L g4113 ( 
.A1(n_3448),
.A2(n_37),
.B(n_38),
.Y(n_4113)
);

INVx2_ASAP7_75t_L g4114 ( 
.A(n_3264),
.Y(n_4114)
);

AND2x2_ASAP7_75t_L g4115 ( 
.A(n_3310),
.B(n_446),
.Y(n_4115)
);

AOI21xp5_ASAP7_75t_L g4116 ( 
.A1(n_3346),
.A2(n_447),
.B(n_446),
.Y(n_4116)
);

AOI22xp5_ASAP7_75t_L g4117 ( 
.A1(n_3240),
.A2(n_448),
.B1(n_449),
.B2(n_447),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_L g4118 ( 
.A(n_3313),
.B(n_447),
.Y(n_4118)
);

AOI21xp5_ASAP7_75t_L g4119 ( 
.A1(n_3353),
.A2(n_3355),
.B(n_3354),
.Y(n_4119)
);

INVx2_ASAP7_75t_L g4120 ( 
.A(n_3287),
.Y(n_4120)
);

BUFx2_ASAP7_75t_L g4121 ( 
.A(n_3309),
.Y(n_4121)
);

NOR2xp33_ASAP7_75t_L g4122 ( 
.A(n_3373),
.B(n_448),
.Y(n_4122)
);

AOI21xp5_ASAP7_75t_L g4123 ( 
.A1(n_3356),
.A2(n_450),
.B(n_449),
.Y(n_4123)
);

A2O1A1Ixp33_ASAP7_75t_L g4124 ( 
.A1(n_3571),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_4124)
);

AOI21xp5_ASAP7_75t_L g4125 ( 
.A1(n_3308),
.A2(n_451),
.B(n_450),
.Y(n_4125)
);

AO21x1_ASAP7_75t_L g4126 ( 
.A1(n_3616),
.A2(n_452),
.B(n_451),
.Y(n_4126)
);

AOI21x1_ASAP7_75t_L g4127 ( 
.A1(n_3464),
.A2(n_3467),
.B(n_3465),
.Y(n_4127)
);

HB1xp67_ASAP7_75t_L g4128 ( 
.A(n_3275),
.Y(n_4128)
);

AOI21xp5_ASAP7_75t_L g4129 ( 
.A1(n_3211),
.A2(n_453),
.B(n_452),
.Y(n_4129)
);

AOI21xp5_ASAP7_75t_L g4130 ( 
.A1(n_3211),
.A2(n_455),
.B(n_454),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_3078),
.B(n_454),
.Y(n_4131)
);

BUFx6f_ASAP7_75t_L g4132 ( 
.A(n_3169),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_3266),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_3284),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_SL g4135 ( 
.A(n_3256),
.B(n_455),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_3332),
.B(n_455),
.Y(n_4136)
);

NAND2x1p5_ASAP7_75t_L g4137 ( 
.A(n_3410),
.B(n_456),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_L g4138 ( 
.A(n_3595),
.B(n_456),
.Y(n_4138)
);

NOR2xp33_ASAP7_75t_L g4139 ( 
.A(n_3107),
.B(n_456),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_3604),
.B(n_457),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_L g4141 ( 
.A(n_3613),
.B(n_3620),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_3623),
.B(n_457),
.Y(n_4142)
);

NOR2x1p5_ASAP7_75t_L g4143 ( 
.A(n_3636),
.B(n_458),
.Y(n_4143)
);

CKINVDCx20_ASAP7_75t_R g4144 ( 
.A(n_3274),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_SL g4145 ( 
.A(n_3533),
.B(n_458),
.Y(n_4145)
);

AOI21xp5_ASAP7_75t_L g4146 ( 
.A1(n_3426),
.A2(n_3439),
.B(n_3291),
.Y(n_4146)
);

OAI21xp5_ASAP7_75t_L g4147 ( 
.A1(n_3231),
.A2(n_39),
.B(n_40),
.Y(n_4147)
);

AOI33xp33_ASAP7_75t_L g4148 ( 
.A1(n_3696),
.A2(n_461),
.A3(n_459),
.B1(n_462),
.B2(n_460),
.B3(n_458),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_L g4149 ( 
.A(n_3634),
.B(n_459),
.Y(n_4149)
);

AOI21xp5_ASAP7_75t_L g4150 ( 
.A1(n_3288),
.A2(n_3407),
.B(n_3053),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_SL g4151 ( 
.A(n_3575),
.B(n_3652),
.Y(n_4151)
);

AOI21xp5_ASAP7_75t_L g4152 ( 
.A1(n_3048),
.A2(n_460),
.B(n_459),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_SL g4153 ( 
.A(n_3665),
.B(n_460),
.Y(n_4153)
);

AOI22xp5_ASAP7_75t_L g4154 ( 
.A1(n_3641),
.A2(n_462),
.B1(n_464),
.B2(n_461),
.Y(n_4154)
);

AND2x2_ASAP7_75t_L g4155 ( 
.A(n_3662),
.B(n_461),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_3663),
.B(n_462),
.Y(n_4156)
);

BUFx3_ASAP7_75t_L g4157 ( 
.A(n_3170),
.Y(n_4157)
);

AOI21xp5_ASAP7_75t_L g4158 ( 
.A1(n_3057),
.A2(n_465),
.B(n_464),
.Y(n_4158)
);

AOI21xp5_ASAP7_75t_L g4159 ( 
.A1(n_3059),
.A2(n_465),
.B(n_464),
.Y(n_4159)
);

OR2x2_ASAP7_75t_L g4160 ( 
.A(n_3272),
.B(n_466),
.Y(n_4160)
);

AOI21xp5_ASAP7_75t_L g4161 ( 
.A1(n_3062),
.A2(n_467),
.B(n_466),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_L g4162 ( 
.A(n_3677),
.B(n_466),
.Y(n_4162)
);

AOI21xp33_ASAP7_75t_L g4163 ( 
.A1(n_3312),
.A2(n_468),
.B(n_467),
.Y(n_4163)
);

NOR2xp33_ASAP7_75t_L g4164 ( 
.A(n_3114),
.B(n_3198),
.Y(n_4164)
);

AOI21xp5_ASAP7_75t_L g4165 ( 
.A1(n_3065),
.A2(n_469),
.B(n_468),
.Y(n_4165)
);

NAND2xp5_ASAP7_75t_L g4166 ( 
.A(n_3679),
.B(n_468),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_3401),
.Y(n_4167)
);

OAI21xp33_ASAP7_75t_SL g4168 ( 
.A1(n_3570),
.A2(n_3643),
.B(n_3586),
.Y(n_4168)
);

NAND2xp5_ASAP7_75t_L g4169 ( 
.A(n_3698),
.B(n_470),
.Y(n_4169)
);

AND2x2_ASAP7_75t_L g4170 ( 
.A(n_3333),
.B(n_470),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_L g4171 ( 
.A(n_3704),
.B(n_470),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_SL g4172 ( 
.A(n_3700),
.B(n_471),
.Y(n_4172)
);

AOI22x1_ASAP7_75t_L g4173 ( 
.A1(n_3480),
.A2(n_472),
.B1(n_473),
.B2(n_471),
.Y(n_4173)
);

A2O1A1Ixp33_ASAP7_75t_L g4174 ( 
.A1(n_3644),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_4174)
);

NOR2xp33_ASAP7_75t_L g4175 ( 
.A(n_3208),
.B(n_472),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_SL g4176 ( 
.A(n_3097),
.B(n_473),
.Y(n_4176)
);

AND2x4_ASAP7_75t_L g4177 ( 
.A(n_3172),
.B(n_473),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_L g4178 ( 
.A(n_3314),
.B(n_3089),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_SL g4179 ( 
.A(n_3097),
.B(n_474),
.Y(n_4179)
);

OAI21x1_ASAP7_75t_L g4180 ( 
.A1(n_3249),
.A2(n_475),
.B(n_474),
.Y(n_4180)
);

OR2x2_ASAP7_75t_L g4181 ( 
.A(n_3092),
.B(n_474),
.Y(n_4181)
);

AOI21xp5_ASAP7_75t_L g4182 ( 
.A1(n_3068),
.A2(n_476),
.B(n_475),
.Y(n_4182)
);

OAI321xp33_ASAP7_75t_L g4183 ( 
.A1(n_3573),
.A2(n_3632),
.A3(n_3586),
.B1(n_3678),
.B2(n_3647),
.C(n_3643),
.Y(n_4183)
);

BUFx6f_ASAP7_75t_L g4184 ( 
.A(n_3169),
.Y(n_4184)
);

OAI21xp5_ASAP7_75t_L g4185 ( 
.A1(n_3236),
.A2(n_39),
.B(n_40),
.Y(n_4185)
);

NAND2xp5_ASAP7_75t_L g4186 ( 
.A(n_3325),
.B(n_475),
.Y(n_4186)
);

O2A1O1Ixp5_ASAP7_75t_L g4187 ( 
.A1(n_3329),
.A2(n_477),
.B(n_478),
.C(n_476),
.Y(n_4187)
);

AND2x2_ASAP7_75t_L g4188 ( 
.A(n_3184),
.B(n_476),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_3339),
.B(n_477),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_L g4190 ( 
.A(n_3668),
.B(n_477),
.Y(n_4190)
);

HB1xp67_ASAP7_75t_L g4191 ( 
.A(n_3309),
.Y(n_4191)
);

INVx2_ASAP7_75t_L g4192 ( 
.A(n_3294),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_3404),
.Y(n_4193)
);

AOI21xp5_ASAP7_75t_L g4194 ( 
.A1(n_3069),
.A2(n_479),
.B(n_478),
.Y(n_4194)
);

AOI21xp5_ASAP7_75t_L g4195 ( 
.A1(n_3070),
.A2(n_480),
.B(n_478),
.Y(n_4195)
);

NAND2xp5_ASAP7_75t_L g4196 ( 
.A(n_3674),
.B(n_480),
.Y(n_4196)
);

AND2x2_ASAP7_75t_L g4197 ( 
.A(n_3184),
.B(n_481),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_L g4198 ( 
.A(n_3699),
.B(n_481),
.Y(n_4198)
);

AOI21xp5_ASAP7_75t_L g4199 ( 
.A1(n_3263),
.A2(n_483),
.B(n_482),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_L g4200 ( 
.A(n_3493),
.B(n_482),
.Y(n_4200)
);

AOI21xp5_ASAP7_75t_L g4201 ( 
.A1(n_3265),
.A2(n_483),
.B(n_482),
.Y(n_4201)
);

NAND2xp5_ASAP7_75t_L g4202 ( 
.A(n_3119),
.B(n_483),
.Y(n_4202)
);

AOI21xp5_ASAP7_75t_L g4203 ( 
.A1(n_3268),
.A2(n_485),
.B(n_484),
.Y(n_4203)
);

AOI21xp5_ASAP7_75t_L g4204 ( 
.A1(n_3273),
.A2(n_485),
.B(n_484),
.Y(n_4204)
);

BUFx3_ASAP7_75t_L g4205 ( 
.A(n_3181),
.Y(n_4205)
);

OAI21xp33_ASAP7_75t_L g4206 ( 
.A1(n_3386),
.A2(n_41),
.B(n_42),
.Y(n_4206)
);

OAI21xp5_ASAP7_75t_L g4207 ( 
.A1(n_3279),
.A2(n_42),
.B(n_43),
.Y(n_4207)
);

NOR2xp33_ASAP7_75t_L g4208 ( 
.A(n_3228),
.B(n_484),
.Y(n_4208)
);

HB1xp67_ASAP7_75t_L g4209 ( 
.A(n_3309),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_3271),
.B(n_3139),
.Y(n_4210)
);

AOI21xp5_ASAP7_75t_L g4211 ( 
.A1(n_3453),
.A2(n_486),
.B(n_485),
.Y(n_4211)
);

NOR3xp33_ASAP7_75t_L g4212 ( 
.A(n_3626),
.B(n_487),
.C(n_486),
.Y(n_4212)
);

BUFx6f_ASAP7_75t_L g4213 ( 
.A(n_3181),
.Y(n_4213)
);

INVx4_ASAP7_75t_L g4214 ( 
.A(n_3181),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_3141),
.B(n_486),
.Y(n_4215)
);

AND2x2_ASAP7_75t_L g4216 ( 
.A(n_3094),
.B(n_487),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_3155),
.B(n_487),
.Y(n_4217)
);

HB1xp67_ASAP7_75t_L g4218 ( 
.A(n_3167),
.Y(n_4218)
);

AOI21xp5_ASAP7_75t_L g4219 ( 
.A1(n_3507),
.A2(n_489),
.B(n_488),
.Y(n_4219)
);

AOI21xp5_ASAP7_75t_L g4220 ( 
.A1(n_3515),
.A2(n_489),
.B(n_488),
.Y(n_4220)
);

BUFx6f_ASAP7_75t_L g4221 ( 
.A(n_3299),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_3163),
.B(n_490),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_L g4223 ( 
.A(n_3165),
.B(n_490),
.Y(n_4223)
);

INVx3_ASAP7_75t_L g4224 ( 
.A(n_3428),
.Y(n_4224)
);

INVx2_ASAP7_75t_L g4225 ( 
.A(n_3300),
.Y(n_4225)
);

OAI21xp5_ASAP7_75t_L g4226 ( 
.A1(n_3160),
.A2(n_42),
.B(n_43),
.Y(n_4226)
);

INVx1_ASAP7_75t_L g4227 ( 
.A(n_3323),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_L g4228 ( 
.A(n_3174),
.B(n_491),
.Y(n_4228)
);

BUFx6f_ASAP7_75t_L g4229 ( 
.A(n_3299),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_3366),
.Y(n_4230)
);

AOI21xp5_ASAP7_75t_L g4231 ( 
.A1(n_3544),
.A2(n_492),
.B(n_491),
.Y(n_4231)
);

AOI21xp5_ASAP7_75t_L g4232 ( 
.A1(n_3349),
.A2(n_3403),
.B(n_3270),
.Y(n_4232)
);

INVx4_ASAP7_75t_L g4233 ( 
.A(n_3299),
.Y(n_4233)
);

OAI21xp5_ASAP7_75t_L g4234 ( 
.A1(n_3409),
.A2(n_42),
.B(n_43),
.Y(n_4234)
);

INVx1_ASAP7_75t_SL g4235 ( 
.A(n_3196),
.Y(n_4235)
);

NAND2xp5_ASAP7_75t_L g4236 ( 
.A(n_3176),
.B(n_3285),
.Y(n_4236)
);

NAND2xp33_ASAP7_75t_L g4237 ( 
.A(n_3637),
.B(n_491),
.Y(n_4237)
);

OAI21xp5_ASAP7_75t_L g4238 ( 
.A1(n_3343),
.A2(n_43),
.B(n_44),
.Y(n_4238)
);

OAI21xp33_ASAP7_75t_L g4239 ( 
.A1(n_3390),
.A2(n_44),
.B(n_45),
.Y(n_4239)
);

AOI21xp5_ASAP7_75t_L g4240 ( 
.A1(n_3295),
.A2(n_493),
.B(n_492),
.Y(n_4240)
);

AOI21xp5_ASAP7_75t_L g4241 ( 
.A1(n_3347),
.A2(n_494),
.B(n_493),
.Y(n_4241)
);

A2O1A1Ixp33_ASAP7_75t_L g4242 ( 
.A1(n_3363),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_4242)
);

AOI33xp33_ASAP7_75t_L g4243 ( 
.A1(n_3434),
.A2(n_496),
.A3(n_494),
.B1(n_497),
.B2(n_495),
.B3(n_493),
.Y(n_4243)
);

AOI21x1_ASAP7_75t_L g4244 ( 
.A1(n_3469),
.A2(n_495),
.B(n_494),
.Y(n_4244)
);

HB1xp67_ASAP7_75t_L g4245 ( 
.A(n_3648),
.Y(n_4245)
);

AND2x2_ASAP7_75t_L g4246 ( 
.A(n_3468),
.B(n_495),
.Y(n_4246)
);

AOI21xp5_ASAP7_75t_L g4247 ( 
.A1(n_3350),
.A2(n_497),
.B(n_496),
.Y(n_4247)
);

AND2x2_ASAP7_75t_L g4248 ( 
.A(n_3664),
.B(n_496),
.Y(n_4248)
);

NAND2xp5_ASAP7_75t_SL g4249 ( 
.A(n_3637),
.B(n_497),
.Y(n_4249)
);

OAI22xp5_ASAP7_75t_L g4250 ( 
.A1(n_3647),
.A2(n_499),
.B1(n_500),
.B2(n_498),
.Y(n_4250)
);

OAI21xp5_ASAP7_75t_L g4251 ( 
.A1(n_3344),
.A2(n_45),
.B(n_46),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_L g4252 ( 
.A(n_3242),
.B(n_498),
.Y(n_4252)
);

OAI21xp33_ASAP7_75t_L g4253 ( 
.A1(n_3382),
.A2(n_46),
.B(n_47),
.Y(n_4253)
);

BUFx6f_ASAP7_75t_L g4254 ( 
.A(n_3480),
.Y(n_4254)
);

AOI21xp5_ASAP7_75t_L g4255 ( 
.A1(n_3326),
.A2(n_499),
.B(n_498),
.Y(n_4255)
);

NOR2xp67_ASAP7_75t_L g4256 ( 
.A(n_3539),
.B(n_500),
.Y(n_4256)
);

AOI21x1_ASAP7_75t_L g4257 ( 
.A1(n_3478),
.A2(n_501),
.B(n_500),
.Y(n_4257)
);

A2O1A1Ixp33_ASAP7_75t_L g4258 ( 
.A1(n_3201),
.A2(n_48),
.B(n_46),
.C(n_47),
.Y(n_4258)
);

NAND2x1p5_ASAP7_75t_L g4259 ( 
.A(n_3104),
.B(n_501),
.Y(n_4259)
);

AOI21xp5_ASAP7_75t_L g4260 ( 
.A1(n_3331),
.A2(n_502),
.B(n_501),
.Y(n_4260)
);

NAND2xp5_ASAP7_75t_L g4261 ( 
.A(n_3352),
.B(n_502),
.Y(n_4261)
);

AOI21xp5_ASAP7_75t_L g4262 ( 
.A1(n_3342),
.A2(n_503),
.B(n_502),
.Y(n_4262)
);

AOI21xp5_ASAP7_75t_L g4263 ( 
.A1(n_3357),
.A2(n_3445),
.B(n_3433),
.Y(n_4263)
);

BUFx6f_ASAP7_75t_L g4264 ( 
.A(n_3428),
.Y(n_4264)
);

OAI22xp5_ASAP7_75t_L g4265 ( 
.A1(n_3678),
.A2(n_504),
.B1(n_505),
.B2(n_503),
.Y(n_4265)
);

A2O1A1Ixp33_ASAP7_75t_L g4266 ( 
.A1(n_3692),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_4266)
);

OAI22xp5_ASAP7_75t_L g4267 ( 
.A1(n_3692),
.A2(n_505),
.B1(n_506),
.B2(n_504),
.Y(n_4267)
);

NOR2xp33_ASAP7_75t_L g4268 ( 
.A(n_3281),
.B(n_504),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_3257),
.B(n_505),
.Y(n_4269)
);

OAI21xp5_ASAP7_75t_L g4270 ( 
.A1(n_3335),
.A2(n_47),
.B(n_48),
.Y(n_4270)
);

INVx2_ASAP7_75t_L g4271 ( 
.A(n_3259),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_L g4272 ( 
.A(n_3087),
.B(n_3215),
.Y(n_4272)
);

NOR2xp33_ASAP7_75t_L g4273 ( 
.A(n_3185),
.B(n_506),
.Y(n_4273)
);

AOI21xp5_ASAP7_75t_L g4274 ( 
.A1(n_3301),
.A2(n_507),
.B(n_506),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_L g4275 ( 
.A(n_3189),
.B(n_507),
.Y(n_4275)
);

O2A1O1Ixp33_ASAP7_75t_L g4276 ( 
.A1(n_3587),
.A2(n_508),
.B(n_509),
.C(n_507),
.Y(n_4276)
);

OAI21xp5_ASAP7_75t_L g4277 ( 
.A1(n_3296),
.A2(n_49),
.B(n_50),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_SL g4278 ( 
.A(n_3637),
.B(n_508),
.Y(n_4278)
);

OAI321xp33_ASAP7_75t_L g4279 ( 
.A1(n_3705),
.A2(n_3238),
.A3(n_3159),
.B1(n_3624),
.B2(n_3609),
.C(n_3591),
.Y(n_4279)
);

INVx1_ASAP7_75t_SL g4280 ( 
.A(n_3135),
.Y(n_4280)
);

OR2x6_ASAP7_75t_L g4281 ( 
.A(n_3569),
.B(n_508),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_L g4282 ( 
.A(n_3214),
.B(n_509),
.Y(n_4282)
);

OAI21xp5_ASAP7_75t_L g4283 ( 
.A1(n_3298),
.A2(n_49),
.B(n_50),
.Y(n_4283)
);

NOR3xp33_ASAP7_75t_L g4284 ( 
.A(n_3627),
.B(n_3635),
.C(n_3630),
.Y(n_4284)
);

NAND2xp5_ASAP7_75t_L g4285 ( 
.A(n_3388),
.B(n_509),
.Y(n_4285)
);

NOR2xp33_ASAP7_75t_L g4286 ( 
.A(n_3164),
.B(n_510),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_SL g4287 ( 
.A(n_3637),
.B(n_510),
.Y(n_4287)
);

BUFx6f_ASAP7_75t_L g4288 ( 
.A(n_3113),
.Y(n_4288)
);

AOI21xp5_ASAP7_75t_L g4289 ( 
.A1(n_3316),
.A2(n_511),
.B(n_510),
.Y(n_4289)
);

AND2x4_ASAP7_75t_L g4290 ( 
.A(n_3172),
.B(n_512),
.Y(n_4290)
);

INVx3_ASAP7_75t_L g4291 ( 
.A(n_3113),
.Y(n_4291)
);

NAND2xp5_ASAP7_75t_L g4292 ( 
.A(n_3364),
.B(n_512),
.Y(n_4292)
);

AOI21xp5_ASAP7_75t_L g4293 ( 
.A1(n_3656),
.A2(n_513),
.B(n_512),
.Y(n_4293)
);

OAI22xp5_ASAP7_75t_L g4294 ( 
.A1(n_3915),
.A2(n_3489),
.B1(n_3492),
.B2(n_3414),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_L g4295 ( 
.A(n_3717),
.B(n_3315),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_SL g4296 ( 
.A(n_3834),
.B(n_3297),
.Y(n_4296)
);

AOI21xp5_ASAP7_75t_L g4297 ( 
.A1(n_3810),
.A2(n_3479),
.B(n_3476),
.Y(n_4297)
);

AND2x2_ASAP7_75t_L g4298 ( 
.A(n_4104),
.B(n_3498),
.Y(n_4298)
);

NAND2xp5_ASAP7_75t_SL g4299 ( 
.A(n_3895),
.B(n_3384),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_3721),
.Y(n_4300)
);

INVx5_ASAP7_75t_L g4301 ( 
.A(n_3794),
.Y(n_4301)
);

AOI21xp5_ASAP7_75t_L g4302 ( 
.A1(n_3930),
.A2(n_3479),
.B(n_3436),
.Y(n_4302)
);

NAND2xp5_ASAP7_75t_L g4303 ( 
.A(n_4073),
.B(n_3429),
.Y(n_4303)
);

BUFx3_ASAP7_75t_L g4304 ( 
.A(n_4144),
.Y(n_4304)
);

BUFx6f_ASAP7_75t_L g4305 ( 
.A(n_3723),
.Y(n_4305)
);

AND2x2_ASAP7_75t_L g4306 ( 
.A(n_3852),
.B(n_3402),
.Y(n_4306)
);

A2O1A1Ixp33_ASAP7_75t_L g4307 ( 
.A1(n_4168),
.A2(n_3483),
.B(n_3666),
.C(n_3660),
.Y(n_4307)
);

A2O1A1Ixp33_ASAP7_75t_L g4308 ( 
.A1(n_3966),
.A2(n_3676),
.B(n_3685),
.C(n_3670),
.Y(n_4308)
);

O2A1O1Ixp33_ASAP7_75t_L g4309 ( 
.A1(n_4141),
.A2(n_3694),
.B(n_3706),
.C(n_3686),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_SL g4310 ( 
.A(n_4121),
.B(n_3761),
.Y(n_4310)
);

NOR2xp33_ASAP7_75t_L g4311 ( 
.A(n_3994),
.B(n_3207),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_3736),
.Y(n_4312)
);

AOI22xp33_ASAP7_75t_L g4313 ( 
.A1(n_4025),
.A2(n_3391),
.B1(n_3435),
.B2(n_3336),
.Y(n_4313)
);

AOI21xp5_ASAP7_75t_L g4314 ( 
.A1(n_4237),
.A2(n_3457),
.B(n_3523),
.Y(n_4314)
);

NOR2xp33_ASAP7_75t_L g4315 ( 
.A(n_3854),
.B(n_3207),
.Y(n_4315)
);

NAND2xp5_ASAP7_75t_SL g4316 ( 
.A(n_4022),
.B(n_3637),
.Y(n_4316)
);

BUFx3_ASAP7_75t_L g4317 ( 
.A(n_3766),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_L g4318 ( 
.A(n_3937),
.B(n_3248),
.Y(n_4318)
);

OAI21x1_ASAP7_75t_L g4319 ( 
.A1(n_4127),
.A2(n_3556),
.B(n_3523),
.Y(n_4319)
);

NOR2xp33_ASAP7_75t_L g4320 ( 
.A(n_3755),
.B(n_3629),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_3745),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_L g4322 ( 
.A(n_4178),
.B(n_3444),
.Y(n_4322)
);

AOI21xp5_ASAP7_75t_L g4323 ( 
.A1(n_3778),
.A2(n_3770),
.B(n_3728),
.Y(n_4323)
);

NOR2xp33_ASAP7_75t_L g4324 ( 
.A(n_3725),
.B(n_3931),
.Y(n_4324)
);

A2O1A1Ixp33_ASAP7_75t_L g4325 ( 
.A1(n_4077),
.A2(n_3477),
.B(n_3474),
.C(n_3470),
.Y(n_4325)
);

AO21x2_ASAP7_75t_L g4326 ( 
.A1(n_4176),
.A2(n_3376),
.B(n_3454),
.Y(n_4326)
);

O2A1O1Ixp33_ASAP7_75t_L g4327 ( 
.A1(n_4236),
.A2(n_3416),
.B(n_3425),
.C(n_3418),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_3756),
.B(n_3321),
.Y(n_4328)
);

A2O1A1Ixp33_ASAP7_75t_L g4329 ( 
.A1(n_4106),
.A2(n_3472),
.B(n_3481),
.C(n_3459),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_SL g4330 ( 
.A(n_4254),
.B(n_3475),
.Y(n_4330)
);

BUFx6f_ASAP7_75t_L g4331 ( 
.A(n_3723),
.Y(n_4331)
);

AOI22xp5_ASAP7_75t_L g4332 ( 
.A1(n_4143),
.A2(n_3218),
.B1(n_3261),
.B2(n_3276),
.Y(n_4332)
);

OAI22xp33_ASAP7_75t_L g4333 ( 
.A1(n_4281),
.A2(n_3305),
.B1(n_3710),
.B2(n_3629),
.Y(n_4333)
);

AOI21xp5_ASAP7_75t_L g4334 ( 
.A1(n_4146),
.A2(n_3590),
.B(n_3556),
.Y(n_4334)
);

OAI21xp33_ASAP7_75t_SL g4335 ( 
.A1(n_3767),
.A2(n_3365),
.B(n_3359),
.Y(n_4335)
);

OAI22xp5_ASAP7_75t_L g4336 ( 
.A1(n_4266),
.A2(n_3397),
.B1(n_3302),
.B2(n_3432),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_L g4337 ( 
.A(n_4227),
.B(n_3351),
.Y(n_4337)
);

CKINVDCx5p33_ASAP7_75t_R g4338 ( 
.A(n_3980),
.Y(n_4338)
);

NAND2xp5_ASAP7_75t_L g4339 ( 
.A(n_4115),
.B(n_3462),
.Y(n_4339)
);

BUFx3_ASAP7_75t_L g4340 ( 
.A(n_3845),
.Y(n_4340)
);

AOI22xp33_ASAP7_75t_L g4341 ( 
.A1(n_4212),
.A2(n_3435),
.B1(n_3336),
.B2(n_3398),
.Y(n_4341)
);

AOI21xp5_ASAP7_75t_L g4342 ( 
.A1(n_4030),
.A2(n_3590),
.B(n_3486),
.Y(n_4342)
);

INVx1_ASAP7_75t_SL g4343 ( 
.A(n_4235),
.Y(n_4343)
);

INVxp67_ASAP7_75t_SL g4344 ( 
.A(n_3746),
.Y(n_4344)
);

OAI22xp5_ASAP7_75t_L g4345 ( 
.A1(n_4281),
.A2(n_3369),
.B1(n_3338),
.B2(n_3105),
.Y(n_4345)
);

AOI21xp5_ASAP7_75t_L g4346 ( 
.A1(n_4150),
.A2(n_3482),
.B(n_3473),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_3718),
.Y(n_4347)
);

AND2x2_ASAP7_75t_L g4348 ( 
.A(n_4246),
.B(n_3292),
.Y(n_4348)
);

NOR2xp33_ASAP7_75t_L g4349 ( 
.A(n_3815),
.B(n_3710),
.Y(n_4349)
);

NOR2xp33_ASAP7_75t_R g4350 ( 
.A(n_3858),
.B(n_3274),
.Y(n_4350)
);

AOI21xp5_ASAP7_75t_L g4351 ( 
.A1(n_3938),
.A2(n_3050),
.B(n_3460),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_4105),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_3750),
.Y(n_4353)
);

AND2x4_ASAP7_75t_SL g4354 ( 
.A(n_3794),
.B(n_3898),
.Y(n_4354)
);

BUFx6f_ASAP7_75t_L g4355 ( 
.A(n_3723),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_3751),
.Y(n_4356)
);

AND2x4_ASAP7_75t_L g4357 ( 
.A(n_3898),
.B(n_4214),
.Y(n_4357)
);

NAND2xp5_ASAP7_75t_SL g4358 ( 
.A(n_4254),
.B(n_3475),
.Y(n_4358)
);

OR2x2_ASAP7_75t_L g4359 ( 
.A(n_3802),
.B(n_3060),
.Y(n_4359)
);

NOR2xp33_ASAP7_75t_L g4360 ( 
.A(n_4191),
.B(n_3408),
.Y(n_4360)
);

AOI21xp5_ASAP7_75t_L g4361 ( 
.A1(n_4007),
.A2(n_3485),
.B(n_3484),
.Y(n_4361)
);

AND2x2_ASAP7_75t_L g4362 ( 
.A(n_4036),
.B(n_3292),
.Y(n_4362)
);

AOI21xp5_ASAP7_75t_L g4363 ( 
.A1(n_4016),
.A2(n_3182),
.B(n_3406),
.Y(n_4363)
);

AND2x2_ASAP7_75t_L g4364 ( 
.A(n_4188),
.B(n_3398),
.Y(n_4364)
);

BUFx2_ASAP7_75t_L g4365 ( 
.A(n_4017),
.Y(n_4365)
);

AOI22xp33_ASAP7_75t_L g4366 ( 
.A1(n_4284),
.A2(n_3293),
.B1(n_3318),
.B2(n_3304),
.Y(n_4366)
);

NAND2xp5_ASAP7_75t_SL g4367 ( 
.A(n_4254),
.B(n_3924),
.Y(n_4367)
);

OAI21xp33_ASAP7_75t_L g4368 ( 
.A1(n_3742),
.A2(n_3307),
.B(n_3303),
.Y(n_4368)
);

INVx2_ASAP7_75t_SL g4369 ( 
.A(n_4213),
.Y(n_4369)
);

AND2x2_ASAP7_75t_L g4370 ( 
.A(n_4197),
.B(n_4089),
.Y(n_4370)
);

NOR3xp33_ASAP7_75t_SL g4371 ( 
.A(n_3788),
.B(n_3822),
.C(n_3818),
.Y(n_4371)
);

BUFx2_ASAP7_75t_L g4372 ( 
.A(n_4017),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_3771),
.Y(n_4373)
);

A2O1A1Ixp33_ASAP7_75t_SL g4374 ( 
.A1(n_3904),
.A2(n_3121),
.B(n_3466),
.C(n_3458),
.Y(n_4374)
);

NAND2xp5_ASAP7_75t_SL g4375 ( 
.A(n_3924),
.B(n_3617),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_3796),
.Y(n_4376)
);

NAND2xp5_ASAP7_75t_L g4377 ( 
.A(n_4167),
.B(n_3131),
.Y(n_4377)
);

CKINVDCx5p33_ASAP7_75t_R g4378 ( 
.A(n_3768),
.Y(n_4378)
);

NAND2xp5_ASAP7_75t_L g4379 ( 
.A(n_4193),
.B(n_3162),
.Y(n_4379)
);

NOR2xp33_ASAP7_75t_R g4380 ( 
.A(n_3768),
.B(n_3408),
.Y(n_4380)
);

AOI21x1_ASAP7_75t_L g4381 ( 
.A1(n_4151),
.A2(n_3042),
.B(n_3137),
.Y(n_4381)
);

NOR2xp33_ASAP7_75t_L g4382 ( 
.A(n_4209),
.B(n_3282),
.Y(n_4382)
);

AOI21xp5_ASAP7_75t_L g4383 ( 
.A1(n_4049),
.A2(n_3148),
.B(n_3146),
.Y(n_4383)
);

INVx2_ASAP7_75t_L g4384 ( 
.A(n_3731),
.Y(n_4384)
);

NOR2xp33_ASAP7_75t_R g4385 ( 
.A(n_4059),
.B(n_3293),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_3798),
.Y(n_4386)
);

NAND2xp5_ASAP7_75t_L g4387 ( 
.A(n_4272),
.B(n_3178),
.Y(n_4387)
);

INVx3_ASAP7_75t_L g4388 ( 
.A(n_4214),
.Y(n_4388)
);

INVx2_ASAP7_75t_L g4389 ( 
.A(n_3732),
.Y(n_4389)
);

CKINVDCx5p33_ASAP7_75t_R g4390 ( 
.A(n_3918),
.Y(n_4390)
);

AOI21xp5_ASAP7_75t_L g4391 ( 
.A1(n_4083),
.A2(n_3394),
.B(n_3374),
.Y(n_4391)
);

A2O1A1Ixp33_ASAP7_75t_L g4392 ( 
.A1(n_4028),
.A2(n_3395),
.B(n_3324),
.C(n_3372),
.Y(n_4392)
);

AOI21xp5_ASAP7_75t_L g4393 ( 
.A1(n_4100),
.A2(n_3244),
.B(n_3216),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_3813),
.Y(n_4394)
);

NAND2xp5_ASAP7_75t_SL g4395 ( 
.A(n_3982),
.B(n_3111),
.Y(n_4395)
);

BUFx3_ASAP7_75t_L g4396 ( 
.A(n_3927),
.Y(n_4396)
);

BUFx6f_ASAP7_75t_L g4397 ( 
.A(n_3752),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_3839),
.Y(n_4398)
);

AO22x1_ASAP7_75t_L g4399 ( 
.A1(n_3806),
.A2(n_3411),
.B1(n_3168),
.B2(n_3461),
.Y(n_4399)
);

NAND2xp5_ASAP7_75t_L g4400 ( 
.A(n_3859),
.B(n_3179),
.Y(n_4400)
);

AND2x2_ASAP7_75t_L g4401 ( 
.A(n_4091),
.B(n_3127),
.Y(n_4401)
);

OR2x6_ASAP7_75t_L g4402 ( 
.A(n_3784),
.B(n_3361),
.Y(n_4402)
);

NOR2xp33_ASAP7_75t_R g4403 ( 
.A(n_3927),
.B(n_3183),
.Y(n_4403)
);

NAND2xp5_ASAP7_75t_SL g4404 ( 
.A(n_3982),
.B(n_3267),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_3868),
.Y(n_4405)
);

O2A1O1Ixp5_ASAP7_75t_SL g4406 ( 
.A1(n_3797),
.A2(n_3202),
.B(n_3262),
.C(n_3362),
.Y(n_4406)
);

AND2x2_ASAP7_75t_L g4407 ( 
.A(n_3811),
.B(n_3289),
.Y(n_4407)
);

OAI22xp5_ASAP7_75t_L g4408 ( 
.A1(n_3919),
.A2(n_3306),
.B1(n_514),
.B2(n_515),
.Y(n_4408)
);

AOI21xp5_ASAP7_75t_L g4409 ( 
.A1(n_4232),
.A2(n_515),
.B(n_513),
.Y(n_4409)
);

AND2x2_ASAP7_75t_L g4410 ( 
.A(n_3833),
.B(n_1150),
.Y(n_4410)
);

AOI21xp5_ASAP7_75t_L g4411 ( 
.A1(n_3830),
.A2(n_516),
.B(n_515),
.Y(n_4411)
);

NOR2xp33_ASAP7_75t_L g4412 ( 
.A(n_3906),
.B(n_516),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_3885),
.Y(n_4413)
);

INVx2_ASAP7_75t_L g4414 ( 
.A(n_3737),
.Y(n_4414)
);

NOR2xp33_ASAP7_75t_L g4415 ( 
.A(n_3842),
.B(n_517),
.Y(n_4415)
);

NOR2x1_ASAP7_75t_L g4416 ( 
.A(n_4099),
.B(n_517),
.Y(n_4416)
);

AOI21xp5_ASAP7_75t_L g4417 ( 
.A1(n_3849),
.A2(n_518),
.B(n_517),
.Y(n_4417)
);

INVx4_ASAP7_75t_L g4418 ( 
.A(n_4233),
.Y(n_4418)
);

NOR2xp33_ASAP7_75t_L g4419 ( 
.A(n_4164),
.B(n_518),
.Y(n_4419)
);

INVx1_ASAP7_75t_SL g4420 ( 
.A(n_3984),
.Y(n_4420)
);

NAND2xp5_ASAP7_75t_L g4421 ( 
.A(n_3939),
.B(n_518),
.Y(n_4421)
);

OAI22xp5_ASAP7_75t_L g4422 ( 
.A1(n_3926),
.A2(n_520),
.B1(n_521),
.B2(n_519),
.Y(n_4422)
);

NAND2x1p5_ASAP7_75t_L g4423 ( 
.A(n_4233),
.B(n_524),
.Y(n_4423)
);

NOR2xp33_ASAP7_75t_R g4424 ( 
.A(n_3724),
.B(n_519),
.Y(n_4424)
);

A2O1A1Ixp33_ASAP7_75t_L g4425 ( 
.A1(n_3860),
.A2(n_521),
.B(n_522),
.C(n_520),
.Y(n_4425)
);

HB1xp67_ASAP7_75t_L g4426 ( 
.A(n_4128),
.Y(n_4426)
);

AOI22xp5_ASAP7_75t_L g4427 ( 
.A1(n_3910),
.A2(n_522),
.B1(n_523),
.B2(n_521),
.Y(n_4427)
);

OA21x2_ASAP7_75t_L g4428 ( 
.A1(n_4180),
.A2(n_523),
.B(n_522),
.Y(n_4428)
);

NAND2xp5_ASAP7_75t_L g4429 ( 
.A(n_3943),
.B(n_523),
.Y(n_4429)
);

AOI22xp5_ASAP7_75t_L g4430 ( 
.A1(n_4038),
.A2(n_526),
.B1(n_527),
.B2(n_525),
.Y(n_4430)
);

AND2x4_ASAP7_75t_L g4431 ( 
.A(n_3950),
.B(n_525),
.Y(n_4431)
);

INVx3_ASAP7_75t_L g4432 ( 
.A(n_3729),
.Y(n_4432)
);

NOR2xp33_ASAP7_75t_SL g4433 ( 
.A(n_4280),
.B(n_525),
.Y(n_4433)
);

NOR2xp33_ASAP7_75t_L g4434 ( 
.A(n_3934),
.B(n_527),
.Y(n_4434)
);

O2A1O1Ixp5_ASAP7_75t_L g4435 ( 
.A1(n_3978),
.A2(n_528),
.B(n_529),
.C(n_527),
.Y(n_4435)
);

NAND3xp33_ASAP7_75t_SL g4436 ( 
.A(n_3956),
.B(n_4095),
.C(n_3850),
.Y(n_4436)
);

AOI22xp5_ASAP7_75t_L g4437 ( 
.A1(n_3825),
.A2(n_529),
.B1(n_530),
.B2(n_528),
.Y(n_4437)
);

AOI21xp5_ASAP7_75t_L g4438 ( 
.A1(n_4046),
.A2(n_530),
.B(n_528),
.Y(n_4438)
);

AOI21xp5_ASAP7_75t_L g4439 ( 
.A1(n_3894),
.A2(n_532),
.B(n_531),
.Y(n_4439)
);

NOR2xp33_ASAP7_75t_SL g4440 ( 
.A(n_3814),
.B(n_531),
.Y(n_4440)
);

HB1xp67_ASAP7_75t_L g4441 ( 
.A(n_3748),
.Y(n_4441)
);

BUFx6f_ASAP7_75t_L g4442 ( 
.A(n_3752),
.Y(n_4442)
);

INVxp67_ASAP7_75t_L g4443 ( 
.A(n_3985),
.Y(n_4443)
);

INVx3_ASAP7_75t_L g4444 ( 
.A(n_3729),
.Y(n_4444)
);

NAND2xp5_ASAP7_75t_L g4445 ( 
.A(n_3954),
.B(n_531),
.Y(n_4445)
);

NAND2xp5_ASAP7_75t_L g4446 ( 
.A(n_3975),
.B(n_532),
.Y(n_4446)
);

NOR2xp33_ASAP7_75t_L g4447 ( 
.A(n_3865),
.B(n_4160),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_4000),
.Y(n_4448)
);

O2A1O1Ixp5_ASAP7_75t_SL g4449 ( 
.A1(n_4145),
.A2(n_533),
.B(n_534),
.C(n_532),
.Y(n_4449)
);

BUFx12f_ASAP7_75t_L g4450 ( 
.A(n_3806),
.Y(n_4450)
);

AOI21xp5_ASAP7_75t_L g4451 ( 
.A1(n_4179),
.A2(n_534),
.B(n_533),
.Y(n_4451)
);

AOI21xp5_ASAP7_75t_L g4452 ( 
.A1(n_4249),
.A2(n_4287),
.B(n_4278),
.Y(n_4452)
);

AND2x4_ASAP7_75t_L g4453 ( 
.A(n_4027),
.B(n_533),
.Y(n_4453)
);

INVx2_ASAP7_75t_L g4454 ( 
.A(n_3781),
.Y(n_4454)
);

AOI21xp5_ASAP7_75t_L g4455 ( 
.A1(n_3760),
.A2(n_535),
.B(n_534),
.Y(n_4455)
);

AOI21xp5_ASAP7_75t_L g4456 ( 
.A1(n_4183),
.A2(n_536),
.B(n_535),
.Y(n_4456)
);

A2O1A1Ixp33_ASAP7_75t_L g4457 ( 
.A1(n_3749),
.A2(n_537),
.B(n_538),
.C(n_536),
.Y(n_4457)
);

INVx1_ASAP7_75t_L g4458 ( 
.A(n_4062),
.Y(n_4458)
);

BUFx2_ASAP7_75t_L g4459 ( 
.A(n_4027),
.Y(n_4459)
);

AOI21xp5_ASAP7_75t_L g4460 ( 
.A1(n_4263),
.A2(n_538),
.B(n_536),
.Y(n_4460)
);

INVx1_ASAP7_75t_SL g4461 ( 
.A(n_4086),
.Y(n_4461)
);

INVxp67_ASAP7_75t_SL g4462 ( 
.A(n_3843),
.Y(n_4462)
);

INVx4_ASAP7_75t_L g4463 ( 
.A(n_4213),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_L g4464 ( 
.A(n_4074),
.B(n_538),
.Y(n_4464)
);

HB1xp67_ASAP7_75t_L g4465 ( 
.A(n_4014),
.Y(n_4465)
);

INVx1_ASAP7_75t_L g4466 ( 
.A(n_4133),
.Y(n_4466)
);

AOI21xp5_ASAP7_75t_L g4467 ( 
.A1(n_4119),
.A2(n_540),
.B(n_539),
.Y(n_4467)
);

INVxp67_ASAP7_75t_L g4468 ( 
.A(n_4102),
.Y(n_4468)
);

AOI21xp5_ASAP7_75t_L g4469 ( 
.A1(n_3726),
.A2(n_540),
.B(n_539),
.Y(n_4469)
);

BUFx3_ASAP7_75t_L g4470 ( 
.A(n_4157),
.Y(n_4470)
);

OAI22xp5_ASAP7_75t_L g4471 ( 
.A1(n_3962),
.A2(n_541),
.B1(n_542),
.B2(n_539),
.Y(n_4471)
);

INVx1_ASAP7_75t_L g4472 ( 
.A(n_4134),
.Y(n_4472)
);

AND2x2_ASAP7_75t_L g4473 ( 
.A(n_4009),
.B(n_4029),
.Y(n_4473)
);

INVx2_ASAP7_75t_L g4474 ( 
.A(n_3787),
.Y(n_4474)
);

NOR2xp33_ASAP7_75t_L g4475 ( 
.A(n_4002),
.B(n_541),
.Y(n_4475)
);

NAND2xp5_ASAP7_75t_L g4476 ( 
.A(n_4155),
.B(n_541),
.Y(n_4476)
);

BUFx2_ASAP7_75t_L g4477 ( 
.A(n_3733),
.Y(n_4477)
);

OAI22xp5_ASAP7_75t_L g4478 ( 
.A1(n_4103),
.A2(n_543),
.B1(n_544),
.B2(n_542),
.Y(n_4478)
);

OAI22xp5_ASAP7_75t_L g4479 ( 
.A1(n_4135),
.A2(n_544),
.B1(n_545),
.B2(n_543),
.Y(n_4479)
);

INVx2_ASAP7_75t_L g4480 ( 
.A(n_3804),
.Y(n_4480)
);

NOR2x1_ASAP7_75t_R g4481 ( 
.A(n_4205),
.B(n_545),
.Y(n_4481)
);

BUFx6f_ASAP7_75t_L g4482 ( 
.A(n_3752),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_3827),
.Y(n_4483)
);

INVx4_ASAP7_75t_L g4484 ( 
.A(n_4213),
.Y(n_4484)
);

AOI21xp5_ASAP7_75t_L g4485 ( 
.A1(n_3911),
.A2(n_3940),
.B(n_3929),
.Y(n_4485)
);

O2A1O1Ixp33_ASAP7_75t_L g4486 ( 
.A1(n_3829),
.A2(n_546),
.B(n_547),
.C(n_545),
.Y(n_4486)
);

NAND3xp33_ASAP7_75t_SL g4487 ( 
.A(n_4137),
.B(n_50),
.C(n_51),
.Y(n_4487)
);

BUFx6f_ASAP7_75t_L g4488 ( 
.A(n_3790),
.Y(n_4488)
);

OAI22xp5_ASAP7_75t_L g4489 ( 
.A1(n_3713),
.A2(n_547),
.B1(n_548),
.B2(n_546),
.Y(n_4489)
);

INVx2_ASAP7_75t_L g4490 ( 
.A(n_3831),
.Y(n_4490)
);

NOR3xp33_ASAP7_75t_SL g4491 ( 
.A(n_4279),
.B(n_1150),
.C(n_1149),
.Y(n_4491)
);

HB1xp67_ASAP7_75t_L g4492 ( 
.A(n_4218),
.Y(n_4492)
);

INVx1_ASAP7_75t_L g4493 ( 
.A(n_3961),
.Y(n_4493)
);

INVxp67_ASAP7_75t_SL g4494 ( 
.A(n_3790),
.Y(n_4494)
);

BUFx2_ASAP7_75t_SL g4495 ( 
.A(n_4221),
.Y(n_4495)
);

OAI22xp5_ASAP7_75t_L g4496 ( 
.A1(n_3890),
.A2(n_547),
.B1(n_548),
.B2(n_546),
.Y(n_4496)
);

O2A1O1Ixp33_ASAP7_75t_L g4497 ( 
.A1(n_4258),
.A2(n_549),
.B(n_550),
.C(n_548),
.Y(n_4497)
);

INVx2_ASAP7_75t_L g4498 ( 
.A(n_3856),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_SL g4499 ( 
.A(n_3933),
.B(n_549),
.Y(n_4499)
);

CKINVDCx5p33_ASAP7_75t_R g4500 ( 
.A(n_4245),
.Y(n_4500)
);

NOR2x1_ASAP7_75t_L g4501 ( 
.A(n_4256),
.B(n_549),
.Y(n_4501)
);

OAI22xp5_ASAP7_75t_L g4502 ( 
.A1(n_4117),
.A2(n_551),
.B1(n_552),
.B2(n_550),
.Y(n_4502)
);

O2A1O1Ixp33_ASAP7_75t_L g4503 ( 
.A1(n_3869),
.A2(n_551),
.B(n_552),
.C(n_550),
.Y(n_4503)
);

OAI22xp5_ASAP7_75t_L g4504 ( 
.A1(n_4075),
.A2(n_552),
.B1(n_553),
.B2(n_551),
.Y(n_4504)
);

BUFx6f_ASAP7_75t_SL g4505 ( 
.A(n_3977),
.Y(n_4505)
);

NOR3xp33_ASAP7_75t_L g4506 ( 
.A(n_3872),
.B(n_554),
.C(n_553),
.Y(n_4506)
);

AOI21xp5_ASAP7_75t_L g4507 ( 
.A1(n_3941),
.A2(n_554),
.B(n_553),
.Y(n_4507)
);

OAI21xp33_ASAP7_75t_L g4508 ( 
.A1(n_4239),
.A2(n_4243),
.B(n_4148),
.Y(n_4508)
);

AOI21xp5_ASAP7_75t_L g4509 ( 
.A1(n_3942),
.A2(n_557),
.B(n_554),
.Y(n_4509)
);

INVx1_ASAP7_75t_SL g4510 ( 
.A(n_3912),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_L g4511 ( 
.A(n_4230),
.B(n_557),
.Y(n_4511)
);

NOR2xp67_ASAP7_75t_L g4512 ( 
.A(n_3733),
.B(n_557),
.Y(n_4512)
);

NOR2xp33_ASAP7_75t_L g4513 ( 
.A(n_3807),
.B(n_558),
.Y(n_4513)
);

BUFx6f_ASAP7_75t_L g4514 ( 
.A(n_3790),
.Y(n_4514)
);

A2O1A1Ixp33_ASAP7_75t_SL g4515 ( 
.A1(n_4268),
.A2(n_52),
.B(n_50),
.C(n_51),
.Y(n_4515)
);

AND2x4_ASAP7_75t_L g4516 ( 
.A(n_3968),
.B(n_558),
.Y(n_4516)
);

NAND2xp5_ASAP7_75t_SL g4517 ( 
.A(n_4051),
.B(n_558),
.Y(n_4517)
);

NAND2xp5_ASAP7_75t_L g4518 ( 
.A(n_3993),
.B(n_559),
.Y(n_4518)
);

O2A1O1Ixp33_ASAP7_75t_L g4519 ( 
.A1(n_3776),
.A2(n_561),
.B(n_562),
.C(n_560),
.Y(n_4519)
);

AOI21xp33_ASAP7_75t_L g4520 ( 
.A1(n_4067),
.A2(n_561),
.B(n_560),
.Y(n_4520)
);

AOI22xp33_ASAP7_75t_L g4521 ( 
.A1(n_3817),
.A2(n_562),
.B1(n_563),
.B2(n_561),
.Y(n_4521)
);

AND2x2_ASAP7_75t_L g4522 ( 
.A(n_3960),
.B(n_4081),
.Y(n_4522)
);

HB1xp67_ASAP7_75t_L g4523 ( 
.A(n_4177),
.Y(n_4523)
);

NOR2xp33_ASAP7_75t_L g4524 ( 
.A(n_3824),
.B(n_563),
.Y(n_4524)
);

BUFx8_ASAP7_75t_L g4525 ( 
.A(n_4221),
.Y(n_4525)
);

INVx4_ASAP7_75t_L g4526 ( 
.A(n_4221),
.Y(n_4526)
);

INVx1_ASAP7_75t_L g4527 ( 
.A(n_3971),
.Y(n_4527)
);

NAND2xp5_ASAP7_75t_L g4528 ( 
.A(n_3711),
.B(n_565),
.Y(n_4528)
);

A2O1A1Ixp33_ASAP7_75t_L g4529 ( 
.A1(n_3758),
.A2(n_566),
.B(n_567),
.C(n_565),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_SL g4530 ( 
.A(n_4051),
.B(n_565),
.Y(n_4530)
);

AND2x2_ASAP7_75t_L g4531 ( 
.A(n_4053),
.B(n_1151),
.Y(n_4531)
);

NOR2xp33_ASAP7_75t_L g4532 ( 
.A(n_3952),
.B(n_3874),
.Y(n_4532)
);

INVx1_ASAP7_75t_L g4533 ( 
.A(n_3979),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_SL g4534 ( 
.A(n_4051),
.B(n_566),
.Y(n_4534)
);

INVx2_ASAP7_75t_L g4535 ( 
.A(n_3875),
.Y(n_4535)
);

AOI21xp5_ASAP7_75t_L g4536 ( 
.A1(n_3946),
.A2(n_567),
.B(n_566),
.Y(n_4536)
);

AOI21xp5_ASAP7_75t_L g4537 ( 
.A1(n_3948),
.A2(n_569),
.B(n_568),
.Y(n_4537)
);

O2A1O1Ixp33_ASAP7_75t_L g4538 ( 
.A1(n_4210),
.A2(n_569),
.B(n_570),
.C(n_568),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_L g4539 ( 
.A(n_4175),
.B(n_568),
.Y(n_4539)
);

NAND2xp5_ASAP7_75t_SL g4540 ( 
.A(n_4041),
.B(n_570),
.Y(n_4540)
);

NOR3xp33_ASAP7_75t_L g4541 ( 
.A(n_3887),
.B(n_571),
.C(n_570),
.Y(n_4541)
);

HB1xp67_ASAP7_75t_L g4542 ( 
.A(n_4177),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_SL g4543 ( 
.A(n_4041),
.B(n_572),
.Y(n_4543)
);

OAI22xp33_ASAP7_75t_L g4544 ( 
.A1(n_3944),
.A2(n_573),
.B1(n_574),
.B2(n_572),
.Y(n_4544)
);

OAI21xp33_ASAP7_75t_SL g4545 ( 
.A1(n_3855),
.A2(n_573),
.B(n_572),
.Y(n_4545)
);

INVx1_ASAP7_75t_L g4546 ( 
.A(n_3983),
.Y(n_4546)
);

OAI21xp5_ASAP7_75t_L g4547 ( 
.A1(n_3779),
.A2(n_575),
.B(n_574),
.Y(n_4547)
);

O2A1O1Ixp5_ASAP7_75t_SL g4548 ( 
.A1(n_4153),
.A2(n_575),
.B(n_576),
.C(n_574),
.Y(n_4548)
);

INVx2_ASAP7_75t_L g4549 ( 
.A(n_3914),
.Y(n_4549)
);

AND2x2_ASAP7_75t_L g4550 ( 
.A(n_3735),
.B(n_1162),
.Y(n_4550)
);

NOR2xp33_ASAP7_75t_R g4551 ( 
.A(n_3739),
.B(n_575),
.Y(n_4551)
);

NAND2xp5_ASAP7_75t_L g4552 ( 
.A(n_4208),
.B(n_576),
.Y(n_4552)
);

INVxp67_ASAP7_75t_L g4553 ( 
.A(n_4122),
.Y(n_4553)
);

NAND2xp5_ASAP7_75t_SL g4554 ( 
.A(n_4058),
.B(n_577),
.Y(n_4554)
);

OAI22xp5_ASAP7_75t_L g4555 ( 
.A1(n_3932),
.A2(n_578),
.B1(n_579),
.B2(n_577),
.Y(n_4555)
);

INVx4_ASAP7_75t_L g4556 ( 
.A(n_4229),
.Y(n_4556)
);

O2A1O1Ixp5_ASAP7_75t_L g4557 ( 
.A1(n_3789),
.A2(n_578),
.B(n_579),
.C(n_577),
.Y(n_4557)
);

NAND2xp5_ASAP7_75t_L g4558 ( 
.A(n_3990),
.B(n_578),
.Y(n_4558)
);

AOI21xp5_ASAP7_75t_L g4559 ( 
.A1(n_3959),
.A2(n_581),
.B(n_580),
.Y(n_4559)
);

NAND2xp5_ASAP7_75t_L g4560 ( 
.A(n_4034),
.B(n_4200),
.Y(n_4560)
);

AND2x2_ASAP7_75t_L g4561 ( 
.A(n_4170),
.B(n_4094),
.Y(n_4561)
);

BUFx6f_ASAP7_75t_L g4562 ( 
.A(n_3799),
.Y(n_4562)
);

INVx2_ASAP7_75t_L g4563 ( 
.A(n_3951),
.Y(n_4563)
);

INVx3_ASAP7_75t_L g4564 ( 
.A(n_3739),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_4271),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_SL g4566 ( 
.A(n_4058),
.B(n_580),
.Y(n_4566)
);

HB1xp67_ASAP7_75t_L g4567 ( 
.A(n_4290),
.Y(n_4567)
);

A2O1A1Ixp33_ASAP7_75t_SL g4568 ( 
.A1(n_4273),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_4568)
);

NAND2xp5_ASAP7_75t_SL g4569 ( 
.A(n_3963),
.B(n_580),
.Y(n_4569)
);

NOR2xp33_ASAP7_75t_SL g4570 ( 
.A(n_3883),
.B(n_581),
.Y(n_4570)
);

AOI21xp5_ASAP7_75t_L g4571 ( 
.A1(n_3964),
.A2(n_583),
.B(n_582),
.Y(n_4571)
);

AOI21xp5_ASAP7_75t_L g4572 ( 
.A1(n_3974),
.A2(n_583),
.B(n_582),
.Y(n_4572)
);

AOI21xp5_ASAP7_75t_L g4573 ( 
.A1(n_3976),
.A2(n_583),
.B(n_582),
.Y(n_4573)
);

A2O1A1Ixp33_ASAP7_75t_L g4574 ( 
.A1(n_3759),
.A2(n_585),
.B(n_586),
.C(n_584),
.Y(n_4574)
);

INVxp67_ASAP7_75t_L g4575 ( 
.A(n_4290),
.Y(n_4575)
);

OAI22xp5_ASAP7_75t_L g4576 ( 
.A1(n_3892),
.A2(n_585),
.B1(n_586),
.B2(n_584),
.Y(n_4576)
);

NAND2xp5_ASAP7_75t_L g4577 ( 
.A(n_4003),
.B(n_584),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_4090),
.Y(n_4578)
);

INVx4_ASAP7_75t_L g4579 ( 
.A(n_4229),
.Y(n_4579)
);

CKINVDCx8_ASAP7_75t_R g4580 ( 
.A(n_4229),
.Y(n_4580)
);

OAI22xp5_ASAP7_75t_SL g4581 ( 
.A1(n_4259),
.A2(n_586),
.B1(n_587),
.B2(n_585),
.Y(n_4581)
);

NOR2xp33_ASAP7_75t_L g4582 ( 
.A(n_3891),
.B(n_587),
.Y(n_4582)
);

INVx3_ASAP7_75t_L g4583 ( 
.A(n_3883),
.Y(n_4583)
);

NAND2xp5_ASAP7_75t_L g4584 ( 
.A(n_4114),
.B(n_588),
.Y(n_4584)
);

OR2x6_ASAP7_75t_L g4585 ( 
.A(n_3801),
.B(n_588),
.Y(n_4585)
);

INVx3_ASAP7_75t_L g4586 ( 
.A(n_4098),
.Y(n_4586)
);

AO22x1_ASAP7_75t_L g4587 ( 
.A1(n_3740),
.A2(n_589),
.B1(n_590),
.B2(n_588),
.Y(n_4587)
);

OAI22xp5_ASAP7_75t_L g4588 ( 
.A1(n_4154),
.A2(n_590),
.B1(n_591),
.B2(n_589),
.Y(n_4588)
);

INVx2_ASAP7_75t_L g4589 ( 
.A(n_4120),
.Y(n_4589)
);

NAND2xp5_ASAP7_75t_L g4590 ( 
.A(n_3712),
.B(n_589),
.Y(n_4590)
);

AOI21xp5_ASAP7_75t_L g4591 ( 
.A1(n_3981),
.A2(n_591),
.B(n_590),
.Y(n_4591)
);

BUFx8_ASAP7_75t_L g4592 ( 
.A(n_4248),
.Y(n_4592)
);

INVx1_ASAP7_75t_L g4593 ( 
.A(n_3953),
.Y(n_4593)
);

CKINVDCx5p33_ASAP7_75t_R g4594 ( 
.A(n_3716),
.Y(n_4594)
);

NAND2xp5_ASAP7_75t_L g4595 ( 
.A(n_3809),
.B(n_591),
.Y(n_4595)
);

INVx1_ASAP7_75t_L g4596 ( 
.A(n_3957),
.Y(n_4596)
);

AOI21xp5_ASAP7_75t_L g4597 ( 
.A1(n_3992),
.A2(n_593),
.B(n_592),
.Y(n_4597)
);

INVx1_ASAP7_75t_L g4598 ( 
.A(n_3820),
.Y(n_4598)
);

NAND2xp5_ASAP7_75t_L g4599 ( 
.A(n_4136),
.B(n_593),
.Y(n_4599)
);

AOI22xp5_ASAP7_75t_L g4600 ( 
.A1(n_3901),
.A2(n_595),
.B1(n_596),
.B2(n_594),
.Y(n_4600)
);

AOI21xp5_ASAP7_75t_L g4601 ( 
.A1(n_3995),
.A2(n_596),
.B(n_594),
.Y(n_4601)
);

BUFx6f_ASAP7_75t_L g4602 ( 
.A(n_3799),
.Y(n_4602)
);

BUFx4f_ASAP7_75t_L g4603 ( 
.A(n_3740),
.Y(n_4603)
);

A2O1A1Ixp33_ASAP7_75t_L g4604 ( 
.A1(n_4234),
.A2(n_596),
.B(n_597),
.C(n_594),
.Y(n_4604)
);

INVx2_ASAP7_75t_L g4605 ( 
.A(n_4192),
.Y(n_4605)
);

NAND2xp5_ASAP7_75t_SL g4606 ( 
.A(n_3799),
.B(n_597),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_3821),
.Y(n_4607)
);

AOI21xp5_ASAP7_75t_L g4608 ( 
.A1(n_3996),
.A2(n_598),
.B(n_597),
.Y(n_4608)
);

AOI22xp5_ASAP7_75t_L g4609 ( 
.A1(n_3917),
.A2(n_599),
.B1(n_600),
.B2(n_598),
.Y(n_4609)
);

AND2x2_ASAP7_75t_L g4610 ( 
.A(n_4216),
.B(n_1152),
.Y(n_4610)
);

NAND2xp5_ASAP7_75t_L g4611 ( 
.A(n_4261),
.B(n_598),
.Y(n_4611)
);

AOI21xp5_ASAP7_75t_L g4612 ( 
.A1(n_3997),
.A2(n_600),
.B(n_599),
.Y(n_4612)
);

BUFx6f_ASAP7_75t_L g4613 ( 
.A(n_3853),
.Y(n_4613)
);

BUFx2_ASAP7_75t_L g4614 ( 
.A(n_3912),
.Y(n_4614)
);

A2O1A1Ixp33_ASAP7_75t_L g4615 ( 
.A1(n_4060),
.A2(n_600),
.B(n_601),
.C(n_599),
.Y(n_4615)
);

AOI21xp5_ASAP7_75t_L g4616 ( 
.A1(n_4010),
.A2(n_602),
.B(n_601),
.Y(n_4616)
);

NAND2xp5_ASAP7_75t_L g4617 ( 
.A(n_4118),
.B(n_601),
.Y(n_4617)
);

NAND2xp5_ASAP7_75t_L g4618 ( 
.A(n_3958),
.B(n_3878),
.Y(n_4618)
);

INVx2_ASAP7_75t_L g4619 ( 
.A(n_4225),
.Y(n_4619)
);

NAND2xp5_ASAP7_75t_L g4620 ( 
.A(n_3786),
.B(n_602),
.Y(n_4620)
);

BUFx12f_ASAP7_75t_L g4621 ( 
.A(n_3720),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_3826),
.Y(n_4622)
);

NAND2xp5_ASAP7_75t_L g4623 ( 
.A(n_3792),
.B(n_602),
.Y(n_4623)
);

NAND2xp5_ASAP7_75t_L g4624 ( 
.A(n_3803),
.B(n_603),
.Y(n_4624)
);

BUFx6f_ASAP7_75t_L g4625 ( 
.A(n_3853),
.Y(n_4625)
);

AOI21xp5_ASAP7_75t_L g4626 ( 
.A1(n_4018),
.A2(n_4042),
.B(n_4031),
.Y(n_4626)
);

BUFx6f_ASAP7_75t_L g4627 ( 
.A(n_3853),
.Y(n_4627)
);

AOI21xp5_ASAP7_75t_L g4628 ( 
.A1(n_4043),
.A2(n_604),
.B(n_603),
.Y(n_4628)
);

AOI21xp5_ASAP7_75t_L g4629 ( 
.A1(n_4047),
.A2(n_604),
.B(n_603),
.Y(n_4629)
);

NAND2xp5_ASAP7_75t_L g4630 ( 
.A(n_4202),
.B(n_604),
.Y(n_4630)
);

NAND2xp5_ASAP7_75t_L g4631 ( 
.A(n_4181),
.B(n_605),
.Y(n_4631)
);

NOR2xp33_ASAP7_75t_L g4632 ( 
.A(n_3900),
.B(n_605),
.Y(n_4632)
);

O2A1O1Ixp5_ASAP7_75t_L g4633 ( 
.A1(n_3836),
.A2(n_607),
.B(n_608),
.C(n_606),
.Y(n_4633)
);

AND2x2_ASAP7_75t_L g4634 ( 
.A(n_3913),
.B(n_1161),
.Y(n_4634)
);

BUFx3_ASAP7_75t_L g4635 ( 
.A(n_4098),
.Y(n_4635)
);

AND2x2_ASAP7_75t_L g4636 ( 
.A(n_3913),
.B(n_3720),
.Y(n_4636)
);

OAI22xp5_ASAP7_75t_L g4637 ( 
.A1(n_4250),
.A2(n_607),
.B1(n_608),
.B2(n_606),
.Y(n_4637)
);

INVx2_ASAP7_75t_L g4638 ( 
.A(n_3873),
.Y(n_4638)
);

NOR2xp33_ASAP7_75t_R g4639 ( 
.A(n_3740),
.B(n_606),
.Y(n_4639)
);

OAI22xp5_ASAP7_75t_L g4640 ( 
.A1(n_4265),
.A2(n_608),
.B1(n_609),
.B2(n_607),
.Y(n_4640)
);

OAI22xp5_ASAP7_75t_L g4641 ( 
.A1(n_4267),
.A2(n_610),
.B1(n_611),
.B2(n_609),
.Y(n_4641)
);

NAND2xp5_ASAP7_75t_L g4642 ( 
.A(n_4285),
.B(n_609),
.Y(n_4642)
);

XOR2xp5_ASAP7_75t_L g4643 ( 
.A(n_3972),
.B(n_51),
.Y(n_4643)
);

NOR2xp33_ASAP7_75t_L g4644 ( 
.A(n_3907),
.B(n_610),
.Y(n_4644)
);

AOI21xp5_ASAP7_75t_L g4645 ( 
.A1(n_4055),
.A2(n_611),
.B(n_610),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_4186),
.B(n_612),
.Y(n_4646)
);

BUFx2_ASAP7_75t_L g4647 ( 
.A(n_3740),
.Y(n_4647)
);

O2A1O1Ixp33_ASAP7_75t_L g4648 ( 
.A1(n_3851),
.A2(n_613),
.B(n_614),
.C(n_612),
.Y(n_4648)
);

HB1xp67_ASAP7_75t_L g4649 ( 
.A(n_3902),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_4189),
.B(n_613),
.Y(n_4650)
);

NOR2xp33_ASAP7_75t_L g4651 ( 
.A(n_3753),
.B(n_613),
.Y(n_4651)
);

BUFx6f_ASAP7_75t_L g4652 ( 
.A(n_3861),
.Y(n_4652)
);

NOR2xp33_ASAP7_75t_L g4653 ( 
.A(n_3947),
.B(n_614),
.Y(n_4653)
);

NOR2xp33_ASAP7_75t_L g4654 ( 
.A(n_3773),
.B(n_614),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_3828),
.Y(n_4655)
);

BUFx2_ASAP7_75t_L g4656 ( 
.A(n_4098),
.Y(n_4656)
);

O2A1O1Ixp33_ASAP7_75t_L g4657 ( 
.A1(n_3903),
.A2(n_616),
.B(n_617),
.C(n_615),
.Y(n_4657)
);

O2A1O1Ixp33_ASAP7_75t_L g4658 ( 
.A1(n_4065),
.A2(n_4068),
.B(n_4071),
.C(n_4066),
.Y(n_4658)
);

CKINVDCx5p33_ASAP7_75t_R g4659 ( 
.A(n_4132),
.Y(n_4659)
);

NOR2x1_ASAP7_75t_L g4660 ( 
.A(n_4172),
.B(n_615),
.Y(n_4660)
);

AOI21xp5_ASAP7_75t_L g4661 ( 
.A1(n_4056),
.A2(n_4076),
.B(n_4064),
.Y(n_4661)
);

BUFx3_ASAP7_75t_L g4662 ( 
.A(n_4132),
.Y(n_4662)
);

OAI22xp5_ASAP7_75t_L g4663 ( 
.A1(n_3905),
.A2(n_616),
.B1(n_617),
.B2(n_615),
.Y(n_4663)
);

BUFx2_ASAP7_75t_L g4664 ( 
.A(n_4132),
.Y(n_4664)
);

OR2x6_ASAP7_75t_L g4665 ( 
.A(n_4184),
.B(n_617),
.Y(n_4665)
);

AND2x2_ASAP7_75t_SL g4666 ( 
.A(n_4184),
.B(n_618),
.Y(n_4666)
);

AOI22xp5_ASAP7_75t_L g4667 ( 
.A1(n_4286),
.A2(n_620),
.B1(n_621),
.B2(n_618),
.Y(n_4667)
);

BUFx3_ASAP7_75t_L g4668 ( 
.A(n_4184),
.Y(n_4668)
);

AOI21x1_ASAP7_75t_L g4669 ( 
.A1(n_3989),
.A2(n_620),
.B(n_618),
.Y(n_4669)
);

O2A1O1Ixp33_ASAP7_75t_L g4670 ( 
.A1(n_4124),
.A2(n_621),
.B(n_622),
.C(n_620),
.Y(n_4670)
);

BUFx6f_ASAP7_75t_L g4671 ( 
.A(n_3861),
.Y(n_4671)
);

CKINVDCx5p33_ASAP7_75t_R g4672 ( 
.A(n_3785),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_3837),
.Y(n_4673)
);

NOR2xp33_ASAP7_75t_L g4674 ( 
.A(n_4139),
.B(n_621),
.Y(n_4674)
);

AO21x1_ASAP7_75t_L g4675 ( 
.A1(n_4008),
.A2(n_624),
.B(n_623),
.Y(n_4675)
);

OAI22xp5_ASAP7_75t_L g4676 ( 
.A1(n_4063),
.A2(n_624),
.B1(n_625),
.B2(n_623),
.Y(n_4676)
);

CKINVDCx5p33_ASAP7_75t_R g4677 ( 
.A(n_3715),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_3838),
.Y(n_4678)
);

INVx2_ASAP7_75t_SL g4679 ( 
.A(n_4264),
.Y(n_4679)
);

AOI21xp5_ASAP7_75t_L g4680 ( 
.A1(n_4080),
.A2(n_624),
.B(n_623),
.Y(n_4680)
);

AOI21xp5_ASAP7_75t_L g4681 ( 
.A1(n_4082),
.A2(n_627),
.B(n_626),
.Y(n_4681)
);

NAND2xp5_ASAP7_75t_L g4682 ( 
.A(n_4292),
.B(n_626),
.Y(n_4682)
);

AOI21xp5_ASAP7_75t_L g4683 ( 
.A1(n_4087),
.A2(n_627),
.B(n_626),
.Y(n_4683)
);

AOI21xp5_ASAP7_75t_L g4684 ( 
.A1(n_4088),
.A2(n_629),
.B(n_628),
.Y(n_4684)
);

O2A1O1Ixp33_ASAP7_75t_L g4685 ( 
.A1(n_4242),
.A2(n_630),
.B(n_631),
.C(n_628),
.Y(n_4685)
);

INVx4_ASAP7_75t_L g4686 ( 
.A(n_4264),
.Y(n_4686)
);

A2O1A1Ixp33_ASAP7_75t_L g4687 ( 
.A1(n_4026),
.A2(n_631),
.B(n_632),
.C(n_630),
.Y(n_4687)
);

NAND3xp33_ASAP7_75t_L g4688 ( 
.A(n_4173),
.B(n_1155),
.C(n_1153),
.Y(n_4688)
);

INVxp33_ASAP7_75t_SL g4689 ( 
.A(n_4024),
.Y(n_4689)
);

NAND2xp5_ASAP7_75t_SL g4690 ( 
.A(n_3861),
.B(n_4032),
.Y(n_4690)
);

INVx2_ASAP7_75t_L g4691 ( 
.A(n_3999),
.Y(n_4691)
);

AOI21xp5_ASAP7_75t_L g4692 ( 
.A1(n_4096),
.A2(n_632),
.B(n_630),
.Y(n_4692)
);

BUFx10_ASAP7_75t_L g4693 ( 
.A(n_3876),
.Y(n_4693)
);

OAI22xp5_ASAP7_75t_L g4694 ( 
.A1(n_4040),
.A2(n_634),
.B1(n_635),
.B2(n_633),
.Y(n_4694)
);

NAND2xp5_ASAP7_75t_L g4695 ( 
.A(n_4131),
.B(n_633),
.Y(n_4695)
);

NOR2xp33_ASAP7_75t_L g4696 ( 
.A(n_4282),
.B(n_4275),
.Y(n_4696)
);

OAI21xp33_ASAP7_75t_L g4697 ( 
.A1(n_4020),
.A2(n_52),
.B(n_53),
.Y(n_4697)
);

OA21x2_ASAP7_75t_L g4698 ( 
.A1(n_3896),
.A2(n_636),
.B(n_634),
.Y(n_4698)
);

OAI22xp5_ASAP7_75t_L g4699 ( 
.A1(n_4226),
.A2(n_636),
.B1(n_637),
.B2(n_634),
.Y(n_4699)
);

NAND2xp5_ASAP7_75t_L g4700 ( 
.A(n_4252),
.B(n_636),
.Y(n_4700)
);

O2A1O1Ixp33_ASAP7_75t_L g4701 ( 
.A1(n_4044),
.A2(n_638),
.B(n_640),
.C(n_637),
.Y(n_4701)
);

NAND2xp5_ASAP7_75t_L g4702 ( 
.A(n_4138),
.B(n_638),
.Y(n_4702)
);

NOR2xp33_ASAP7_75t_R g4703 ( 
.A(n_3902),
.B(n_640),
.Y(n_4703)
);

INVx5_ASAP7_75t_L g4704 ( 
.A(n_3876),
.Y(n_4704)
);

INVx1_ASAP7_75t_L g4705 ( 
.A(n_3844),
.Y(n_4705)
);

AOI21xp5_ASAP7_75t_L g4706 ( 
.A1(n_4101),
.A2(n_642),
.B(n_641),
.Y(n_4706)
);

NAND2xp5_ASAP7_75t_L g4707 ( 
.A(n_4140),
.B(n_641),
.Y(n_4707)
);

INVx4_ASAP7_75t_L g4708 ( 
.A(n_4264),
.Y(n_4708)
);

INVx2_ASAP7_75t_L g4709 ( 
.A(n_4054),
.Y(n_4709)
);

BUFx3_ASAP7_75t_L g4710 ( 
.A(n_3908),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_SL g4711 ( 
.A(n_3876),
.B(n_641),
.Y(n_4711)
);

AOI21xp5_ASAP7_75t_L g4712 ( 
.A1(n_4107),
.A2(n_643),
.B(n_642),
.Y(n_4712)
);

NAND2xp5_ASAP7_75t_L g4713 ( 
.A(n_4142),
.B(n_642),
.Y(n_4713)
);

OAI21xp33_ASAP7_75t_SL g4714 ( 
.A1(n_4070),
.A2(n_644),
.B(n_643),
.Y(n_4714)
);

O2A1O1Ixp33_ASAP7_75t_L g4715 ( 
.A1(n_3719),
.A2(n_644),
.B(n_645),
.C(n_643),
.Y(n_4715)
);

BUFx6f_ASAP7_75t_L g4716 ( 
.A(n_3970),
.Y(n_4716)
);

NAND2xp5_ASAP7_75t_L g4717 ( 
.A(n_4149),
.B(n_645),
.Y(n_4717)
);

O2A1O1Ixp33_ASAP7_75t_L g4718 ( 
.A1(n_3897),
.A2(n_646),
.B(n_647),
.C(n_645),
.Y(n_4718)
);

OAI22xp5_ASAP7_75t_L g4719 ( 
.A1(n_4006),
.A2(n_647),
.B1(n_648),
.B2(n_646),
.Y(n_4719)
);

NOR2x1_ASAP7_75t_L g4720 ( 
.A(n_4079),
.B(n_646),
.Y(n_4720)
);

AOI21xp33_ASAP7_75t_L g4721 ( 
.A1(n_4110),
.A2(n_650),
.B(n_649),
.Y(n_4721)
);

BUFx6f_ASAP7_75t_L g4722 ( 
.A(n_3970),
.Y(n_4722)
);

O2A1O1Ixp33_ASAP7_75t_L g4723 ( 
.A1(n_4215),
.A2(n_651),
.B(n_652),
.C(n_650),
.Y(n_4723)
);

NOR2xp67_ASAP7_75t_L g4724 ( 
.A(n_4061),
.B(n_651),
.Y(n_4724)
);

AOI21xp5_ASAP7_75t_L g4725 ( 
.A1(n_4111),
.A2(n_652),
.B(n_651),
.Y(n_4725)
);

CKINVDCx5p33_ASAP7_75t_R g4726 ( 
.A(n_3782),
.Y(n_4726)
);

AND2x2_ASAP7_75t_L g4727 ( 
.A(n_3808),
.B(n_1158),
.Y(n_4727)
);

NAND2xp5_ASAP7_75t_L g4728 ( 
.A(n_4156),
.B(n_652),
.Y(n_4728)
);

NAND2xp5_ASAP7_75t_SL g4729 ( 
.A(n_3970),
.B(n_653),
.Y(n_4729)
);

AOI21xp5_ASAP7_75t_L g4730 ( 
.A1(n_4112),
.A2(n_654),
.B(n_653),
.Y(n_4730)
);

AOI21xp5_ASAP7_75t_L g4731 ( 
.A1(n_4019),
.A2(n_654),
.B(n_653),
.Y(n_4731)
);

NAND2xp5_ASAP7_75t_L g4732 ( 
.A(n_4162),
.B(n_654),
.Y(n_4732)
);

OR2x2_ASAP7_75t_L g4733 ( 
.A(n_3727),
.B(n_655),
.Y(n_4733)
);

AOI21xp5_ASAP7_75t_L g4734 ( 
.A1(n_3780),
.A2(n_656),
.B(n_655),
.Y(n_4734)
);

AOI21xp5_ASAP7_75t_L g4735 ( 
.A1(n_3763),
.A2(n_656),
.B(n_655),
.Y(n_4735)
);

A2O1A1Ixp33_ASAP7_75t_L g4736 ( 
.A1(n_4078),
.A2(n_657),
.B(n_658),
.C(n_656),
.Y(n_4736)
);

O2A1O1Ixp33_ASAP7_75t_L g4737 ( 
.A1(n_4217),
.A2(n_658),
.B(n_659),
.C(n_657),
.Y(n_4737)
);

A2O1A1Ixp33_ASAP7_75t_SL g4738 ( 
.A1(n_4052),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_4738)
);

INVx2_ASAP7_75t_L g4739 ( 
.A(n_4092),
.Y(n_4739)
);

INVx2_ASAP7_75t_L g4740 ( 
.A(n_4032),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_3847),
.Y(n_4741)
);

CKINVDCx20_ASAP7_75t_R g4742 ( 
.A(n_4032),
.Y(n_4742)
);

NAND2xp5_ASAP7_75t_SL g4743 ( 
.A(n_3908),
.B(n_658),
.Y(n_4743)
);

NAND2xp5_ASAP7_75t_L g4744 ( 
.A(n_4166),
.B(n_659),
.Y(n_4744)
);

NOR2xp33_ASAP7_75t_SL g4745 ( 
.A(n_3777),
.B(n_4206),
.Y(n_4745)
);

AOI22xp33_ASAP7_75t_SL g4746 ( 
.A1(n_4277),
.A2(n_660),
.B1(n_661),
.B2(n_659),
.Y(n_4746)
);

INVx5_ASAP7_75t_L g4747 ( 
.A(n_3922),
.Y(n_4747)
);

INVx2_ASAP7_75t_L g4748 ( 
.A(n_4244),
.Y(n_4748)
);

NOR3xp33_ASAP7_75t_SL g4749 ( 
.A(n_4269),
.B(n_4171),
.C(n_4169),
.Y(n_4749)
);

OAI21xp5_ASAP7_75t_L g4750 ( 
.A1(n_4174),
.A2(n_661),
.B(n_660),
.Y(n_4750)
);

O2A1O1Ixp33_ASAP7_75t_L g4751 ( 
.A1(n_4222),
.A2(n_663),
.B(n_664),
.C(n_662),
.Y(n_4751)
);

CKINVDCx5p33_ASAP7_75t_R g4752 ( 
.A(n_4288),
.Y(n_4752)
);

A2O1A1Ixp33_ASAP7_75t_L g4753 ( 
.A1(n_3741),
.A2(n_663),
.B(n_664),
.C(n_662),
.Y(n_4753)
);

A2O1A1Ixp33_ASAP7_75t_L g4754 ( 
.A1(n_3764),
.A2(n_663),
.B(n_665),
.C(n_662),
.Y(n_4754)
);

O2A1O1Ixp33_ASAP7_75t_L g4755 ( 
.A1(n_4223),
.A2(n_666),
.B(n_667),
.C(n_665),
.Y(n_4755)
);

AOI21xp5_ASAP7_75t_L g4756 ( 
.A1(n_4228),
.A2(n_666),
.B(n_665),
.Y(n_4756)
);

NAND2xp5_ASAP7_75t_L g4757 ( 
.A(n_3734),
.B(n_667),
.Y(n_4757)
);

HB1xp67_ASAP7_75t_L g4758 ( 
.A(n_3922),
.Y(n_4758)
);

NAND2xp5_ASAP7_75t_L g4759 ( 
.A(n_3744),
.B(n_667),
.Y(n_4759)
);

NAND3xp33_ASAP7_75t_L g4760 ( 
.A(n_3819),
.B(n_1164),
.C(n_1162),
.Y(n_4760)
);

INVx2_ASAP7_75t_SL g4761 ( 
.A(n_4224),
.Y(n_4761)
);

BUFx8_ASAP7_75t_L g4762 ( 
.A(n_4288),
.Y(n_4762)
);

AND2x2_ASAP7_75t_L g4763 ( 
.A(n_3754),
.B(n_1162),
.Y(n_4763)
);

AOI21xp5_ASAP7_75t_L g4764 ( 
.A1(n_3769),
.A2(n_669),
.B(n_668),
.Y(n_4764)
);

NAND2x1p5_ASAP7_75t_L g4765 ( 
.A(n_3925),
.B(n_669),
.Y(n_4765)
);

AOI21xp5_ASAP7_75t_L g4766 ( 
.A1(n_3775),
.A2(n_669),
.B(n_668),
.Y(n_4766)
);

O2A1O1Ixp5_ASAP7_75t_L g4767 ( 
.A1(n_3840),
.A2(n_670),
.B(n_671),
.C(n_668),
.Y(n_4767)
);

CKINVDCx6p67_ASAP7_75t_R g4768 ( 
.A(n_3986),
.Y(n_4768)
);

NAND2xp5_ASAP7_75t_L g4769 ( 
.A(n_3757),
.B(n_670),
.Y(n_4769)
);

AOI21xp5_ASAP7_75t_L g4770 ( 
.A1(n_3791),
.A2(n_673),
.B(n_672),
.Y(n_4770)
);

INVx2_ASAP7_75t_L g4771 ( 
.A(n_4257),
.Y(n_4771)
);

NAND2xp5_ASAP7_75t_L g4772 ( 
.A(n_3762),
.B(n_672),
.Y(n_4772)
);

INVx2_ASAP7_75t_SL g4773 ( 
.A(n_4224),
.Y(n_4773)
);

AOI21xp5_ASAP7_75t_L g4774 ( 
.A1(n_3793),
.A2(n_674),
.B(n_672),
.Y(n_4774)
);

BUFx4f_ASAP7_75t_L g4775 ( 
.A(n_4288),
.Y(n_4775)
);

BUFx3_ASAP7_75t_L g4776 ( 
.A(n_3925),
.Y(n_4776)
);

INVxp67_ASAP7_75t_L g4777 ( 
.A(n_4084),
.Y(n_4777)
);

OAI21xp33_ASAP7_75t_L g4778 ( 
.A1(n_3881),
.A2(n_54),
.B(n_55),
.Y(n_4778)
);

HB1xp67_ASAP7_75t_L g4779 ( 
.A(n_3867),
.Y(n_4779)
);

AOI21xp5_ASAP7_75t_L g4780 ( 
.A1(n_3795),
.A2(n_676),
.B(n_675),
.Y(n_4780)
);

OAI22x1_ASAP7_75t_L g4781 ( 
.A1(n_3991),
.A2(n_4045),
.B1(n_4011),
.B2(n_3864),
.Y(n_4781)
);

AOI22xp5_ASAP7_75t_L g4782 ( 
.A1(n_3857),
.A2(n_676),
.B1(n_677),
.B2(n_675),
.Y(n_4782)
);

A2O1A1Ixp33_ASAP7_75t_L g4783 ( 
.A1(n_3832),
.A2(n_677),
.B(n_679),
.C(n_675),
.Y(n_4783)
);

OAI22xp5_ASAP7_75t_L g4784 ( 
.A1(n_3880),
.A2(n_679),
.B1(n_680),
.B2(n_677),
.Y(n_4784)
);

NOR2xp33_ASAP7_75t_L g4785 ( 
.A(n_3765),
.B(n_680),
.Y(n_4785)
);

AND2x6_ASAP7_75t_L g4786 ( 
.A(n_4291),
.B(n_683),
.Y(n_4786)
);

AOI21xp33_ASAP7_75t_L g4787 ( 
.A1(n_3783),
.A2(n_682),
.B(n_681),
.Y(n_4787)
);

AOI22xp33_ASAP7_75t_L g4788 ( 
.A1(n_3921),
.A2(n_682),
.B1(n_683),
.B2(n_681),
.Y(n_4788)
);

NAND2xp5_ASAP7_75t_L g4789 ( 
.A(n_4238),
.B(n_681),
.Y(n_4789)
);

NOR2xp33_ASAP7_75t_L g4790 ( 
.A(n_4163),
.B(n_683),
.Y(n_4790)
);

A2O1A1Ixp33_ASAP7_75t_L g4791 ( 
.A1(n_3899),
.A2(n_685),
.B(n_686),
.C(n_684),
.Y(n_4791)
);

AOI21xp5_ASAP7_75t_L g4792 ( 
.A1(n_3945),
.A2(n_685),
.B(n_684),
.Y(n_4792)
);

O2A1O1Ixp33_ASAP7_75t_L g4793 ( 
.A1(n_3862),
.A2(n_686),
.B(n_687),
.C(n_685),
.Y(n_4793)
);

OA21x2_ASAP7_75t_L g4794 ( 
.A1(n_4129),
.A2(n_687),
.B(n_686),
.Y(n_4794)
);

AOI21xp5_ASAP7_75t_L g4795 ( 
.A1(n_3955),
.A2(n_689),
.B(n_688),
.Y(n_4795)
);

AOI221xp5_ASAP7_75t_L g4796 ( 
.A1(n_4147),
.A2(n_690),
.B1(n_691),
.B2(n_689),
.C(n_688),
.Y(n_4796)
);

AO22x1_ASAP7_75t_L g4797 ( 
.A1(n_4283),
.A2(n_690),
.B1(n_691),
.B2(n_688),
.Y(n_4797)
);

AND2x2_ASAP7_75t_L g4798 ( 
.A(n_4251),
.B(n_1149),
.Y(n_4798)
);

AOI21xp5_ASAP7_75t_L g4799 ( 
.A1(n_4185),
.A2(n_693),
.B(n_691),
.Y(n_4799)
);

AOI22xp5_ASAP7_75t_L g4800 ( 
.A1(n_4190),
.A2(n_694),
.B1(n_695),
.B2(n_693),
.Y(n_4800)
);

AOI22xp33_ASAP7_75t_L g4801 ( 
.A1(n_4012),
.A2(n_695),
.B1(n_696),
.B2(n_694),
.Y(n_4801)
);

BUFx6f_ASAP7_75t_L g4802 ( 
.A(n_4291),
.Y(n_4802)
);

NOR3xp33_ASAP7_75t_SL g4803 ( 
.A(n_4207),
.B(n_1155),
.C(n_1153),
.Y(n_4803)
);

A2O1A1Ixp33_ASAP7_75t_L g4804 ( 
.A1(n_4113),
.A2(n_695),
.B(n_696),
.C(n_694),
.Y(n_4804)
);

AOI22xp33_ASAP7_75t_L g4805 ( 
.A1(n_4126),
.A2(n_698),
.B1(n_699),
.B2(n_697),
.Y(n_4805)
);

AOI21xp5_ASAP7_75t_L g4806 ( 
.A1(n_4130),
.A2(n_698),
.B(n_697),
.Y(n_4806)
);

INVx1_ASAP7_75t_L g4807 ( 
.A(n_3870),
.Y(n_4807)
);

BUFx6f_ASAP7_75t_L g4808 ( 
.A(n_4196),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_3877),
.Y(n_4809)
);

INVx1_ASAP7_75t_L g4810 ( 
.A(n_3879),
.Y(n_4810)
);

NAND2xp5_ASAP7_75t_L g4811 ( 
.A(n_3884),
.B(n_697),
.Y(n_4811)
);

INVx2_ASAP7_75t_L g4812 ( 
.A(n_3886),
.Y(n_4812)
);

NAND2xp5_ASAP7_75t_L g4813 ( 
.A(n_3888),
.B(n_699),
.Y(n_4813)
);

INVx1_ASAP7_75t_L g4814 ( 
.A(n_4198),
.Y(n_4814)
);

BUFx6f_ASAP7_75t_L g4815 ( 
.A(n_4035),
.Y(n_4815)
);

NAND2xp5_ASAP7_75t_L g4816 ( 
.A(n_4270),
.B(n_699),
.Y(n_4816)
);

CKINVDCx5p33_ASAP7_75t_R g4817 ( 
.A(n_4293),
.Y(n_4817)
);

A2O1A1Ixp33_ASAP7_75t_L g4818 ( 
.A1(n_4085),
.A2(n_701),
.B(n_702),
.C(n_700),
.Y(n_4818)
);

INVxp67_ASAP7_75t_SL g4819 ( 
.A(n_4276),
.Y(n_4819)
);

INVx2_ASAP7_75t_L g4820 ( 
.A(n_4187),
.Y(n_4820)
);

OR2x2_ASAP7_75t_L g4821 ( 
.A(n_3772),
.B(n_700),
.Y(n_4821)
);

O2A1O1Ixp33_ASAP7_75t_L g4822 ( 
.A1(n_3969),
.A2(n_701),
.B(n_702),
.C(n_700),
.Y(n_4822)
);

OAI22xp5_ASAP7_75t_L g4823 ( 
.A1(n_4253),
.A2(n_702),
.B1(n_703),
.B2(n_701),
.Y(n_4823)
);

AO21x1_ASAP7_75t_L g4824 ( 
.A1(n_3714),
.A2(n_704),
.B(n_703),
.Y(n_4824)
);

NOR2x1_ASAP7_75t_L g4825 ( 
.A(n_3738),
.B(n_704),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_3965),
.Y(n_4826)
);

AOI21xp5_ASAP7_75t_L g4827 ( 
.A1(n_3722),
.A2(n_705),
.B(n_704),
.Y(n_4827)
);

NOR2xp33_ASAP7_75t_L g4828 ( 
.A(n_4199),
.B(n_4201),
.Y(n_4828)
);

OAI22xp5_ASAP7_75t_L g4829 ( 
.A1(n_4021),
.A2(n_706),
.B1(n_707),
.B2(n_705),
.Y(n_4829)
);

NAND2xp5_ASAP7_75t_L g4830 ( 
.A(n_4203),
.B(n_706),
.Y(n_4830)
);

INVx1_ASAP7_75t_L g4831 ( 
.A(n_3747),
.Y(n_4831)
);

AOI221xp5_ASAP7_75t_L g4832 ( 
.A1(n_4204),
.A2(n_4159),
.B1(n_4161),
.B2(n_4158),
.C(n_4152),
.Y(n_4832)
);

O2A1O1Ixp33_ASAP7_75t_L g4833 ( 
.A1(n_3936),
.A2(n_707),
.B(n_708),
.C(n_706),
.Y(n_4833)
);

INVx1_ASAP7_75t_L g4834 ( 
.A(n_3800),
.Y(n_4834)
);

INVx5_ASAP7_75t_L g4835 ( 
.A(n_3730),
.Y(n_4835)
);

AOI21xp5_ASAP7_75t_L g4836 ( 
.A1(n_3935),
.A2(n_709),
.B(n_708),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_L g4837 ( 
.A(n_4165),
.B(n_708),
.Y(n_4837)
);

AND2x4_ASAP7_75t_L g4838 ( 
.A(n_4182),
.B(n_709),
.Y(n_4838)
);

NOR2xp33_ASAP7_75t_L g4839 ( 
.A(n_4194),
.B(n_709),
.Y(n_4839)
);

BUFx2_ASAP7_75t_L g4840 ( 
.A(n_4057),
.Y(n_4840)
);

BUFx2_ASAP7_75t_L g4841 ( 
.A(n_4219),
.Y(n_4841)
);

NAND2x1p5_ASAP7_75t_L g4842 ( 
.A(n_4220),
.B(n_712),
.Y(n_4842)
);

NOR2xp33_ASAP7_75t_L g4843 ( 
.A(n_4195),
.B(n_710),
.Y(n_4843)
);

NOR2x1_ASAP7_75t_L g4844 ( 
.A(n_4211),
.B(n_710),
.Y(n_4844)
);

NAND2xp5_ASAP7_75t_L g4845 ( 
.A(n_4241),
.B(n_710),
.Y(n_4845)
);

AOI21xp5_ASAP7_75t_L g4846 ( 
.A1(n_3743),
.A2(n_712),
.B(n_711),
.Y(n_4846)
);

NOR2x1_ASAP7_75t_SL g4847 ( 
.A(n_4231),
.B(n_1155),
.Y(n_4847)
);

AOI21xp5_ASAP7_75t_L g4848 ( 
.A1(n_3967),
.A2(n_712),
.B(n_711),
.Y(n_4848)
);

NOR2xp33_ASAP7_75t_L g4849 ( 
.A(n_4247),
.B(n_713),
.Y(n_4849)
);

A2O1A1Ixp33_ASAP7_75t_L g4850 ( 
.A1(n_4072),
.A2(n_4097),
.B(n_4108),
.C(n_4093),
.Y(n_4850)
);

CKINVDCx20_ASAP7_75t_R g4851 ( 
.A(n_4255),
.Y(n_4851)
);

AOI21xp5_ASAP7_75t_L g4852 ( 
.A1(n_3973),
.A2(n_715),
.B(n_714),
.Y(n_4852)
);

NOR2xp33_ASAP7_75t_L g4853 ( 
.A(n_4260),
.B(n_714),
.Y(n_4853)
);

AOI21xp5_ASAP7_75t_L g4854 ( 
.A1(n_3987),
.A2(n_716),
.B(n_715),
.Y(n_4854)
);

AOI22xp5_ASAP7_75t_L g4855 ( 
.A1(n_4262),
.A2(n_716),
.B1(n_717),
.B2(n_715),
.Y(n_4855)
);

INVx1_ASAP7_75t_L g4856 ( 
.A(n_3805),
.Y(n_4856)
);

AOI22xp5_ASAP7_75t_L g4857 ( 
.A1(n_4240),
.A2(n_717),
.B1(n_718),
.B2(n_716),
.Y(n_4857)
);

NAND2xp5_ASAP7_75t_SL g4858 ( 
.A(n_3812),
.B(n_718),
.Y(n_4858)
);

NOR2xp33_ASAP7_75t_L g4859 ( 
.A(n_3949),
.B(n_718),
.Y(n_4859)
);

OAI22xp5_ASAP7_75t_L g4860 ( 
.A1(n_3816),
.A2(n_3823),
.B1(n_3841),
.B2(n_3835),
.Y(n_4860)
);

NAND2xp5_ASAP7_75t_SL g4861 ( 
.A(n_3846),
.B(n_719),
.Y(n_4861)
);

AND2x4_ASAP7_75t_L g4862 ( 
.A(n_3988),
.B(n_720),
.Y(n_4862)
);

NAND2xp5_ASAP7_75t_L g4863 ( 
.A(n_3848),
.B(n_720),
.Y(n_4863)
);

AOI22xp33_ASAP7_75t_L g4864 ( 
.A1(n_3774),
.A2(n_721),
.B1(n_722),
.B2(n_720),
.Y(n_4864)
);

INVx1_ASAP7_75t_L g4865 ( 
.A(n_3863),
.Y(n_4865)
);

AO32x2_ASAP7_75t_L g4866 ( 
.A1(n_3866),
.A2(n_723),
.A3(n_724),
.B1(n_722),
.B2(n_721),
.Y(n_4866)
);

AND2x2_ASAP7_75t_L g4867 ( 
.A(n_4306),
.B(n_721),
.Y(n_4867)
);

INVx3_ASAP7_75t_L g4868 ( 
.A(n_4354),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4300),
.Y(n_4869)
);

A2O1A1Ixp33_ASAP7_75t_L g4870 ( 
.A1(n_4603),
.A2(n_4327),
.B(n_4724),
.C(n_4508),
.Y(n_4870)
);

OAI21x1_ASAP7_75t_L g4871 ( 
.A1(n_4323),
.A2(n_4015),
.B(n_4001),
.Y(n_4871)
);

O2A1O1Ixp5_ASAP7_75t_SL g4872 ( 
.A1(n_4310),
.A2(n_723),
.B(n_724),
.C(n_722),
.Y(n_4872)
);

OAI21x1_ASAP7_75t_L g4873 ( 
.A1(n_4342),
.A2(n_4004),
.B(n_3998),
.Y(n_4873)
);

AOI22xp5_ASAP7_75t_L g4874 ( 
.A1(n_4689),
.A2(n_4048),
.B1(n_3923),
.B2(n_3882),
.Y(n_4874)
);

BUFx6f_ASAP7_75t_L g4875 ( 
.A(n_4580),
.Y(n_4875)
);

AOI221x1_ASAP7_75t_L g4876 ( 
.A1(n_4294),
.A2(n_4037),
.B1(n_4039),
.B2(n_4033),
.C(n_4023),
.Y(n_4876)
);

O2A1O1Ixp5_ASAP7_75t_L g4877 ( 
.A1(n_4316),
.A2(n_3889),
.B(n_3893),
.C(n_3871),
.Y(n_4877)
);

BUFx12f_ASAP7_75t_L g4878 ( 
.A(n_4450),
.Y(n_4878)
);

OAI21x1_ASAP7_75t_L g4879 ( 
.A1(n_4748),
.A2(n_4013),
.B(n_4005),
.Y(n_4879)
);

AOI21xp5_ASAP7_75t_L g4880 ( 
.A1(n_4297),
.A2(n_3916),
.B(n_3909),
.Y(n_4880)
);

INVx4_ASAP7_75t_L g4881 ( 
.A(n_4301),
.Y(n_4881)
);

INVx3_ASAP7_75t_L g4882 ( 
.A(n_4418),
.Y(n_4882)
);

OAI21xp5_ASAP7_75t_L g4883 ( 
.A1(n_4557),
.A2(n_3928),
.B(n_3920),
.Y(n_4883)
);

AOI221xp5_ASAP7_75t_L g4884 ( 
.A1(n_4696),
.A2(n_4069),
.B1(n_4050),
.B2(n_4289),
.C(n_4274),
.Y(n_4884)
);

OA22x2_ASAP7_75t_L g4885 ( 
.A1(n_4585),
.A2(n_724),
.B1(n_725),
.B2(n_723),
.Y(n_4885)
);

NAND2xp5_ASAP7_75t_L g4886 ( 
.A(n_4483),
.B(n_725),
.Y(n_4886)
);

CKINVDCx6p67_ASAP7_75t_R g4887 ( 
.A(n_4396),
.Y(n_4887)
);

AOI21xp5_ASAP7_75t_L g4888 ( 
.A1(n_4302),
.A2(n_4123),
.B(n_4109),
.Y(n_4888)
);

AOI21xp5_ASAP7_75t_L g4889 ( 
.A1(n_4690),
.A2(n_4116),
.B(n_4125),
.Y(n_4889)
);

AOI221x1_ASAP7_75t_L g4890 ( 
.A1(n_4778),
.A2(n_727),
.B1(n_728),
.B2(n_726),
.C(n_725),
.Y(n_4890)
);

BUFx6f_ASAP7_75t_L g4891 ( 
.A(n_4357),
.Y(n_4891)
);

BUFx6f_ASAP7_75t_L g4892 ( 
.A(n_4470),
.Y(n_4892)
);

NAND2xp5_ASAP7_75t_L g4893 ( 
.A(n_4473),
.B(n_726),
.Y(n_4893)
);

NAND2xp5_ASAP7_75t_L g4894 ( 
.A(n_4322),
.B(n_727),
.Y(n_4894)
);

BUFx6f_ASAP7_75t_L g4895 ( 
.A(n_4301),
.Y(n_4895)
);

OAI22xp5_ASAP7_75t_L g4896 ( 
.A1(n_4677),
.A2(n_729),
.B1(n_730),
.B2(n_728),
.Y(n_4896)
);

NAND2xp5_ASAP7_75t_L g4897 ( 
.A(n_4370),
.B(n_728),
.Y(n_4897)
);

AOI21xp5_ASAP7_75t_L g4898 ( 
.A1(n_4334),
.A2(n_4314),
.B(n_4452),
.Y(n_4898)
);

NAND2x1p5_ASAP7_75t_L g4899 ( 
.A(n_4301),
.B(n_729),
.Y(n_4899)
);

CKINVDCx5p33_ASAP7_75t_R g4900 ( 
.A(n_4350),
.Y(n_4900)
);

NAND2xp5_ASAP7_75t_L g4901 ( 
.A(n_4303),
.B(n_730),
.Y(n_4901)
);

OAI21xp33_ASAP7_75t_SL g4902 ( 
.A1(n_4666),
.A2(n_731),
.B(n_730),
.Y(n_4902)
);

NAND3x1_ASAP7_75t_L g4903 ( 
.A(n_4320),
.B(n_732),
.C(n_731),
.Y(n_4903)
);

AOI21xp5_ASAP7_75t_L g4904 ( 
.A1(n_4346),
.A2(n_732),
.B(n_731),
.Y(n_4904)
);

NOR3xp33_ASAP7_75t_L g4905 ( 
.A(n_4333),
.B(n_743),
.C(n_735),
.Y(n_4905)
);

NAND2xp5_ASAP7_75t_SL g4906 ( 
.A(n_4639),
.B(n_733),
.Y(n_4906)
);

AOI21x1_ASAP7_75t_L g4907 ( 
.A1(n_4771),
.A2(n_734),
.B(n_733),
.Y(n_4907)
);

AOI22xp5_ASAP7_75t_L g4908 ( 
.A1(n_4349),
.A2(n_1144),
.B1(n_1145),
.B2(n_1143),
.Y(n_4908)
);

NOR2xp33_ASAP7_75t_L g4909 ( 
.A(n_4315),
.B(n_734),
.Y(n_4909)
);

NAND2xp5_ASAP7_75t_L g4910 ( 
.A(n_4312),
.B(n_4321),
.Y(n_4910)
);

INVx4_ASAP7_75t_L g4911 ( 
.A(n_4338),
.Y(n_4911)
);

OAI21xp5_ASAP7_75t_L g4912 ( 
.A1(n_4767),
.A2(n_736),
.B(n_735),
.Y(n_4912)
);

OAI21xp5_ASAP7_75t_L g4913 ( 
.A1(n_4688),
.A2(n_738),
.B(n_737),
.Y(n_4913)
);

BUFx3_ASAP7_75t_L g4914 ( 
.A(n_4525),
.Y(n_4914)
);

NOR2xp67_ASAP7_75t_SL g4915 ( 
.A(n_4621),
.B(n_737),
.Y(n_4915)
);

AND2x4_ASAP7_75t_L g4916 ( 
.A(n_4463),
.B(n_737),
.Y(n_4916)
);

O2A1O1Ixp33_ASAP7_75t_L g4917 ( 
.A1(n_4392),
.A2(n_740),
.B(n_741),
.C(n_739),
.Y(n_4917)
);

AO21x1_ASAP7_75t_L g4918 ( 
.A1(n_4570),
.A2(n_740),
.B(n_739),
.Y(n_4918)
);

INVx1_ASAP7_75t_L g4919 ( 
.A(n_4352),
.Y(n_4919)
);

AOI21xp5_ASAP7_75t_SL g4920 ( 
.A1(n_4665),
.A2(n_741),
.B(n_740),
.Y(n_4920)
);

INVx1_ASAP7_75t_L g4921 ( 
.A(n_4353),
.Y(n_4921)
);

AOI221x1_ASAP7_75t_L g4922 ( 
.A1(n_4456),
.A2(n_4436),
.B1(n_4697),
.B2(n_4781),
.C(n_4532),
.Y(n_4922)
);

OAI21xp5_ASAP7_75t_SL g4923 ( 
.A1(n_4487),
.A2(n_1156),
.B(n_1153),
.Y(n_4923)
);

AOI21xp5_ASAP7_75t_L g4924 ( 
.A1(n_4485),
.A2(n_743),
.B(n_742),
.Y(n_4924)
);

BUFx6f_ASAP7_75t_L g4925 ( 
.A(n_4317),
.Y(n_4925)
);

INVx1_ASAP7_75t_L g4926 ( 
.A(n_4356),
.Y(n_4926)
);

OR2x6_ASAP7_75t_L g4927 ( 
.A(n_4399),
.B(n_743),
.Y(n_4927)
);

AND2x2_ASAP7_75t_L g4928 ( 
.A(n_4522),
.B(n_744),
.Y(n_4928)
);

CKINVDCx20_ASAP7_75t_R g4929 ( 
.A(n_4390),
.Y(n_4929)
);

NOR2xp33_ASAP7_75t_L g4930 ( 
.A(n_4440),
.B(n_744),
.Y(n_4930)
);

AOI221x1_ASAP7_75t_L g4931 ( 
.A1(n_4626),
.A2(n_747),
.B1(n_748),
.B2(n_746),
.C(n_745),
.Y(n_4931)
);

OA21x2_ASAP7_75t_L g4932 ( 
.A1(n_4691),
.A2(n_746),
.B(n_745),
.Y(n_4932)
);

NAND2xp5_ASAP7_75t_L g4933 ( 
.A(n_4373),
.B(n_746),
.Y(n_4933)
);

OAI22x1_ASAP7_75t_L g4934 ( 
.A1(n_4643),
.A2(n_748),
.B1(n_749),
.B2(n_747),
.Y(n_4934)
);

NOR2xp67_ASAP7_75t_L g4935 ( 
.A(n_4388),
.B(n_750),
.Y(n_4935)
);

NAND2xp5_ASAP7_75t_L g4936 ( 
.A(n_4376),
.B(n_747),
.Y(n_4936)
);

INVx5_ASAP7_75t_L g4937 ( 
.A(n_4665),
.Y(n_4937)
);

OAI21x1_ASAP7_75t_L g4938 ( 
.A1(n_4638),
.A2(n_750),
.B(n_749),
.Y(n_4938)
);

BUFx6f_ASAP7_75t_L g4939 ( 
.A(n_4340),
.Y(n_4939)
);

BUFx6f_ASAP7_75t_L g4940 ( 
.A(n_4484),
.Y(n_4940)
);

OAI22x1_ASAP7_75t_L g4941 ( 
.A1(n_4462),
.A2(n_751),
.B1(n_752),
.B2(n_749),
.Y(n_4941)
);

OR2x2_ASAP7_75t_L g4942 ( 
.A(n_4339),
.B(n_751),
.Y(n_4942)
);

NOR2xp33_ASAP7_75t_L g4943 ( 
.A(n_4311),
.B(n_751),
.Y(n_4943)
);

OAI21x1_ASAP7_75t_L g4944 ( 
.A1(n_4709),
.A2(n_753),
.B(n_752),
.Y(n_4944)
);

NAND2x1_ASAP7_75t_L g4945 ( 
.A(n_4647),
.B(n_753),
.Y(n_4945)
);

NOR2xp33_ASAP7_75t_L g4946 ( 
.A(n_4481),
.B(n_753),
.Y(n_4946)
);

AND2x2_ASAP7_75t_L g4947 ( 
.A(n_4410),
.B(n_4561),
.Y(n_4947)
);

OA21x2_ASAP7_75t_L g4948 ( 
.A1(n_4739),
.A2(n_4865),
.B(n_4856),
.Y(n_4948)
);

NAND2xp5_ASAP7_75t_L g4949 ( 
.A(n_4386),
.B(n_754),
.Y(n_4949)
);

OAI21x1_ASAP7_75t_L g4950 ( 
.A1(n_4319),
.A2(n_755),
.B(n_754),
.Y(n_4950)
);

AOI21xp5_ASAP7_75t_L g4951 ( 
.A1(n_4661),
.A2(n_756),
.B(n_755),
.Y(n_4951)
);

BUFx3_ASAP7_75t_L g4952 ( 
.A(n_4304),
.Y(n_4952)
);

NAND2xp5_ASAP7_75t_L g4953 ( 
.A(n_4394),
.B(n_4398),
.Y(n_4953)
);

AOI22xp5_ASAP7_75t_L g4954 ( 
.A1(n_4324),
.A2(n_1152),
.B1(n_1157),
.B2(n_1150),
.Y(n_4954)
);

CKINVDCx11_ASAP7_75t_R g4955 ( 
.A(n_4402),
.Y(n_4955)
);

INVx1_ASAP7_75t_L g4956 ( 
.A(n_4405),
.Y(n_4956)
);

AOI21xp5_ASAP7_75t_L g4957 ( 
.A1(n_4860),
.A2(n_757),
.B(n_756),
.Y(n_4957)
);

O2A1O1Ixp33_ASAP7_75t_L g4958 ( 
.A1(n_4368),
.A2(n_4515),
.B(n_4308),
.C(n_4568),
.Y(n_4958)
);

BUFx12f_ASAP7_75t_L g4959 ( 
.A(n_4378),
.Y(n_4959)
);

OAI21x1_ASAP7_75t_L g4960 ( 
.A1(n_4831),
.A2(n_758),
.B(n_757),
.Y(n_4960)
);

OAI21x1_ASAP7_75t_L g4961 ( 
.A1(n_4834),
.A2(n_758),
.B(n_757),
.Y(n_4961)
);

NAND2xp5_ASAP7_75t_L g4962 ( 
.A(n_4413),
.B(n_759),
.Y(n_4962)
);

AOI221xp5_ASAP7_75t_L g4963 ( 
.A1(n_4785),
.A2(n_761),
.B1(n_762),
.B2(n_760),
.C(n_759),
.Y(n_4963)
);

A2O1A1Ixp33_ASAP7_75t_L g4964 ( 
.A1(n_4658),
.A2(n_760),
.B(n_761),
.C(n_759),
.Y(n_4964)
);

NOR4xp25_ASAP7_75t_L g4965 ( 
.A(n_4443),
.B(n_762),
.C(n_763),
.D(n_760),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4448),
.Y(n_4966)
);

NAND2xp5_ASAP7_75t_L g4967 ( 
.A(n_4458),
.B(n_762),
.Y(n_4967)
);

OAI21x1_ASAP7_75t_L g4968 ( 
.A1(n_4826),
.A2(n_764),
.B(n_763),
.Y(n_4968)
);

INVx2_ASAP7_75t_L g4969 ( 
.A(n_4347),
.Y(n_4969)
);

AND2x4_ASAP7_75t_L g4970 ( 
.A(n_4526),
.B(n_763),
.Y(n_4970)
);

NOR2xp33_ASAP7_75t_L g4971 ( 
.A(n_4298),
.B(n_4295),
.Y(n_4971)
);

NAND2xp5_ASAP7_75t_SL g4972 ( 
.A(n_4703),
.B(n_764),
.Y(n_4972)
);

OAI21xp33_ASAP7_75t_L g4973 ( 
.A1(n_4424),
.A2(n_766),
.B(n_765),
.Y(n_4973)
);

OR2x2_ASAP7_75t_L g4974 ( 
.A(n_4426),
.B(n_765),
.Y(n_4974)
);

INVx1_ASAP7_75t_L g4975 ( 
.A(n_4466),
.Y(n_4975)
);

OAI21xp5_ASAP7_75t_L g4976 ( 
.A1(n_4435),
.A2(n_766),
.B(n_765),
.Y(n_4976)
);

AOI21x1_ASAP7_75t_L g4977 ( 
.A1(n_4296),
.A2(n_767),
.B(n_766),
.Y(n_4977)
);

OAI21x1_ASAP7_75t_L g4978 ( 
.A1(n_4669),
.A2(n_768),
.B(n_767),
.Y(n_4978)
);

AOI21x1_ASAP7_75t_SL g4979 ( 
.A1(n_4539),
.A2(n_769),
.B(n_768),
.Y(n_4979)
);

NAND2xp5_ASAP7_75t_L g4980 ( 
.A(n_4472),
.B(n_768),
.Y(n_4980)
);

AOI21xp5_ASAP7_75t_SL g4981 ( 
.A1(n_4736),
.A2(n_770),
.B(n_769),
.Y(n_4981)
);

A2O1A1Ixp33_ASAP7_75t_L g4982 ( 
.A1(n_4803),
.A2(n_770),
.B(n_771),
.C(n_769),
.Y(n_4982)
);

AOI21xp5_ASAP7_75t_L g4983 ( 
.A1(n_4335),
.A2(n_771),
.B(n_770),
.Y(n_4983)
);

AO32x2_ASAP7_75t_L g4984 ( 
.A1(n_4581),
.A2(n_774),
.A3(n_775),
.B1(n_773),
.B2(n_772),
.Y(n_4984)
);

AND2x2_ASAP7_75t_L g4985 ( 
.A(n_4401),
.B(n_772),
.Y(n_4985)
);

OR2x2_ASAP7_75t_L g4986 ( 
.A(n_4465),
.B(n_772),
.Y(n_4986)
);

INVx1_ASAP7_75t_L g4987 ( 
.A(n_4493),
.Y(n_4987)
);

OAI21xp5_ASAP7_75t_L g4988 ( 
.A1(n_4633),
.A2(n_4307),
.B(n_4760),
.Y(n_4988)
);

NAND2xp5_ASAP7_75t_L g4989 ( 
.A(n_4527),
.B(n_773),
.Y(n_4989)
);

BUFx2_ASAP7_75t_L g4990 ( 
.A(n_4742),
.Y(n_4990)
);

NAND2xp5_ASAP7_75t_L g4991 ( 
.A(n_4533),
.B(n_773),
.Y(n_4991)
);

OAI21x1_ASAP7_75t_L g4992 ( 
.A1(n_4740),
.A2(n_775),
.B(n_774),
.Y(n_4992)
);

OA21x2_ASAP7_75t_L g4993 ( 
.A1(n_4841),
.A2(n_776),
.B(n_775),
.Y(n_4993)
);

AOI21xp5_ASAP7_75t_L g4994 ( 
.A1(n_4494),
.A2(n_777),
.B(n_776),
.Y(n_4994)
);

AOI21xp5_ASAP7_75t_L g4995 ( 
.A1(n_4828),
.A2(n_4351),
.B(n_4850),
.Y(n_4995)
);

NAND2xp5_ASAP7_75t_L g4996 ( 
.A(n_4546),
.B(n_776),
.Y(n_4996)
);

CKINVDCx20_ASAP7_75t_R g4997 ( 
.A(n_4403),
.Y(n_4997)
);

AOI221xp5_ASAP7_75t_SL g4998 ( 
.A1(n_4777),
.A2(n_57),
.B1(n_54),
.B2(n_56),
.C(n_58),
.Y(n_4998)
);

NAND2x1p5_ASAP7_75t_L g4999 ( 
.A(n_4556),
.B(n_777),
.Y(n_4999)
);

NAND2xp5_ASAP7_75t_SL g5000 ( 
.A(n_4385),
.B(n_777),
.Y(n_5000)
);

NAND2xp5_ASAP7_75t_L g5001 ( 
.A(n_4565),
.B(n_778),
.Y(n_5001)
);

INVx1_ASAP7_75t_L g5002 ( 
.A(n_4578),
.Y(n_5002)
);

HB1xp67_ASAP7_75t_L g5003 ( 
.A(n_4492),
.Y(n_5003)
);

OAI21xp5_ASAP7_75t_L g5004 ( 
.A1(n_4770),
.A2(n_4780),
.B(n_4774),
.Y(n_5004)
);

INVx2_ASAP7_75t_L g5005 ( 
.A(n_4384),
.Y(n_5005)
);

AND2x2_ASAP7_75t_L g5006 ( 
.A(n_4550),
.B(n_778),
.Y(n_5006)
);

NAND3xp33_ASAP7_75t_SL g5007 ( 
.A(n_4551),
.B(n_54),
.C(n_56),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4593),
.Y(n_5008)
);

AOI21xp5_ASAP7_75t_L g5009 ( 
.A1(n_4361),
.A2(n_779),
.B(n_778),
.Y(n_5009)
);

AOI21xp5_ASAP7_75t_L g5010 ( 
.A1(n_4840),
.A2(n_780),
.B(n_779),
.Y(n_5010)
);

NAND2xp5_ASAP7_75t_L g5011 ( 
.A(n_4598),
.B(n_779),
.Y(n_5011)
);

INVxp67_ASAP7_75t_L g5012 ( 
.A(n_4433),
.Y(n_5012)
);

AND2x2_ASAP7_75t_L g5013 ( 
.A(n_4362),
.B(n_780),
.Y(n_5013)
);

OAI21x1_ASAP7_75t_L g5014 ( 
.A1(n_4409),
.A2(n_781),
.B(n_780),
.Y(n_5014)
);

O2A1O1Ixp33_ASAP7_75t_L g5015 ( 
.A1(n_4738),
.A2(n_783),
.B(n_784),
.C(n_782),
.Y(n_5015)
);

NAND3xp33_ASAP7_75t_L g5016 ( 
.A(n_4749),
.B(n_784),
.C(n_783),
.Y(n_5016)
);

NAND2xp5_ASAP7_75t_L g5017 ( 
.A(n_4607),
.B(n_783),
.Y(n_5017)
);

OAI21x1_ASAP7_75t_SL g5018 ( 
.A1(n_4675),
.A2(n_786),
.B(n_785),
.Y(n_5018)
);

AOI21xp5_ASAP7_75t_L g5019 ( 
.A1(n_4367),
.A2(n_786),
.B(n_785),
.Y(n_5019)
);

AOI21x1_ASAP7_75t_L g5020 ( 
.A1(n_4299),
.A2(n_4587),
.B(n_4797),
.Y(n_5020)
);

AOI21xp5_ASAP7_75t_L g5021 ( 
.A1(n_4835),
.A2(n_786),
.B(n_785),
.Y(n_5021)
);

AOI21xp5_ASAP7_75t_L g5022 ( 
.A1(n_4835),
.A2(n_788),
.B(n_787),
.Y(n_5022)
);

CKINVDCx20_ASAP7_75t_R g5023 ( 
.A(n_4380),
.Y(n_5023)
);

INVx2_ASAP7_75t_L g5024 ( 
.A(n_4389),
.Y(n_5024)
);

NAND3xp33_ASAP7_75t_L g5025 ( 
.A(n_4491),
.B(n_788),
.C(n_787),
.Y(n_5025)
);

INVx1_ASAP7_75t_L g5026 ( 
.A(n_4596),
.Y(n_5026)
);

AND2x2_ASAP7_75t_L g5027 ( 
.A(n_4634),
.B(n_789),
.Y(n_5027)
);

NAND2xp5_ASAP7_75t_L g5028 ( 
.A(n_4622),
.B(n_789),
.Y(n_5028)
);

HB1xp67_ASAP7_75t_L g5029 ( 
.A(n_4441),
.Y(n_5029)
);

NOR2xp33_ASAP7_75t_L g5030 ( 
.A(n_4360),
.B(n_790),
.Y(n_5030)
);

AND2x4_ASAP7_75t_L g5031 ( 
.A(n_4579),
.B(n_4635),
.Y(n_5031)
);

INVx2_ASAP7_75t_L g5032 ( 
.A(n_4414),
.Y(n_5032)
);

AND2x4_ASAP7_75t_L g5033 ( 
.A(n_4662),
.B(n_790),
.Y(n_5033)
);

INVx3_ASAP7_75t_L g5034 ( 
.A(n_4402),
.Y(n_5034)
);

AOI221xp5_ASAP7_75t_SL g5035 ( 
.A1(n_4553),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.C(n_59),
.Y(n_5035)
);

OAI21x1_ASAP7_75t_L g5036 ( 
.A1(n_4820),
.A2(n_791),
.B(n_790),
.Y(n_5036)
);

INVx2_ASAP7_75t_SL g5037 ( 
.A(n_4659),
.Y(n_5037)
);

OAI21xp5_ASAP7_75t_L g5038 ( 
.A1(n_4792),
.A2(n_4799),
.B(n_4795),
.Y(n_5038)
);

NAND2xp5_ASAP7_75t_L g5039 ( 
.A(n_4655),
.B(n_791),
.Y(n_5039)
);

OAI21xp5_ASAP7_75t_L g5040 ( 
.A1(n_4455),
.A2(n_792),
.B(n_791),
.Y(n_5040)
);

OAI21xp33_ASAP7_75t_L g5041 ( 
.A1(n_4745),
.A2(n_793),
.B(n_792),
.Y(n_5041)
);

OAI21x1_ASAP7_75t_L g5042 ( 
.A1(n_4848),
.A2(n_794),
.B(n_793),
.Y(n_5042)
);

AOI21xp5_ASAP7_75t_L g5043 ( 
.A1(n_4835),
.A2(n_794),
.B(n_793),
.Y(n_5043)
);

AOI21xp5_ASAP7_75t_L g5044 ( 
.A1(n_4330),
.A2(n_795),
.B(n_794),
.Y(n_5044)
);

A2O1A1Ixp33_ASAP7_75t_L g5045 ( 
.A1(n_4670),
.A2(n_796),
.B(n_797),
.C(n_795),
.Y(n_5045)
);

BUFx2_ASAP7_75t_L g5046 ( 
.A(n_4762),
.Y(n_5046)
);

NAND2xp5_ASAP7_75t_L g5047 ( 
.A(n_4673),
.B(n_795),
.Y(n_5047)
);

A2O1A1Ixp33_ASAP7_75t_L g5048 ( 
.A1(n_4519),
.A2(n_797),
.B(n_798),
.C(n_796),
.Y(n_5048)
);

INVx2_ASAP7_75t_L g5049 ( 
.A(n_4454),
.Y(n_5049)
);

AOI21xp5_ASAP7_75t_L g5050 ( 
.A1(n_4358),
.A2(n_797),
.B(n_796),
.Y(n_5050)
);

OAI21x1_ASAP7_75t_L g5051 ( 
.A1(n_4460),
.A2(n_4548),
.B(n_4449),
.Y(n_5051)
);

OAI21x1_ASAP7_75t_L g5052 ( 
.A1(n_4428),
.A2(n_799),
.B(n_798),
.Y(n_5052)
);

NAND2xp5_ASAP7_75t_L g5053 ( 
.A(n_4678),
.B(n_798),
.Y(n_5053)
);

AOI21xp5_ASAP7_75t_L g5054 ( 
.A1(n_4326),
.A2(n_801),
.B(n_800),
.Y(n_5054)
);

OAI21x1_ASAP7_75t_L g5055 ( 
.A1(n_4428),
.A2(n_801),
.B(n_800),
.Y(n_5055)
);

OAI22xp5_ASAP7_75t_L g5056 ( 
.A1(n_4313),
.A2(n_802),
.B1(n_803),
.B2(n_801),
.Y(n_5056)
);

AOI21xp5_ASAP7_75t_L g5057 ( 
.A1(n_4819),
.A2(n_804),
.B(n_802),
.Y(n_5057)
);

OA21x2_ASAP7_75t_L g5058 ( 
.A1(n_4750),
.A2(n_4787),
.B(n_4832),
.Y(n_5058)
);

NAND2xp5_ASAP7_75t_L g5059 ( 
.A(n_4705),
.B(n_804),
.Y(n_5059)
);

OAI21xp5_ASAP7_75t_L g5060 ( 
.A1(n_4783),
.A2(n_806),
.B(n_805),
.Y(n_5060)
);

AOI21xp5_ASAP7_75t_L g5061 ( 
.A1(n_4336),
.A2(n_806),
.B(n_805),
.Y(n_5061)
);

O2A1O1Ixp5_ASAP7_75t_L g5062 ( 
.A1(n_4824),
.A2(n_806),
.B(n_807),
.C(n_805),
.Y(n_5062)
);

INVx2_ASAP7_75t_L g5063 ( 
.A(n_4474),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_4480),
.Y(n_5064)
);

AND2x4_ASAP7_75t_L g5065 ( 
.A(n_4668),
.B(n_807),
.Y(n_5065)
);

AND2x4_ASAP7_75t_L g5066 ( 
.A(n_4585),
.B(n_807),
.Y(n_5066)
);

AOI21xp5_ASAP7_75t_L g5067 ( 
.A1(n_4858),
.A2(n_809),
.B(n_808),
.Y(n_5067)
);

OAI22xp5_ASAP7_75t_L g5068 ( 
.A1(n_4341),
.A2(n_809),
.B1(n_810),
.B2(n_808),
.Y(n_5068)
);

NOR4xp25_ASAP7_75t_L g5069 ( 
.A(n_4468),
.B(n_809),
.C(n_810),
.D(n_808),
.Y(n_5069)
);

BUFx10_ASAP7_75t_L g5070 ( 
.A(n_4594),
.Y(n_5070)
);

AOI22xp33_ASAP7_75t_L g5071 ( 
.A1(n_4505),
.A2(n_812),
.B1(n_813),
.B2(n_811),
.Y(n_5071)
);

INVx1_ASAP7_75t_L g5072 ( 
.A(n_4490),
.Y(n_5072)
);

OAI21x1_ASAP7_75t_L g5073 ( 
.A1(n_4825),
.A2(n_813),
.B(n_811),
.Y(n_5073)
);

OAI21x1_ASAP7_75t_L g5074 ( 
.A1(n_4318),
.A2(n_4406),
.B(n_4698),
.Y(n_5074)
);

AOI21xp5_ASAP7_75t_SL g5075 ( 
.A1(n_4516),
.A2(n_813),
.B(n_811),
.Y(n_5075)
);

AOI21xp5_ASAP7_75t_L g5076 ( 
.A1(n_4861),
.A2(n_815),
.B(n_814),
.Y(n_5076)
);

OAI21x1_ASAP7_75t_L g5077 ( 
.A1(n_4698),
.A2(n_816),
.B(n_815),
.Y(n_5077)
);

AOI21xp5_ASAP7_75t_L g5078 ( 
.A1(n_4498),
.A2(n_816),
.B(n_815),
.Y(n_5078)
);

BUFx6f_ASAP7_75t_L g5079 ( 
.A(n_4656),
.Y(n_5079)
);

AOI21xp5_ASAP7_75t_L g5080 ( 
.A1(n_4535),
.A2(n_4563),
.B(n_4549),
.Y(n_5080)
);

NAND3xp33_ASAP7_75t_L g5081 ( 
.A(n_4653),
.B(n_817),
.C(n_816),
.Y(n_5081)
);

CKINVDCx16_ASAP7_75t_R g5082 ( 
.A(n_4495),
.Y(n_5082)
);

AOI22xp5_ASAP7_75t_L g5083 ( 
.A1(n_4726),
.A2(n_1148),
.B1(n_1152),
.B2(n_1147),
.Y(n_5083)
);

OR2x6_ASAP7_75t_L g5084 ( 
.A(n_4423),
.B(n_817),
.Y(n_5084)
);

OA21x2_ASAP7_75t_L g5085 ( 
.A1(n_4520),
.A2(n_818),
.B(n_817),
.Y(n_5085)
);

AOI21xp5_ASAP7_75t_L g5086 ( 
.A1(n_4589),
.A2(n_819),
.B(n_818),
.Y(n_5086)
);

NOR2xp33_ASAP7_75t_SL g5087 ( 
.A(n_4592),
.B(n_1159),
.Y(n_5087)
);

INVx2_ASAP7_75t_SL g5088 ( 
.A(n_4420),
.Y(n_5088)
);

AOI21xp5_ASAP7_75t_L g5089 ( 
.A1(n_4363),
.A2(n_820),
.B(n_819),
.Y(n_5089)
);

OAI22x1_ASAP7_75t_L g5090 ( 
.A1(n_4344),
.A2(n_820),
.B1(n_821),
.B2(n_819),
.Y(n_5090)
);

INVx4_ASAP7_75t_L g5091 ( 
.A(n_4752),
.Y(n_5091)
);

OAI21x1_ASAP7_75t_L g5092 ( 
.A1(n_4391),
.A2(n_821),
.B(n_820),
.Y(n_5092)
);

INVx2_ASAP7_75t_L g5093 ( 
.A(n_4605),
.Y(n_5093)
);

INVx1_ASAP7_75t_L g5094 ( 
.A(n_4619),
.Y(n_5094)
);

AOI21xp33_ASAP7_75t_L g5095 ( 
.A1(n_4309),
.A2(n_823),
.B(n_822),
.Y(n_5095)
);

AOI21xp5_ASAP7_75t_L g5096 ( 
.A1(n_4329),
.A2(n_823),
.B(n_822),
.Y(n_5096)
);

INVxp67_ASAP7_75t_L g5097 ( 
.A(n_4387),
.Y(n_5097)
);

OAI21xp5_ASAP7_75t_L g5098 ( 
.A1(n_4791),
.A2(n_823),
.B(n_822),
.Y(n_5098)
);

AOI21xp5_ASAP7_75t_SL g5099 ( 
.A1(n_4516),
.A2(n_825),
.B(n_824),
.Y(n_5099)
);

AND2x4_ASAP7_75t_L g5100 ( 
.A(n_4369),
.B(n_824),
.Y(n_5100)
);

INVx2_ASAP7_75t_L g5101 ( 
.A(n_4812),
.Y(n_5101)
);

NOR2xp67_ASAP7_75t_L g5102 ( 
.A(n_4545),
.B(n_827),
.Y(n_5102)
);

OAI22xp5_ASAP7_75t_L g5103 ( 
.A1(n_4371),
.A2(n_825),
.B1(n_826),
.B2(n_824),
.Y(n_5103)
);

OAI21x1_ASAP7_75t_L g5104 ( 
.A1(n_4842),
.A2(n_826),
.B(n_825),
.Y(n_5104)
);

NAND2xp5_ASAP7_75t_L g5105 ( 
.A(n_4741),
.B(n_827),
.Y(n_5105)
);

NAND3xp33_ASAP7_75t_L g5106 ( 
.A(n_4674),
.B(n_829),
.C(n_828),
.Y(n_5106)
);

INVx3_ASAP7_75t_L g5107 ( 
.A(n_4461),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_4377),
.Y(n_5108)
);

INVx4_ASAP7_75t_L g5109 ( 
.A(n_4365),
.Y(n_5109)
);

INVx2_ASAP7_75t_SL g5110 ( 
.A(n_4664),
.Y(n_5110)
);

OR2x2_ASAP7_75t_L g5111 ( 
.A(n_4343),
.B(n_828),
.Y(n_5111)
);

OAI21x1_ASAP7_75t_L g5112 ( 
.A1(n_4411),
.A2(n_829),
.B(n_828),
.Y(n_5112)
);

NAND2xp5_ASAP7_75t_L g5113 ( 
.A(n_4807),
.B(n_829),
.Y(n_5113)
);

AOI21xp5_ASAP7_75t_L g5114 ( 
.A1(n_4305),
.A2(n_831),
.B(n_830),
.Y(n_5114)
);

OAI21x1_ASAP7_75t_L g5115 ( 
.A1(n_4417),
.A2(n_831),
.B(n_830),
.Y(n_5115)
);

AOI21x1_ASAP7_75t_L g5116 ( 
.A1(n_4375),
.A2(n_832),
.B(n_830),
.Y(n_5116)
);

AOI21x1_ASAP7_75t_L g5117 ( 
.A1(n_4512),
.A2(n_833),
.B(n_832),
.Y(n_5117)
);

INVx2_ASAP7_75t_L g5118 ( 
.A(n_4794),
.Y(n_5118)
);

NOR2xp67_ASAP7_75t_L g5119 ( 
.A(n_4453),
.B(n_835),
.Y(n_5119)
);

OAI21xp5_ASAP7_75t_SL g5120 ( 
.A1(n_4746),
.A2(n_1147),
.B(n_1146),
.Y(n_5120)
);

NAND2xp5_ASAP7_75t_L g5121 ( 
.A(n_4809),
.B(n_832),
.Y(n_5121)
);

OAI21x1_ASAP7_75t_L g5122 ( 
.A1(n_4438),
.A2(n_834),
.B(n_833),
.Y(n_5122)
);

AOI22xp5_ASAP7_75t_L g5123 ( 
.A1(n_4851),
.A2(n_4524),
.B1(n_4434),
.B2(n_4415),
.Y(n_5123)
);

AOI22xp5_ASAP7_75t_L g5124 ( 
.A1(n_4475),
.A2(n_1157),
.B1(n_1160),
.B2(n_1148),
.Y(n_5124)
);

OAI21xp5_ASAP7_75t_L g5125 ( 
.A1(n_4818),
.A2(n_835),
.B(n_833),
.Y(n_5125)
);

A2O1A1Ixp33_ASAP7_75t_L g5126 ( 
.A1(n_4648),
.A2(n_836),
.B(n_837),
.C(n_835),
.Y(n_5126)
);

OAI21x1_ASAP7_75t_L g5127 ( 
.A1(n_4844),
.A2(n_837),
.B(n_836),
.Y(n_5127)
);

NAND2xp5_ASAP7_75t_L g5128 ( 
.A(n_4810),
.B(n_838),
.Y(n_5128)
);

INVx3_ASAP7_75t_L g5129 ( 
.A(n_4432),
.Y(n_5129)
);

BUFx12f_ASAP7_75t_L g5130 ( 
.A(n_4500),
.Y(n_5130)
);

OAI21x1_ASAP7_75t_L g5131 ( 
.A1(n_4852),
.A2(n_839),
.B(n_838),
.Y(n_5131)
);

OAI21xp5_ASAP7_75t_L g5132 ( 
.A1(n_4687),
.A2(n_840),
.B(n_839),
.Y(n_5132)
);

INVxp67_ASAP7_75t_L g5133 ( 
.A(n_4337),
.Y(n_5133)
);

OR2x2_ASAP7_75t_L g5134 ( 
.A(n_4510),
.B(n_839),
.Y(n_5134)
);

A2O1A1Ixp33_ASAP7_75t_L g5135 ( 
.A1(n_4701),
.A2(n_841),
.B(n_842),
.C(n_840),
.Y(n_5135)
);

O2A1O1Ixp33_ASAP7_75t_L g5136 ( 
.A1(n_4779),
.A2(n_841),
.B(n_842),
.C(n_840),
.Y(n_5136)
);

AND2x2_ASAP7_75t_L g5137 ( 
.A(n_4348),
.B(n_843),
.Y(n_5137)
);

OAI21x1_ASAP7_75t_L g5138 ( 
.A1(n_4854),
.A2(n_844),
.B(n_843),
.Y(n_5138)
);

OAI21xp5_ASAP7_75t_L g5139 ( 
.A1(n_4735),
.A2(n_845),
.B(n_844),
.Y(n_5139)
);

AOI21xp5_ASAP7_75t_L g5140 ( 
.A1(n_4305),
.A2(n_846),
.B(n_845),
.Y(n_5140)
);

OAI21x1_ASAP7_75t_L g5141 ( 
.A1(n_4794),
.A2(n_847),
.B(n_845),
.Y(n_5141)
);

BUFx6f_ASAP7_75t_L g5142 ( 
.A(n_4775),
.Y(n_5142)
);

OAI21x1_ASAP7_75t_L g5143 ( 
.A1(n_4836),
.A2(n_848),
.B(n_847),
.Y(n_5143)
);

INVx1_ASAP7_75t_L g5144 ( 
.A(n_4379),
.Y(n_5144)
);

INVxp67_ASAP7_75t_SL g5145 ( 
.A(n_4523),
.Y(n_5145)
);

AOI21xp5_ASAP7_75t_L g5146 ( 
.A1(n_4305),
.A2(n_848),
.B(n_847),
.Y(n_5146)
);

CKINVDCx20_ASAP7_75t_R g5147 ( 
.A(n_4614),
.Y(n_5147)
);

AND2x4_ASAP7_75t_L g5148 ( 
.A(n_4453),
.B(n_849),
.Y(n_5148)
);

NAND2xp5_ASAP7_75t_SL g5149 ( 
.A(n_4704),
.B(n_849),
.Y(n_5149)
);

NAND2xp5_ASAP7_75t_L g5150 ( 
.A(n_4618),
.B(n_849),
.Y(n_5150)
);

NAND2xp5_ASAP7_75t_L g5151 ( 
.A(n_4814),
.B(n_850),
.Y(n_5151)
);

AOI21xp5_ASAP7_75t_L g5152 ( 
.A1(n_4331),
.A2(n_851),
.B(n_850),
.Y(n_5152)
);

BUFx2_ASAP7_75t_R g5153 ( 
.A(n_4395),
.Y(n_5153)
);

NOR2xp33_ASAP7_75t_L g5154 ( 
.A(n_4672),
.B(n_850),
.Y(n_5154)
);

BUFx4_ASAP7_75t_SL g5155 ( 
.A(n_4359),
.Y(n_5155)
);

AOI21xp5_ASAP7_75t_L g5156 ( 
.A1(n_4331),
.A2(n_852),
.B(n_851),
.Y(n_5156)
);

AOI21xp5_ASAP7_75t_SL g5157 ( 
.A1(n_4425),
.A2(n_852),
.B(n_851),
.Y(n_5157)
);

OAI21x1_ASAP7_75t_SL g5158 ( 
.A1(n_4547),
.A2(n_853),
.B(n_852),
.Y(n_5158)
);

BUFx2_ASAP7_75t_L g5159 ( 
.A(n_4372),
.Y(n_5159)
);

A2O1A1Ixp33_ASAP7_75t_L g5160 ( 
.A1(n_4718),
.A2(n_854),
.B(n_855),
.C(n_853),
.Y(n_5160)
);

O2A1O1Ixp33_ASAP7_75t_SL g5161 ( 
.A1(n_4604),
.A2(n_855),
.B(n_856),
.C(n_854),
.Y(n_5161)
);

INVxp67_ASAP7_75t_L g5162 ( 
.A(n_4447),
.Y(n_5162)
);

NAND2xp5_ASAP7_75t_L g5163 ( 
.A(n_4610),
.B(n_854),
.Y(n_5163)
);

AND2x2_ASAP7_75t_L g5164 ( 
.A(n_4531),
.B(n_856),
.Y(n_5164)
);

AND2x4_ASAP7_75t_L g5165 ( 
.A(n_4636),
.B(n_856),
.Y(n_5165)
);

AND2x2_ASAP7_75t_L g5166 ( 
.A(n_4364),
.B(n_857),
.Y(n_5166)
);

INVx2_ASAP7_75t_L g5167 ( 
.A(n_4693),
.Y(n_5167)
);

INVx1_ASAP7_75t_L g5168 ( 
.A(n_4421),
.Y(n_5168)
);

INVx3_ASAP7_75t_SL g5169 ( 
.A(n_4431),
.Y(n_5169)
);

NAND2xp5_ASAP7_75t_L g5170 ( 
.A(n_4542),
.B(n_4567),
.Y(n_5170)
);

AOI21xp5_ASAP7_75t_L g5171 ( 
.A1(n_4331),
.A2(n_858),
.B(n_857),
.Y(n_5171)
);

AO31x2_ASAP7_75t_L g5172 ( 
.A1(n_4847),
.A2(n_858),
.A3(n_859),
.B(n_857),
.Y(n_5172)
);

OAI21x1_ASAP7_75t_L g5173 ( 
.A1(n_4467),
.A2(n_4734),
.B(n_4806),
.Y(n_5173)
);

NAND2xp5_ASAP7_75t_SL g5174 ( 
.A(n_4704),
.B(n_4747),
.Y(n_5174)
);

AOI21x1_ASAP7_75t_L g5175 ( 
.A1(n_4569),
.A2(n_859),
.B(n_858),
.Y(n_5175)
);

INVx1_ASAP7_75t_L g5176 ( 
.A(n_4429),
.Y(n_5176)
);

HB1xp67_ASAP7_75t_L g5177 ( 
.A(n_4459),
.Y(n_5177)
);

NAND2xp5_ASAP7_75t_L g5178 ( 
.A(n_4560),
.B(n_859),
.Y(n_5178)
);

NAND3xp33_ASAP7_75t_L g5179 ( 
.A(n_4419),
.B(n_861),
.C(n_860),
.Y(n_5179)
);

INVx1_ASAP7_75t_L g5180 ( 
.A(n_4445),
.Y(n_5180)
);

OAI21x1_ASAP7_75t_L g5181 ( 
.A1(n_4863),
.A2(n_861),
.B(n_860),
.Y(n_5181)
);

BUFx3_ASAP7_75t_L g5182 ( 
.A(n_4477),
.Y(n_5182)
);

AOI21xp5_ASAP7_75t_L g5183 ( 
.A1(n_4355),
.A2(n_861),
.B(n_860),
.Y(n_5183)
);

OAI21x1_ASAP7_75t_L g5184 ( 
.A1(n_4765),
.A2(n_863),
.B(n_862),
.Y(n_5184)
);

INVx1_ASAP7_75t_L g5185 ( 
.A(n_4446),
.Y(n_5185)
);

AND2x2_ASAP7_75t_L g5186 ( 
.A(n_4407),
.B(n_862),
.Y(n_5186)
);

AOI21xp5_ASAP7_75t_L g5187 ( 
.A1(n_4355),
.A2(n_863),
.B(n_862),
.Y(n_5187)
);

AOI21xp5_ASAP7_75t_L g5188 ( 
.A1(n_4355),
.A2(n_4442),
.B(n_4397),
.Y(n_5188)
);

AO32x2_ASAP7_75t_L g5189 ( 
.A1(n_4699),
.A2(n_865),
.A3(n_866),
.B1(n_864),
.B2(n_863),
.Y(n_5189)
);

INVx3_ASAP7_75t_L g5190 ( 
.A(n_4444),
.Y(n_5190)
);

BUFx6f_ASAP7_75t_L g5191 ( 
.A(n_4704),
.Y(n_5191)
);

AO32x2_ASAP7_75t_L g5192 ( 
.A1(n_4676),
.A2(n_4784),
.A3(n_4504),
.B1(n_4588),
.B2(n_4719),
.Y(n_5192)
);

AND2x2_ASAP7_75t_L g5193 ( 
.A(n_4400),
.B(n_4763),
.Y(n_5193)
);

OAI21x1_ASAP7_75t_L g5194 ( 
.A1(n_4731),
.A2(n_865),
.B(n_864),
.Y(n_5194)
);

AND2x2_ASAP7_75t_L g5195 ( 
.A(n_4513),
.B(n_866),
.Y(n_5195)
);

NAND2xp5_ASAP7_75t_L g5196 ( 
.A(n_4798),
.B(n_866),
.Y(n_5196)
);

HB1xp67_ASAP7_75t_L g5197 ( 
.A(n_4575),
.Y(n_5197)
);

OAI21x1_ASAP7_75t_L g5198 ( 
.A1(n_4451),
.A2(n_868),
.B(n_867),
.Y(n_5198)
);

NOR2xp33_ASAP7_75t_L g5199 ( 
.A(n_4328),
.B(n_867),
.Y(n_5199)
);

NAND2xp5_ASAP7_75t_L g5200 ( 
.A(n_4464),
.B(n_867),
.Y(n_5200)
);

OAI21x1_ASAP7_75t_L g5201 ( 
.A1(n_4649),
.A2(n_869),
.B(n_868),
.Y(n_5201)
);

NAND2xp5_ASAP7_75t_L g5202 ( 
.A(n_4511),
.B(n_868),
.Y(n_5202)
);

AO32x2_ASAP7_75t_L g5203 ( 
.A1(n_4496),
.A2(n_888),
.A3(n_896),
.B1(n_880),
.B2(n_872),
.Y(n_5203)
);

NOR2xp33_ASAP7_75t_L g5204 ( 
.A(n_4404),
.B(n_869),
.Y(n_5204)
);

OR2x6_ASAP7_75t_L g5205 ( 
.A(n_4416),
.B(n_869),
.Y(n_5205)
);

NAND2xp5_ASAP7_75t_L g5206 ( 
.A(n_4590),
.B(n_870),
.Y(n_5206)
);

INVx1_ASAP7_75t_L g5207 ( 
.A(n_4558),
.Y(n_5207)
);

NAND2x1p5_ASAP7_75t_L g5208 ( 
.A(n_4586),
.B(n_870),
.Y(n_5208)
);

INVx1_ASAP7_75t_L g5209 ( 
.A(n_4577),
.Y(n_5209)
);

NAND3xp33_ASAP7_75t_SL g5210 ( 
.A(n_4506),
.B(n_56),
.C(n_57),
.Y(n_5210)
);

NAND2xp5_ASAP7_75t_L g5211 ( 
.A(n_4476),
.B(n_870),
.Y(n_5211)
);

AOI221x1_ASAP7_75t_L g5212 ( 
.A1(n_4541),
.A2(n_874),
.B1(n_875),
.B2(n_873),
.C(n_871),
.Y(n_5212)
);

AO31x2_ASAP7_75t_L g5213 ( 
.A1(n_4754),
.A2(n_4804),
.A3(n_4615),
.B(n_4753),
.Y(n_5213)
);

OAI21x1_ASAP7_75t_L g5214 ( 
.A1(n_4758),
.A2(n_873),
.B(n_871),
.Y(n_5214)
);

AOI21x1_ASAP7_75t_L g5215 ( 
.A1(n_4540),
.A2(n_874),
.B(n_871),
.Y(n_5215)
);

NOR2xp33_ASAP7_75t_L g5216 ( 
.A(n_4332),
.B(n_874),
.Y(n_5216)
);

HB1xp67_ASAP7_75t_L g5217 ( 
.A(n_4710),
.Y(n_5217)
);

OAI21x1_ASAP7_75t_L g5218 ( 
.A1(n_4606),
.A2(n_876),
.B(n_875),
.Y(n_5218)
);

OAI21x1_ASAP7_75t_L g5219 ( 
.A1(n_4711),
.A2(n_877),
.B(n_876),
.Y(n_5219)
);

AO31x2_ASAP7_75t_L g5220 ( 
.A1(n_4489),
.A2(n_4823),
.A3(n_4529),
.B(n_4574),
.Y(n_5220)
);

AOI21xp5_ASAP7_75t_L g5221 ( 
.A1(n_4397),
.A2(n_877),
.B(n_876),
.Y(n_5221)
);

INVx2_ASAP7_75t_L g5222 ( 
.A(n_4397),
.Y(n_5222)
);

OAI21x1_ASAP7_75t_L g5223 ( 
.A1(n_4729),
.A2(n_4766),
.B(n_4764),
.Y(n_5223)
);

NAND2xp5_ASAP7_75t_L g5224 ( 
.A(n_4790),
.B(n_878),
.Y(n_5224)
);

INVx2_ASAP7_75t_SL g5225 ( 
.A(n_4564),
.Y(n_5225)
);

NOR2xp67_ASAP7_75t_L g5226 ( 
.A(n_4430),
.B(n_883),
.Y(n_5226)
);

OAI21x1_ASAP7_75t_L g5227 ( 
.A1(n_4720),
.A2(n_879),
.B(n_878),
.Y(n_5227)
);

AND2x2_ASAP7_75t_L g5228 ( 
.A(n_4412),
.B(n_879),
.Y(n_5228)
);

INVx1_ASAP7_75t_L g5229 ( 
.A(n_4584),
.Y(n_5229)
);

O2A1O1Ixp33_ASAP7_75t_L g5230 ( 
.A1(n_4552),
.A2(n_881),
.B(n_882),
.C(n_879),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_4786),
.Y(n_5231)
);

AOI221x1_ASAP7_75t_L g5232 ( 
.A1(n_4721),
.A2(n_884),
.B1(n_885),
.B2(n_883),
.C(n_881),
.Y(n_5232)
);

INVx3_ASAP7_75t_L g5233 ( 
.A(n_4583),
.Y(n_5233)
);

AOI22xp5_ASAP7_75t_L g5234 ( 
.A1(n_4654),
.A2(n_884),
.B1(n_886),
.B2(n_881),
.Y(n_5234)
);

AOI21xp5_ASAP7_75t_L g5235 ( 
.A1(n_4442),
.A2(n_886),
.B(n_884),
.Y(n_5235)
);

INVx2_ASAP7_75t_SL g5236 ( 
.A(n_4776),
.Y(n_5236)
);

BUFx2_ASAP7_75t_L g5237 ( 
.A(n_4686),
.Y(n_5237)
);

AOI21xp5_ASAP7_75t_L g5238 ( 
.A1(n_4442),
.A2(n_888),
.B(n_887),
.Y(n_5238)
);

AND2x2_ASAP7_75t_L g5239 ( 
.A(n_4518),
.B(n_889),
.Y(n_5239)
);

INVx1_ASAP7_75t_L g5240 ( 
.A(n_4786),
.Y(n_5240)
);

NOR2xp33_ASAP7_75t_L g5241 ( 
.A(n_4382),
.B(n_890),
.Y(n_5241)
);

AO21x2_ASAP7_75t_L g5242 ( 
.A1(n_4782),
.A2(n_891),
.B(n_890),
.Y(n_5242)
);

AO21x2_ASAP7_75t_L g5243 ( 
.A1(n_4743),
.A2(n_891),
.B(n_890),
.Y(n_5243)
);

INVx1_ASAP7_75t_L g5244 ( 
.A(n_4786),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_4786),
.Y(n_5245)
);

INVx4_ASAP7_75t_L g5246 ( 
.A(n_4708),
.Y(n_5246)
);

NAND3xp33_ASAP7_75t_L g5247 ( 
.A(n_4651),
.B(n_4632),
.C(n_4582),
.Y(n_5247)
);

BUFx6f_ASAP7_75t_L g5248 ( 
.A(n_4482),
.Y(n_5248)
);

OA22x2_ASAP7_75t_L g5249 ( 
.A1(n_4437),
.A2(n_893),
.B1(n_894),
.B2(n_892),
.Y(n_5249)
);

INVx5_ASAP7_75t_L g5250 ( 
.A(n_4482),
.Y(n_5250)
);

INVx1_ASAP7_75t_L g5251 ( 
.A(n_4866),
.Y(n_5251)
);

NAND2xp5_ASAP7_75t_L g5252 ( 
.A(n_4789),
.B(n_892),
.Y(n_5252)
);

INVx2_ASAP7_75t_L g5253 ( 
.A(n_4482),
.Y(n_5253)
);

NAND2xp5_ASAP7_75t_L g5254 ( 
.A(n_4816),
.B(n_892),
.Y(n_5254)
);

A2O1A1Ixp33_ASAP7_75t_L g5255 ( 
.A1(n_4715),
.A2(n_894),
.B(n_895),
.C(n_893),
.Y(n_5255)
);

INVxp67_ASAP7_75t_L g5256 ( 
.A(n_4501),
.Y(n_5256)
);

AOI21xp5_ASAP7_75t_SL g5257 ( 
.A1(n_4538),
.A2(n_895),
.B(n_893),
.Y(n_5257)
);

INVx3_ASAP7_75t_L g5258 ( 
.A(n_4768),
.Y(n_5258)
);

A2O1A1Ixp33_ASAP7_75t_L g5259 ( 
.A1(n_4497),
.A2(n_897),
.B(n_898),
.C(n_896),
.Y(n_5259)
);

NAND2xp5_ASAP7_75t_SL g5260 ( 
.A(n_4747),
.B(n_897),
.Y(n_5260)
);

AOI221xp5_ASAP7_75t_L g5261 ( 
.A1(n_4544),
.A2(n_899),
.B1(n_900),
.B2(n_898),
.C(n_897),
.Y(n_5261)
);

NAND2xp5_ASAP7_75t_L g5262 ( 
.A(n_4646),
.B(n_4650),
.Y(n_5262)
);

INVx3_ASAP7_75t_L g5263 ( 
.A(n_4802),
.Y(n_5263)
);

AOI221xp5_ASAP7_75t_SL g5264 ( 
.A1(n_4383),
.A2(n_4393),
.B1(n_4756),
.B2(n_4509),
.C(n_4536),
.Y(n_5264)
);

A2O1A1Ixp33_ASAP7_75t_L g5265 ( 
.A1(n_4657),
.A2(n_899),
.B(n_901),
.C(n_898),
.Y(n_5265)
);

NOR2xp33_ASAP7_75t_L g5266 ( 
.A(n_4366),
.B(n_901),
.Y(n_5266)
);

OAI22x1_ASAP7_75t_L g5267 ( 
.A1(n_4427),
.A2(n_902),
.B1(n_903),
.B2(n_901),
.Y(n_5267)
);

AOI21xp5_ASAP7_75t_L g5268 ( 
.A1(n_4488),
.A2(n_4562),
.B(n_4514),
.Y(n_5268)
);

NAND2xp5_ASAP7_75t_SL g5269 ( 
.A(n_4747),
.B(n_902),
.Y(n_5269)
);

OR2x2_ASAP7_75t_L g5270 ( 
.A(n_4733),
.B(n_903),
.Y(n_5270)
);

AOI221x1_ASAP7_75t_L g5271 ( 
.A1(n_4644),
.A2(n_905),
.B1(n_906),
.B2(n_904),
.C(n_903),
.Y(n_5271)
);

INVx1_ASAP7_75t_L g5272 ( 
.A(n_4866),
.Y(n_5272)
);

OAI21x1_ASAP7_75t_L g5273 ( 
.A1(n_4846),
.A2(n_905),
.B(n_904),
.Y(n_5273)
);

O2A1O1Ixp33_ASAP7_75t_L g5274 ( 
.A1(n_4499),
.A2(n_905),
.B(n_906),
.C(n_904),
.Y(n_5274)
);

INVx2_ASAP7_75t_SL g5275 ( 
.A(n_4802),
.Y(n_5275)
);

NAND2xp5_ASAP7_75t_L g5276 ( 
.A(n_4617),
.B(n_907),
.Y(n_5276)
);

AOI22xp5_ASAP7_75t_L g5277 ( 
.A1(n_4345),
.A2(n_1143),
.B1(n_1144),
.B2(n_1142),
.Y(n_5277)
);

OAI21x1_ASAP7_75t_L g5278 ( 
.A1(n_4827),
.A2(n_908),
.B(n_907),
.Y(n_5278)
);

OAI21xp5_ASAP7_75t_L g5279 ( 
.A1(n_4833),
.A2(n_910),
.B(n_908),
.Y(n_5279)
);

OR2x6_ASAP7_75t_L g5280 ( 
.A(n_4838),
.B(n_908),
.Y(n_5280)
);

AO21x1_ASAP7_75t_L g5281 ( 
.A1(n_4543),
.A2(n_4566),
.B(n_4554),
.Y(n_5281)
);

O2A1O1Ixp33_ASAP7_75t_L g5282 ( 
.A1(n_4325),
.A2(n_911),
.B(n_912),
.C(n_910),
.Y(n_5282)
);

AOI21xp5_ASAP7_75t_SL g5283 ( 
.A1(n_4457),
.A2(n_913),
.B(n_912),
.Y(n_5283)
);

OAI21x1_ASAP7_75t_L g5284 ( 
.A1(n_4381),
.A2(n_913),
.B(n_912),
.Y(n_5284)
);

INVx1_ASAP7_75t_L g5285 ( 
.A(n_4866),
.Y(n_5285)
);

HB1xp67_ASAP7_75t_L g5286 ( 
.A(n_4802),
.Y(n_5286)
);

OAI21xp5_ASAP7_75t_L g5287 ( 
.A1(n_4822),
.A2(n_915),
.B(n_914),
.Y(n_5287)
);

NAND2xp5_ASAP7_75t_L g5288 ( 
.A(n_4727),
.B(n_4631),
.Y(n_5288)
);

OAI22xp5_ASAP7_75t_L g5289 ( 
.A1(n_4521),
.A2(n_4788),
.B1(n_4805),
.B2(n_4801),
.Y(n_5289)
);

AOI21xp5_ASAP7_75t_L g5290 ( 
.A1(n_4488),
.A2(n_915),
.B(n_914),
.Y(n_5290)
);

AOI22xp5_ASAP7_75t_L g5291 ( 
.A1(n_4849),
.A2(n_1164),
.B1(n_1160),
.B2(n_916),
.Y(n_5291)
);

CKINVDCx20_ASAP7_75t_R g5292 ( 
.A(n_4817),
.Y(n_5292)
);

AOI21xp5_ASAP7_75t_L g5293 ( 
.A1(n_4488),
.A2(n_916),
.B(n_914),
.Y(n_5293)
);

BUFx3_ASAP7_75t_L g5294 ( 
.A(n_4679),
.Y(n_5294)
);

INVx2_ASAP7_75t_SL g5295 ( 
.A(n_4761),
.Y(n_5295)
);

NAND2xp5_ASAP7_75t_L g5296 ( 
.A(n_4528),
.B(n_916),
.Y(n_5296)
);

NAND2xp5_ASAP7_75t_L g5297 ( 
.A(n_4702),
.B(n_917),
.Y(n_5297)
);

AND2x2_ASAP7_75t_L g5298 ( 
.A(n_4838),
.B(n_4757),
.Y(n_5298)
);

OAI22xp5_ASAP7_75t_L g5299 ( 
.A1(n_4660),
.A2(n_918),
.B1(n_919),
.B2(n_917),
.Y(n_5299)
);

NAND2xp5_ASAP7_75t_L g5300 ( 
.A(n_4707),
.B(n_918),
.Y(n_5300)
);

OAI21xp33_ASAP7_75t_L g5301 ( 
.A1(n_4667),
.A2(n_919),
.B(n_918),
.Y(n_5301)
);

AOI211x1_ASAP7_75t_L g5302 ( 
.A1(n_4507),
.A2(n_921),
.B(n_922),
.C(n_920),
.Y(n_5302)
);

INVx1_ASAP7_75t_L g5303 ( 
.A(n_4808),
.Y(n_5303)
);

AOI221x1_ASAP7_75t_L g5304 ( 
.A1(n_4537),
.A2(n_922),
.B1(n_923),
.B2(n_921),
.C(n_920),
.Y(n_5304)
);

INVx1_ASAP7_75t_L g5305 ( 
.A(n_4808),
.Y(n_5305)
);

HB1xp67_ASAP7_75t_L g5306 ( 
.A(n_4773),
.Y(n_5306)
);

OR2x6_ASAP7_75t_L g5307 ( 
.A(n_4439),
.B(n_920),
.Y(n_5307)
);

AOI21xp5_ASAP7_75t_L g5308 ( 
.A1(n_4514),
.A2(n_922),
.B(n_921),
.Y(n_5308)
);

INVx3_ASAP7_75t_SL g5309 ( 
.A(n_4514),
.Y(n_5309)
);

INVxp67_ASAP7_75t_L g5310 ( 
.A(n_4759),
.Y(n_5310)
);

AOI21xp5_ASAP7_75t_L g5311 ( 
.A1(n_4562),
.A2(n_924),
.B(n_923),
.Y(n_5311)
);

AOI21xp5_ASAP7_75t_L g5312 ( 
.A1(n_4562),
.A2(n_4613),
.B(n_4602),
.Y(n_5312)
);

OAI21x1_ASAP7_75t_L g5313 ( 
.A1(n_4830),
.A2(n_924),
.B(n_923),
.Y(n_5313)
);

AND2x2_ASAP7_75t_L g5314 ( 
.A(n_4769),
.B(n_4772),
.Y(n_5314)
);

NAND2xp5_ASAP7_75t_L g5315 ( 
.A(n_4713),
.B(n_924),
.Y(n_5315)
);

OAI21x1_ASAP7_75t_L g5316 ( 
.A1(n_4837),
.A2(n_926),
.B(n_925),
.Y(n_5316)
);

NOR2xp33_ASAP7_75t_L g5317 ( 
.A(n_4717),
.B(n_925),
.Y(n_5317)
);

INVx1_ASAP7_75t_SL g5318 ( 
.A(n_4602),
.Y(n_5318)
);

INVx1_ASAP7_75t_L g5319 ( 
.A(n_4808),
.Y(n_5319)
);

AND2x2_ASAP7_75t_L g5320 ( 
.A(n_4728),
.B(n_4732),
.Y(n_5320)
);

AO32x2_ASAP7_75t_L g5321 ( 
.A1(n_4502),
.A2(n_928),
.A3(n_929),
.B1(n_927),
.B2(n_926),
.Y(n_5321)
);

OAI21xp5_ASAP7_75t_L g5322 ( 
.A1(n_4685),
.A2(n_4737),
.B(n_4723),
.Y(n_5322)
);

INVx3_ASAP7_75t_L g5323 ( 
.A(n_4602),
.Y(n_5323)
);

O2A1O1Ixp5_ASAP7_75t_L g5324 ( 
.A1(n_4517),
.A2(n_4530),
.B(n_4534),
.C(n_4663),
.Y(n_5324)
);

OAI21xp5_ASAP7_75t_L g5325 ( 
.A1(n_4751),
.A2(n_928),
.B(n_926),
.Y(n_5325)
);

AOI21xp5_ASAP7_75t_L g5326 ( 
.A1(n_4613),
.A2(n_929),
.B(n_928),
.Y(n_5326)
);

OAI21xp33_ASAP7_75t_L g5327 ( 
.A1(n_4600),
.A2(n_930),
.B(n_929),
.Y(n_5327)
);

INVx1_ASAP7_75t_L g5328 ( 
.A(n_4821),
.Y(n_5328)
);

NAND2xp5_ASAP7_75t_L g5329 ( 
.A(n_4744),
.B(n_930),
.Y(n_5329)
);

OAI21xp5_ASAP7_75t_L g5330 ( 
.A1(n_4755),
.A2(n_931),
.B(n_930),
.Y(n_5330)
);

NAND2xp5_ASAP7_75t_L g5331 ( 
.A(n_4611),
.B(n_931),
.Y(n_5331)
);

OAI21xp5_ASAP7_75t_L g5332 ( 
.A1(n_4793),
.A2(n_933),
.B(n_931),
.Y(n_5332)
);

AND2x2_ASAP7_75t_L g5333 ( 
.A(n_4609),
.B(n_933),
.Y(n_5333)
);

AOI21xp5_ASAP7_75t_L g5334 ( 
.A1(n_4613),
.A2(n_934),
.B(n_933),
.Y(n_5334)
);

AND2x4_ASAP7_75t_L g5335 ( 
.A(n_4862),
.B(n_934),
.Y(n_5335)
);

OAI21x1_ASAP7_75t_L g5336 ( 
.A1(n_4469),
.A2(n_935),
.B(n_934),
.Y(n_5336)
);

AOI21xp5_ASAP7_75t_L g5337 ( 
.A1(n_4625),
.A2(n_937),
.B(n_936),
.Y(n_5337)
);

OAI22xp5_ASAP7_75t_L g5338 ( 
.A1(n_4800),
.A2(n_4857),
.B1(n_4796),
.B2(n_4637),
.Y(n_5338)
);

OAI21x1_ASAP7_75t_L g5339 ( 
.A1(n_4559),
.A2(n_4572),
.B(n_4571),
.Y(n_5339)
);

AO31x2_ASAP7_75t_L g5340 ( 
.A1(n_4829),
.A2(n_937),
.A3(n_938),
.B(n_936),
.Y(n_5340)
);

AOI21x1_ASAP7_75t_L g5341 ( 
.A1(n_4862),
.A2(n_937),
.B(n_936),
.Y(n_5341)
);

INVx2_ASAP7_75t_SL g5342 ( 
.A(n_4625),
.Y(n_5342)
);

NAND2xp5_ASAP7_75t_L g5343 ( 
.A(n_4599),
.B(n_938),
.Y(n_5343)
);

CKINVDCx5p33_ASAP7_75t_R g5344 ( 
.A(n_4555),
.Y(n_5344)
);

AND2x4_ASAP7_75t_L g5345 ( 
.A(n_4625),
.B(n_938),
.Y(n_5345)
);

INVx1_ASAP7_75t_L g5346 ( 
.A(n_4869),
.Y(n_5346)
);

OAI21x1_ASAP7_75t_L g5347 ( 
.A1(n_4871),
.A2(n_4628),
.B(n_4601),
.Y(n_5347)
);

NAND2xp5_ASAP7_75t_L g5348 ( 
.A(n_5101),
.B(n_4595),
.Y(n_5348)
);

AOI22x1_ASAP7_75t_L g5349 ( 
.A1(n_4934),
.A2(n_4900),
.B1(n_5046),
.B2(n_5082),
.Y(n_5349)
);

OR2x2_ASAP7_75t_L g5350 ( 
.A(n_5003),
.B(n_4811),
.Y(n_5350)
);

NAND2xp5_ASAP7_75t_L g5351 ( 
.A(n_5328),
.B(n_4620),
.Y(n_5351)
);

INVx1_ASAP7_75t_L g5352 ( 
.A(n_4919),
.Y(n_5352)
);

OAI21x1_ASAP7_75t_L g5353 ( 
.A1(n_4898),
.A2(n_4683),
.B(n_4612),
.Y(n_5353)
);

BUFx2_ASAP7_75t_L g5354 ( 
.A(n_5109),
.Y(n_5354)
);

NOR2xp67_ASAP7_75t_L g5355 ( 
.A(n_4882),
.B(n_4714),
.Y(n_5355)
);

OA21x2_ASAP7_75t_L g5356 ( 
.A1(n_4995),
.A2(n_4591),
.B(n_4573),
.Y(n_5356)
);

BUFx3_ASAP7_75t_L g5357 ( 
.A(n_4914),
.Y(n_5357)
);

INVx1_ASAP7_75t_L g5358 ( 
.A(n_4921),
.Y(n_5358)
);

AND2x2_ASAP7_75t_L g5359 ( 
.A(n_4947),
.B(n_4627),
.Y(n_5359)
);

INVx3_ASAP7_75t_L g5360 ( 
.A(n_4868),
.Y(n_5360)
);

NAND3xp33_ASAP7_75t_L g5361 ( 
.A(n_4922),
.B(n_4624),
.C(n_4623),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_4926),
.Y(n_5362)
);

AOI222xp33_ASAP7_75t_L g5363 ( 
.A1(n_5007),
.A2(n_4839),
.B1(n_4843),
.B2(n_4853),
.C1(n_4576),
.C2(n_4640),
.Y(n_5363)
);

INVx1_ASAP7_75t_L g5364 ( 
.A(n_4956),
.Y(n_5364)
);

AOI22xp33_ASAP7_75t_L g5365 ( 
.A1(n_4905),
.A2(n_4641),
.B1(n_4694),
.B2(n_4859),
.Y(n_5365)
);

O2A1O1Ixp33_ASAP7_75t_SL g5366 ( 
.A1(n_4870),
.A2(n_4374),
.B(n_4486),
.C(n_4503),
.Y(n_5366)
);

INVx2_ASAP7_75t_SL g5367 ( 
.A(n_4892),
.Y(n_5367)
);

OAI21xp5_ASAP7_75t_L g5368 ( 
.A1(n_4902),
.A2(n_4608),
.B(n_4597),
.Y(n_5368)
);

OAI22xp33_ASAP7_75t_L g5369 ( 
.A1(n_5280),
.A2(n_4855),
.B1(n_4815),
.B2(n_4845),
.Y(n_5369)
);

OAI21x1_ASAP7_75t_L g5370 ( 
.A1(n_5074),
.A2(n_4680),
.B(n_4616),
.Y(n_5370)
);

OAI21x1_ASAP7_75t_L g5371 ( 
.A1(n_5188),
.A2(n_4645),
.B(n_4629),
.Y(n_5371)
);

INVx3_ASAP7_75t_L g5372 ( 
.A(n_4940),
.Y(n_5372)
);

NAND2xp5_ASAP7_75t_L g5373 ( 
.A(n_4987),
.B(n_4695),
.Y(n_5373)
);

AOI22xp5_ASAP7_75t_L g5374 ( 
.A1(n_5280),
.A2(n_4408),
.B1(n_4479),
.B2(n_4478),
.Y(n_5374)
);

OAI21x1_ASAP7_75t_L g5375 ( 
.A1(n_5268),
.A2(n_4712),
.B(n_4684),
.Y(n_5375)
);

AOI21xp33_ASAP7_75t_L g5376 ( 
.A1(n_4958),
.A2(n_4682),
.B(n_4642),
.Y(n_5376)
);

OAI21x1_ASAP7_75t_L g5377 ( 
.A1(n_5312),
.A2(n_4730),
.B(n_4692),
.Y(n_5377)
);

INVx2_ASAP7_75t_L g5378 ( 
.A(n_4969),
.Y(n_5378)
);

AO31x2_ASAP7_75t_L g5379 ( 
.A1(n_5118),
.A2(n_4422),
.A3(n_4471),
.B(n_4681),
.Y(n_5379)
);

OAI21x1_ASAP7_75t_L g5380 ( 
.A1(n_4879),
.A2(n_4706),
.B(n_4725),
.Y(n_5380)
);

INVx3_ASAP7_75t_L g5381 ( 
.A(n_4940),
.Y(n_5381)
);

BUFx2_ASAP7_75t_L g5382 ( 
.A(n_5182),
.Y(n_5382)
);

AOI22xp33_ASAP7_75t_L g5383 ( 
.A1(n_4973),
.A2(n_4815),
.B1(n_4630),
.B2(n_4700),
.Y(n_5383)
);

INVx1_ASAP7_75t_L g5384 ( 
.A(n_4966),
.Y(n_5384)
);

INVx2_ASAP7_75t_L g5385 ( 
.A(n_5005),
.Y(n_5385)
);

AND2x2_ASAP7_75t_L g5386 ( 
.A(n_5193),
.B(n_4627),
.Y(n_5386)
);

OR2x6_ASAP7_75t_L g5387 ( 
.A(n_4927),
.B(n_5084),
.Y(n_5387)
);

AND2x4_ASAP7_75t_L g5388 ( 
.A(n_4891),
.B(n_4627),
.Y(n_5388)
);

INVx3_ASAP7_75t_L g5389 ( 
.A(n_4891),
.Y(n_5389)
);

OAI21xp5_ASAP7_75t_L g5390 ( 
.A1(n_4923),
.A2(n_4813),
.B(n_4864),
.Y(n_5390)
);

INVx1_ASAP7_75t_L g5391 ( 
.A(n_4975),
.Y(n_5391)
);

OR2x2_ASAP7_75t_L g5392 ( 
.A(n_5029),
.B(n_939),
.Y(n_5392)
);

OR2x6_ASAP7_75t_L g5393 ( 
.A(n_4927),
.B(n_4815),
.Y(n_5393)
);

OAI21xp5_ASAP7_75t_L g5394 ( 
.A1(n_5016),
.A2(n_940),
.B(n_939),
.Y(n_5394)
);

INVx2_ASAP7_75t_L g5395 ( 
.A(n_5024),
.Y(n_5395)
);

NAND2xp5_ASAP7_75t_L g5396 ( 
.A(n_5108),
.B(n_4652),
.Y(n_5396)
);

OAI21xp5_ASAP7_75t_L g5397 ( 
.A1(n_5119),
.A2(n_940),
.B(n_939),
.Y(n_5397)
);

O2A1O1Ixp33_ASAP7_75t_SL g5398 ( 
.A1(n_4997),
.A2(n_942),
.B(n_943),
.C(n_941),
.Y(n_5398)
);

INVx1_ASAP7_75t_L g5399 ( 
.A(n_4910),
.Y(n_5399)
);

INVx1_ASAP7_75t_L g5400 ( 
.A(n_4953),
.Y(n_5400)
);

INVx1_ASAP7_75t_L g5401 ( 
.A(n_5002),
.Y(n_5401)
);

AND2x2_ASAP7_75t_L g5402 ( 
.A(n_4867),
.B(n_4652),
.Y(n_5402)
);

AND2x2_ASAP7_75t_L g5403 ( 
.A(n_5298),
.B(n_4652),
.Y(n_5403)
);

OAI22xp5_ASAP7_75t_L g5404 ( 
.A1(n_5226),
.A2(n_4722),
.B1(n_4716),
.B2(n_4671),
.Y(n_5404)
);

INVx2_ASAP7_75t_L g5405 ( 
.A(n_5032),
.Y(n_5405)
);

OAI21x1_ASAP7_75t_L g5406 ( 
.A1(n_4873),
.A2(n_4716),
.B(n_4671),
.Y(n_5406)
);

INVx2_ASAP7_75t_L g5407 ( 
.A(n_5049),
.Y(n_5407)
);

INVx2_ASAP7_75t_L g5408 ( 
.A(n_5063),
.Y(n_5408)
);

HB1xp67_ASAP7_75t_L g5409 ( 
.A(n_5177),
.Y(n_5409)
);

AOI22xp33_ASAP7_75t_L g5410 ( 
.A1(n_5247),
.A2(n_4716),
.B1(n_4722),
.B2(n_4671),
.Y(n_5410)
);

OAI21x1_ASAP7_75t_L g5411 ( 
.A1(n_5077),
.A2(n_4722),
.B(n_943),
.Y(n_5411)
);

AOI21xp5_ASAP7_75t_L g5412 ( 
.A1(n_4880),
.A2(n_943),
.B(n_942),
.Y(n_5412)
);

BUFx3_ASAP7_75t_L g5413 ( 
.A(n_4892),
.Y(n_5413)
);

OAI21x1_ASAP7_75t_L g5414 ( 
.A1(n_4950),
.A2(n_5141),
.B(n_4888),
.Y(n_5414)
);

INVx2_ASAP7_75t_L g5415 ( 
.A(n_5093),
.Y(n_5415)
);

AO21x2_ASAP7_75t_L g5416 ( 
.A1(n_5021),
.A2(n_945),
.B(n_944),
.Y(n_5416)
);

INVx1_ASAP7_75t_L g5417 ( 
.A(n_5008),
.Y(n_5417)
);

OAI21x1_ASAP7_75t_L g5418 ( 
.A1(n_5052),
.A2(n_5055),
.B(n_4938),
.Y(n_5418)
);

HB1xp67_ASAP7_75t_L g5419 ( 
.A(n_5159),
.Y(n_5419)
);

NAND2xp5_ASAP7_75t_L g5420 ( 
.A(n_5144),
.B(n_944),
.Y(n_5420)
);

OAI21x1_ASAP7_75t_SL g5421 ( 
.A1(n_4918),
.A2(n_946),
.B(n_945),
.Y(n_5421)
);

INVx1_ASAP7_75t_L g5422 ( 
.A(n_5026),
.Y(n_5422)
);

OAI21x1_ASAP7_75t_SL g5423 ( 
.A1(n_5020),
.A2(n_946),
.B(n_945),
.Y(n_5423)
);

OAI21x1_ASAP7_75t_SL g5424 ( 
.A1(n_4881),
.A2(n_5341),
.B(n_5281),
.Y(n_5424)
);

INVx2_ASAP7_75t_L g5425 ( 
.A(n_5064),
.Y(n_5425)
);

NAND2xp33_ASAP7_75t_R g5426 ( 
.A(n_5066),
.B(n_5084),
.Y(n_5426)
);

OAI21x1_ASAP7_75t_L g5427 ( 
.A1(n_5223),
.A2(n_948),
.B(n_947),
.Y(n_5427)
);

NAND3x1_ASAP7_75t_L g5428 ( 
.A(n_5258),
.B(n_949),
.C(n_947),
.Y(n_5428)
);

AOI22xp33_ASAP7_75t_SL g5429 ( 
.A1(n_4937),
.A2(n_949),
.B1(n_950),
.B2(n_947),
.Y(n_5429)
);

AOI21xp5_ASAP7_75t_L g5430 ( 
.A1(n_5004),
.A2(n_951),
.B(n_950),
.Y(n_5430)
);

XOR2xp5_ASAP7_75t_L g5431 ( 
.A(n_4929),
.B(n_57),
.Y(n_5431)
);

BUFx2_ASAP7_75t_SL g5432 ( 
.A(n_5023),
.Y(n_5432)
);

AOI21x1_ASAP7_75t_L g5433 ( 
.A1(n_4993),
.A2(n_5174),
.B(n_4945),
.Y(n_5433)
);

INVx2_ASAP7_75t_L g5434 ( 
.A(n_5072),
.Y(n_5434)
);

OAI21x1_ASAP7_75t_L g5435 ( 
.A1(n_4944),
.A2(n_951),
.B(n_950),
.Y(n_5435)
);

OAI21x1_ASAP7_75t_L g5436 ( 
.A1(n_4907),
.A2(n_953),
.B(n_952),
.Y(n_5436)
);

INVx1_ASAP7_75t_L g5437 ( 
.A(n_5094),
.Y(n_5437)
);

AND2x4_ASAP7_75t_L g5438 ( 
.A(n_5031),
.B(n_5110),
.Y(n_5438)
);

BUFx6f_ASAP7_75t_L g5439 ( 
.A(n_4895),
.Y(n_5439)
);

INVx2_ASAP7_75t_L g5440 ( 
.A(n_4948),
.Y(n_5440)
);

INVx1_ASAP7_75t_L g5441 ( 
.A(n_5197),
.Y(n_5441)
);

OAI21xp5_ASAP7_75t_L g5442 ( 
.A1(n_5179),
.A2(n_954),
.B(n_953),
.Y(n_5442)
);

OR2x2_ASAP7_75t_L g5443 ( 
.A(n_5097),
.B(n_1164),
.Y(n_5443)
);

NOR2xp33_ASAP7_75t_SL g5444 ( 
.A(n_5087),
.B(n_954),
.Y(n_5444)
);

AND2x4_ASAP7_75t_L g5445 ( 
.A(n_5237),
.B(n_954),
.Y(n_5445)
);

CKINVDCx20_ASAP7_75t_R g5446 ( 
.A(n_4887),
.Y(n_5446)
);

BUFx2_ASAP7_75t_L g5447 ( 
.A(n_5286),
.Y(n_5447)
);

INVx2_ASAP7_75t_L g5448 ( 
.A(n_4948),
.Y(n_5448)
);

A2O1A1Ixp33_ASAP7_75t_L g5449 ( 
.A1(n_5120),
.A2(n_956),
.B(n_957),
.C(n_955),
.Y(n_5449)
);

OAI221xp5_ASAP7_75t_L g5450 ( 
.A1(n_5123),
.A2(n_957),
.B1(n_958),
.B2(n_956),
.C(n_955),
.Y(n_5450)
);

AO31x2_ASAP7_75t_L g5451 ( 
.A1(n_5251),
.A2(n_956),
.A3(n_958),
.B(n_955),
.Y(n_5451)
);

OAI21x1_ASAP7_75t_L g5452 ( 
.A1(n_4877),
.A2(n_4979),
.B(n_4968),
.Y(n_5452)
);

BUFx6f_ASAP7_75t_L g5453 ( 
.A(n_4895),
.Y(n_5453)
);

INVx2_ASAP7_75t_L g5454 ( 
.A(n_5303),
.Y(n_5454)
);

BUFx6f_ASAP7_75t_L g5455 ( 
.A(n_4875),
.Y(n_5455)
);

INVx1_ASAP7_75t_L g5456 ( 
.A(n_5145),
.Y(n_5456)
);

AND2x2_ASAP7_75t_SL g5457 ( 
.A(n_5148),
.B(n_958),
.Y(n_5457)
);

O2A1O1Ixp33_ASAP7_75t_L g5458 ( 
.A1(n_4972),
.A2(n_960),
.B(n_961),
.C(n_959),
.Y(n_5458)
);

OAI21x1_ASAP7_75t_L g5459 ( 
.A1(n_4960),
.A2(n_960),
.B(n_959),
.Y(n_5459)
);

OAI21x1_ASAP7_75t_L g5460 ( 
.A1(n_4961),
.A2(n_960),
.B(n_959),
.Y(n_5460)
);

O2A1O1Ixp33_ASAP7_75t_L g5461 ( 
.A1(n_4906),
.A2(n_962),
.B(n_963),
.C(n_961),
.Y(n_5461)
);

OAI22xp5_ASAP7_75t_L g5462 ( 
.A1(n_5205),
.A2(n_962),
.B1(n_963),
.B2(n_961),
.Y(n_5462)
);

CKINVDCx11_ASAP7_75t_R g5463 ( 
.A(n_4878),
.Y(n_5463)
);

OAI22xp5_ASAP7_75t_L g5464 ( 
.A1(n_5205),
.A2(n_965),
.B1(n_966),
.B2(n_964),
.Y(n_5464)
);

BUFx2_ASAP7_75t_L g5465 ( 
.A(n_5248),
.Y(n_5465)
);

INVx1_ASAP7_75t_L g5466 ( 
.A(n_5170),
.Y(n_5466)
);

OA21x2_ASAP7_75t_L g5467 ( 
.A1(n_4988),
.A2(n_965),
.B(n_964),
.Y(n_5467)
);

CKINVDCx11_ASAP7_75t_R g5468 ( 
.A(n_4959),
.Y(n_5468)
);

NOR2xp33_ASAP7_75t_L g5469 ( 
.A(n_5012),
.B(n_58),
.Y(n_5469)
);

INVx2_ASAP7_75t_SL g5470 ( 
.A(n_4925),
.Y(n_5470)
);

NAND2x1p5_ASAP7_75t_L g5471 ( 
.A(n_4925),
.B(n_964),
.Y(n_5471)
);

O2A1O1Ixp33_ASAP7_75t_SL g5472 ( 
.A1(n_5000),
.A2(n_4982),
.B(n_4930),
.C(n_5256),
.Y(n_5472)
);

OA21x2_ASAP7_75t_L g5473 ( 
.A1(n_5272),
.A2(n_966),
.B(n_965),
.Y(n_5473)
);

INVx2_ASAP7_75t_L g5474 ( 
.A(n_5305),
.Y(n_5474)
);

BUFx3_ASAP7_75t_L g5475 ( 
.A(n_4939),
.Y(n_5475)
);

INVx2_ASAP7_75t_L g5476 ( 
.A(n_5319),
.Y(n_5476)
);

OAI21x1_ASAP7_75t_L g5477 ( 
.A1(n_5036),
.A2(n_968),
.B(n_967),
.Y(n_5477)
);

AND2x4_ASAP7_75t_L g5478 ( 
.A(n_5147),
.B(n_967),
.Y(n_5478)
);

OAI22xp5_ASAP7_75t_L g5479 ( 
.A1(n_5102),
.A2(n_968),
.B1(n_969),
.B2(n_967),
.Y(n_5479)
);

OAI21x1_ASAP7_75t_L g5480 ( 
.A1(n_5054),
.A2(n_5339),
.B(n_4978),
.Y(n_5480)
);

BUFx2_ASAP7_75t_L g5481 ( 
.A(n_5248),
.Y(n_5481)
);

NAND2xp5_ASAP7_75t_L g5482 ( 
.A(n_5168),
.B(n_1160),
.Y(n_5482)
);

BUFx10_ASAP7_75t_L g5483 ( 
.A(n_4939),
.Y(n_5483)
);

OAI21x1_ASAP7_75t_L g5484 ( 
.A1(n_5173),
.A2(n_970),
.B(n_969),
.Y(n_5484)
);

OAI21x1_ASAP7_75t_L g5485 ( 
.A1(n_4957),
.A2(n_971),
.B(n_970),
.Y(n_5485)
);

O2A1O1Ixp33_ASAP7_75t_SL g5486 ( 
.A1(n_4964),
.A2(n_971),
.B(n_972),
.C(n_970),
.Y(n_5486)
);

INVx1_ASAP7_75t_L g5487 ( 
.A(n_4974),
.Y(n_5487)
);

AO21x2_ASAP7_75t_L g5488 ( 
.A1(n_5022),
.A2(n_5043),
.B(n_4965),
.Y(n_5488)
);

AOI21xp33_ASAP7_75t_L g5489 ( 
.A1(n_5264),
.A2(n_972),
.B(n_971),
.Y(n_5489)
);

INVx1_ASAP7_75t_L g5490 ( 
.A(n_4986),
.Y(n_5490)
);

OAI21x1_ASAP7_75t_L g5491 ( 
.A1(n_4883),
.A2(n_973),
.B(n_972),
.Y(n_5491)
);

AOI222xp33_ASAP7_75t_L g5492 ( 
.A1(n_5216),
.A2(n_976),
.B1(n_974),
.B2(n_977),
.C1(n_975),
.C2(n_973),
.Y(n_5492)
);

AOI221xp5_ASAP7_75t_L g5493 ( 
.A1(n_5069),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.C(n_61),
.Y(n_5493)
);

AND2x2_ASAP7_75t_L g5494 ( 
.A(n_4928),
.B(n_59),
.Y(n_5494)
);

OAI21x1_ASAP7_75t_L g5495 ( 
.A1(n_5222),
.A2(n_974),
.B(n_973),
.Y(n_5495)
);

OAI22xp5_ASAP7_75t_SL g5496 ( 
.A1(n_5292),
.A2(n_975),
.B1(n_976),
.B2(n_974),
.Y(n_5496)
);

AO21x2_ASAP7_75t_L g5497 ( 
.A1(n_5285),
.A2(n_976),
.B(n_975),
.Y(n_5497)
);

BUFx2_ASAP7_75t_R g5498 ( 
.A(n_4952),
.Y(n_5498)
);

OAI21x1_ASAP7_75t_L g5499 ( 
.A1(n_5253),
.A2(n_4992),
.B(n_5080),
.Y(n_5499)
);

OAI21xp5_ASAP7_75t_L g5500 ( 
.A1(n_4920),
.A2(n_978),
.B(n_977),
.Y(n_5500)
);

INVx2_ASAP7_75t_L g5501 ( 
.A(n_4932),
.Y(n_5501)
);

CKINVDCx16_ASAP7_75t_R g5502 ( 
.A(n_5070),
.Y(n_5502)
);

AND2x2_ASAP7_75t_L g5503 ( 
.A(n_5006),
.B(n_60),
.Y(n_5503)
);

OAI21x1_ASAP7_75t_L g5504 ( 
.A1(n_4889),
.A2(n_978),
.B(n_977),
.Y(n_5504)
);

INVx1_ASAP7_75t_L g5505 ( 
.A(n_5306),
.Y(n_5505)
);

AND2x4_ASAP7_75t_L g5506 ( 
.A(n_5236),
.B(n_978),
.Y(n_5506)
);

INVx1_ASAP7_75t_SL g5507 ( 
.A(n_5155),
.Y(n_5507)
);

BUFx8_ASAP7_75t_L g5508 ( 
.A(n_5130),
.Y(n_5508)
);

NAND2x1p5_ASAP7_75t_L g5509 ( 
.A(n_4875),
.B(n_979),
.Y(n_5509)
);

OA21x2_ASAP7_75t_L g5510 ( 
.A1(n_4876),
.A2(n_980),
.B(n_979),
.Y(n_5510)
);

INVx5_ASAP7_75t_L g5511 ( 
.A(n_5191),
.Y(n_5511)
);

INVx1_ASAP7_75t_L g5512 ( 
.A(n_5133),
.Y(n_5512)
);

OAI21x1_ASAP7_75t_L g5513 ( 
.A1(n_5284),
.A2(n_981),
.B(n_980),
.Y(n_5513)
);

OAI21x1_ASAP7_75t_L g5514 ( 
.A1(n_5038),
.A2(n_5323),
.B(n_5092),
.Y(n_5514)
);

INVx4_ASAP7_75t_L g5515 ( 
.A(n_4955),
.Y(n_5515)
);

INVx1_ASAP7_75t_L g5516 ( 
.A(n_4933),
.Y(n_5516)
);

OA21x2_ASAP7_75t_L g5517 ( 
.A1(n_4890),
.A2(n_982),
.B(n_981),
.Y(n_5517)
);

NAND2xp5_ASAP7_75t_L g5518 ( 
.A(n_5176),
.B(n_981),
.Y(n_5518)
);

OAI21xp5_ASAP7_75t_L g5519 ( 
.A1(n_5081),
.A2(n_983),
.B(n_982),
.Y(n_5519)
);

NOR2x1_ASAP7_75t_SL g5520 ( 
.A(n_4937),
.B(n_982),
.Y(n_5520)
);

BUFx6f_ASAP7_75t_L g5521 ( 
.A(n_5191),
.Y(n_5521)
);

AO21x2_ASAP7_75t_L g5522 ( 
.A1(n_5018),
.A2(n_984),
.B(n_983),
.Y(n_5522)
);

INVx2_ASAP7_75t_L g5523 ( 
.A(n_4932),
.Y(n_5523)
);

INVx3_ASAP7_75t_L g5524 ( 
.A(n_5246),
.Y(n_5524)
);

OAI21x1_ASAP7_75t_L g5525 ( 
.A1(n_5051),
.A2(n_985),
.B(n_983),
.Y(n_5525)
);

INVx2_ASAP7_75t_L g5526 ( 
.A(n_5318),
.Y(n_5526)
);

CKINVDCx11_ASAP7_75t_R g5527 ( 
.A(n_4911),
.Y(n_5527)
);

OAI21x1_ASAP7_75t_SL g5528 ( 
.A1(n_5158),
.A2(n_986),
.B(n_985),
.Y(n_5528)
);

INVx1_ASAP7_75t_L g5529 ( 
.A(n_4936),
.Y(n_5529)
);

OA21x2_ASAP7_75t_L g5530 ( 
.A1(n_4931),
.A2(n_987),
.B(n_986),
.Y(n_5530)
);

OAI22xp5_ASAP7_75t_L g5531 ( 
.A1(n_4937),
.A2(n_987),
.B1(n_988),
.B2(n_986),
.Y(n_5531)
);

OAI22xp5_ASAP7_75t_L g5532 ( 
.A1(n_5075),
.A2(n_989),
.B1(n_990),
.B2(n_988),
.Y(n_5532)
);

BUFx8_ASAP7_75t_SL g5533 ( 
.A(n_4990),
.Y(n_5533)
);

INVx2_ASAP7_75t_L g5534 ( 
.A(n_4993),
.Y(n_5534)
);

AO31x2_ASAP7_75t_L g5535 ( 
.A1(n_5231),
.A2(n_990),
.A3(n_991),
.B(n_989),
.Y(n_5535)
);

AOI22xp33_ASAP7_75t_SL g5536 ( 
.A1(n_4885),
.A2(n_990),
.B1(n_992),
.B2(n_989),
.Y(n_5536)
);

BUFx3_ASAP7_75t_L g5537 ( 
.A(n_5107),
.Y(n_5537)
);

OAI22xp5_ASAP7_75t_L g5538 ( 
.A1(n_5099),
.A2(n_993),
.B1(n_994),
.B2(n_992),
.Y(n_5538)
);

INVx2_ASAP7_75t_SL g5539 ( 
.A(n_5091),
.Y(n_5539)
);

NOR2x1_ASAP7_75t_L g5540 ( 
.A(n_5034),
.B(n_993),
.Y(n_5540)
);

INVx2_ASAP7_75t_L g5541 ( 
.A(n_5079),
.Y(n_5541)
);

OA21x2_ASAP7_75t_L g5542 ( 
.A1(n_4983),
.A2(n_995),
.B(n_994),
.Y(n_5542)
);

AOI221xp5_ASAP7_75t_SL g5543 ( 
.A1(n_4946),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.C(n_63),
.Y(n_5543)
);

NAND2xp5_ASAP7_75t_SL g5544 ( 
.A(n_5079),
.B(n_996),
.Y(n_5544)
);

AOI21xp5_ASAP7_75t_L g5545 ( 
.A1(n_5058),
.A2(n_997),
.B(n_996),
.Y(n_5545)
);

OA21x2_ASAP7_75t_L g5546 ( 
.A1(n_5062),
.A2(n_998),
.B(n_997),
.Y(n_5546)
);

INVx1_ASAP7_75t_L g5547 ( 
.A(n_4949),
.Y(n_5547)
);

OAI21x1_ASAP7_75t_L g5548 ( 
.A1(n_5117),
.A2(n_998),
.B(n_997),
.Y(n_5548)
);

OAI22xp5_ASAP7_75t_L g5549 ( 
.A1(n_4935),
.A2(n_5277),
.B1(n_5335),
.B2(n_5344),
.Y(n_5549)
);

OAI21xp5_ASAP7_75t_L g5550 ( 
.A1(n_5106),
.A2(n_1000),
.B(n_999),
.Y(n_5550)
);

OR2x6_ASAP7_75t_L g5551 ( 
.A(n_4899),
.B(n_999),
.Y(n_5551)
);

OAI21x1_ASAP7_75t_L g5552 ( 
.A1(n_5194),
.A2(n_1000),
.B(n_999),
.Y(n_5552)
);

OAI21x1_ASAP7_75t_L g5553 ( 
.A1(n_5116),
.A2(n_1002),
.B(n_1001),
.Y(n_5553)
);

AND2x4_ASAP7_75t_L g5554 ( 
.A(n_5217),
.B(n_1001),
.Y(n_5554)
);

BUFx2_ASAP7_75t_L g5555 ( 
.A(n_5309),
.Y(n_5555)
);

INVx1_ASAP7_75t_L g5556 ( 
.A(n_4962),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_4967),
.Y(n_5557)
);

AOI22xp33_ASAP7_75t_L g5558 ( 
.A1(n_5249),
.A2(n_5210),
.B1(n_5338),
.B2(n_5327),
.Y(n_5558)
);

NAND3xp33_ASAP7_75t_L g5559 ( 
.A(n_4998),
.B(n_1002),
.C(n_1001),
.Y(n_5559)
);

INVx1_ASAP7_75t_L g5560 ( 
.A(n_4980),
.Y(n_5560)
);

INVx1_ASAP7_75t_L g5561 ( 
.A(n_5180),
.Y(n_5561)
);

INVx3_ASAP7_75t_L g5562 ( 
.A(n_5142),
.Y(n_5562)
);

HB1xp67_ASAP7_75t_L g5563 ( 
.A(n_5294),
.Y(n_5563)
);

AOI22xp33_ASAP7_75t_L g5564 ( 
.A1(n_5301),
.A2(n_1003),
.B1(n_1004),
.B2(n_1002),
.Y(n_5564)
);

AND2x4_ASAP7_75t_L g5565 ( 
.A(n_5088),
.B(n_1004),
.Y(n_5565)
);

AOI22xp33_ASAP7_75t_L g5566 ( 
.A1(n_5289),
.A2(n_1006),
.B1(n_1007),
.B2(n_1005),
.Y(n_5566)
);

OAI21x1_ASAP7_75t_L g5567 ( 
.A1(n_5073),
.A2(n_1006),
.B(n_1005),
.Y(n_5567)
);

CKINVDCx5p33_ASAP7_75t_R g5568 ( 
.A(n_5037),
.Y(n_5568)
);

AO21x2_ASAP7_75t_L g5569 ( 
.A1(n_4913),
.A2(n_1008),
.B(n_1007),
.Y(n_5569)
);

AOI22xp33_ASAP7_75t_SL g5570 ( 
.A1(n_5240),
.A2(n_1008),
.B1(n_1009),
.B2(n_1007),
.Y(n_5570)
);

OAI21x1_ASAP7_75t_L g5571 ( 
.A1(n_5201),
.A2(n_1009),
.B(n_1008),
.Y(n_5571)
);

INVx2_ASAP7_75t_SL g5572 ( 
.A(n_5142),
.Y(n_5572)
);

INVx2_ASAP7_75t_L g5573 ( 
.A(n_5342),
.Y(n_5573)
);

AO21x2_ASAP7_75t_L g5574 ( 
.A1(n_5095),
.A2(n_1010),
.B(n_1009),
.Y(n_5574)
);

INVx2_ASAP7_75t_L g5575 ( 
.A(n_5275),
.Y(n_5575)
);

OAI21x1_ASAP7_75t_L g5576 ( 
.A1(n_5214),
.A2(n_1011),
.B(n_1010),
.Y(n_5576)
);

AOI21xp5_ASAP7_75t_SL g5577 ( 
.A1(n_5041),
.A2(n_1012),
.B(n_1011),
.Y(n_5577)
);

INVx2_ASAP7_75t_L g5578 ( 
.A(n_5209),
.Y(n_5578)
);

OAI21x1_ASAP7_75t_L g5579 ( 
.A1(n_5263),
.A2(n_1012),
.B(n_1011),
.Y(n_5579)
);

OAI22xp5_ASAP7_75t_L g5580 ( 
.A1(n_5307),
.A2(n_1013),
.B1(n_1014),
.B2(n_1012),
.Y(n_5580)
);

AND2x4_ASAP7_75t_L g5581 ( 
.A(n_5295),
.B(n_1013),
.Y(n_5581)
);

INVx2_ASAP7_75t_L g5582 ( 
.A(n_5229),
.Y(n_5582)
);

INVxp67_ASAP7_75t_SL g5583 ( 
.A(n_5244),
.Y(n_5583)
);

NAND2xp33_ASAP7_75t_R g5584 ( 
.A(n_4916),
.B(n_4970),
.Y(n_5584)
);

INVx1_ASAP7_75t_L g5585 ( 
.A(n_5185),
.Y(n_5585)
);

INVx4_ASAP7_75t_L g5586 ( 
.A(n_5169),
.Y(n_5586)
);

INVx2_ASAP7_75t_SL g5587 ( 
.A(n_5167),
.Y(n_5587)
);

INVx1_ASAP7_75t_L g5588 ( 
.A(n_5207),
.Y(n_5588)
);

AND2x4_ASAP7_75t_L g5589 ( 
.A(n_5245),
.B(n_1013),
.Y(n_5589)
);

OAI21x1_ASAP7_75t_L g5590 ( 
.A1(n_5215),
.A2(n_1015),
.B(n_1014),
.Y(n_5590)
);

OAI21x1_ASAP7_75t_L g5591 ( 
.A1(n_4977),
.A2(n_1015),
.B(n_1014),
.Y(n_5591)
);

OAI22xp5_ASAP7_75t_L g5592 ( 
.A1(n_5307),
.A2(n_1017),
.B1(n_1018),
.B2(n_1016),
.Y(n_5592)
);

BUFx12f_ASAP7_75t_L g5593 ( 
.A(n_4999),
.Y(n_5593)
);

A2O1A1Ixp33_ASAP7_75t_L g5594 ( 
.A1(n_5282),
.A2(n_1017),
.B(n_1018),
.C(n_1016),
.Y(n_5594)
);

OAI21x1_ASAP7_75t_L g5595 ( 
.A1(n_5181),
.A2(n_1019),
.B(n_1017),
.Y(n_5595)
);

INVx2_ASAP7_75t_L g5596 ( 
.A(n_5250),
.Y(n_5596)
);

OAI21xp5_ASAP7_75t_L g5597 ( 
.A1(n_5025),
.A2(n_1020),
.B(n_1019),
.Y(n_5597)
);

INVx2_ASAP7_75t_L g5598 ( 
.A(n_5250),
.Y(n_5598)
);

AO21x2_ASAP7_75t_L g5599 ( 
.A1(n_5260),
.A2(n_1021),
.B(n_1020),
.Y(n_5599)
);

A2O1A1Ixp33_ASAP7_75t_L g5600 ( 
.A1(n_4917),
.A2(n_1022),
.B(n_1023),
.C(n_1020),
.Y(n_5600)
);

BUFx2_ASAP7_75t_L g5601 ( 
.A(n_5250),
.Y(n_5601)
);

OAI21x1_ASAP7_75t_L g5602 ( 
.A1(n_4872),
.A2(n_1023),
.B(n_1022),
.Y(n_5602)
);

NOR2xp33_ASAP7_75t_L g5603 ( 
.A(n_4971),
.B(n_61),
.Y(n_5603)
);

OAI21xp5_ASAP7_75t_L g5604 ( 
.A1(n_5035),
.A2(n_1025),
.B(n_1024),
.Y(n_5604)
);

OAI22xp5_ASAP7_75t_L g5605 ( 
.A1(n_5083),
.A2(n_1025),
.B1(n_1026),
.B2(n_1024),
.Y(n_5605)
);

INVx1_ASAP7_75t_L g5606 ( 
.A(n_5134),
.Y(n_5606)
);

OAI21x1_ASAP7_75t_SL g5607 ( 
.A1(n_5061),
.A2(n_5330),
.B(n_5325),
.Y(n_5607)
);

AO32x2_ASAP7_75t_L g5608 ( 
.A1(n_5103),
.A2(n_1028),
.A3(n_1029),
.B1(n_1027),
.B2(n_1024),
.Y(n_5608)
);

OAI21xp5_ASAP7_75t_L g5609 ( 
.A1(n_5257),
.A2(n_1029),
.B(n_1027),
.Y(n_5609)
);

OA21x2_ASAP7_75t_L g5610 ( 
.A1(n_4904),
.A2(n_1030),
.B(n_1029),
.Y(n_5610)
);

AOI221xp5_ASAP7_75t_L g5611 ( 
.A1(n_4896),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.C(n_64),
.Y(n_5611)
);

AOI22xp33_ASAP7_75t_L g5612 ( 
.A1(n_5266),
.A2(n_1031),
.B1(n_1032),
.B2(n_1030),
.Y(n_5612)
);

INVx1_ASAP7_75t_L g5613 ( 
.A(n_5111),
.Y(n_5613)
);

INVx1_ASAP7_75t_SL g5614 ( 
.A(n_5153),
.Y(n_5614)
);

NAND2xp5_ASAP7_75t_L g5615 ( 
.A(n_5320),
.B(n_1030),
.Y(n_5615)
);

INVx1_ASAP7_75t_L g5616 ( 
.A(n_4989),
.Y(n_5616)
);

INVx1_ASAP7_75t_L g5617 ( 
.A(n_4991),
.Y(n_5617)
);

INVx1_ASAP7_75t_L g5618 ( 
.A(n_4996),
.Y(n_5618)
);

OAI21x1_ASAP7_75t_L g5619 ( 
.A1(n_5313),
.A2(n_1032),
.B(n_1031),
.Y(n_5619)
);

OAI21x1_ASAP7_75t_L g5620 ( 
.A1(n_5316),
.A2(n_1033),
.B(n_1032),
.Y(n_5620)
);

OAI21x1_ASAP7_75t_L g5621 ( 
.A1(n_5218),
.A2(n_1034),
.B(n_1033),
.Y(n_5621)
);

INVx1_ASAP7_75t_L g5622 ( 
.A(n_5001),
.Y(n_5622)
);

OAI21x1_ASAP7_75t_L g5623 ( 
.A1(n_5219),
.A2(n_1035),
.B(n_1034),
.Y(n_5623)
);

INVx1_ASAP7_75t_SL g5624 ( 
.A(n_5033),
.Y(n_5624)
);

INVx2_ASAP7_75t_SL g5625 ( 
.A(n_5065),
.Y(n_5625)
);

INVx2_ASAP7_75t_L g5626 ( 
.A(n_5345),
.Y(n_5626)
);

OAI21x1_ASAP7_75t_L g5627 ( 
.A1(n_5127),
.A2(n_1035),
.B(n_1034),
.Y(n_5627)
);

OAI21x1_ASAP7_75t_L g5628 ( 
.A1(n_5089),
.A2(n_5227),
.B(n_5104),
.Y(n_5628)
);

INVx2_ASAP7_75t_L g5629 ( 
.A(n_5100),
.Y(n_5629)
);

OAI21x1_ASAP7_75t_L g5630 ( 
.A1(n_5324),
.A2(n_1037),
.B(n_1036),
.Y(n_5630)
);

INVx2_ASAP7_75t_SL g5631 ( 
.A(n_5225),
.Y(n_5631)
);

AOI22xp33_ASAP7_75t_L g5632 ( 
.A1(n_5333),
.A2(n_1037),
.B1(n_1038),
.B2(n_1036),
.Y(n_5632)
);

OAI21xp5_ASAP7_75t_L g5633 ( 
.A1(n_5010),
.A2(n_1037),
.B(n_1036),
.Y(n_5633)
);

BUFx2_ASAP7_75t_SL g5634 ( 
.A(n_5129),
.Y(n_5634)
);

INVx1_ASAP7_75t_L g5635 ( 
.A(n_4886),
.Y(n_5635)
);

INVx1_ASAP7_75t_L g5636 ( 
.A(n_5011),
.Y(n_5636)
);

INVx1_ASAP7_75t_L g5637 ( 
.A(n_5017),
.Y(n_5637)
);

AO21x2_ASAP7_75t_L g5638 ( 
.A1(n_5269),
.A2(n_1039),
.B(n_1038),
.Y(n_5638)
);

AND2x4_ASAP7_75t_L g5639 ( 
.A(n_5190),
.B(n_1039),
.Y(n_5639)
);

OR2x6_ASAP7_75t_L g5640 ( 
.A(n_5208),
.B(n_1039),
.Y(n_5640)
);

OAI21x1_ASAP7_75t_L g5641 ( 
.A1(n_5175),
.A2(n_1041),
.B(n_1040),
.Y(n_5641)
);

BUFx3_ASAP7_75t_L g5642 ( 
.A(n_5233),
.Y(n_5642)
);

OAI21x1_ASAP7_75t_L g5643 ( 
.A1(n_5184),
.A2(n_1041),
.B(n_1040),
.Y(n_5643)
);

AO21x2_ASAP7_75t_L g5644 ( 
.A1(n_5149),
.A2(n_1041),
.B(n_1040),
.Y(n_5644)
);

BUFx2_ASAP7_75t_L g5645 ( 
.A(n_5172),
.Y(n_5645)
);

OAI21x1_ASAP7_75t_L g5646 ( 
.A1(n_5322),
.A2(n_1043),
.B(n_1042),
.Y(n_5646)
);

AND2x4_ASAP7_75t_L g5647 ( 
.A(n_5165),
.B(n_1042),
.Y(n_5647)
);

OA21x2_ASAP7_75t_L g5648 ( 
.A1(n_4912),
.A2(n_1043),
.B(n_1042),
.Y(n_5648)
);

NOR2xp33_ASAP7_75t_L g5649 ( 
.A(n_5162),
.B(n_63),
.Y(n_5649)
);

OAI21x1_ASAP7_75t_L g5650 ( 
.A1(n_5058),
.A2(n_1044),
.B(n_1043),
.Y(n_5650)
);

AOI22xp33_ASAP7_75t_L g5651 ( 
.A1(n_4909),
.A2(n_1045),
.B1(n_1046),
.B2(n_1044),
.Y(n_5651)
);

OAI21x1_ASAP7_75t_L g5652 ( 
.A1(n_5014),
.A2(n_1045),
.B(n_1044),
.Y(n_5652)
);

OAI22xp5_ASAP7_75t_L g5653 ( 
.A1(n_5071),
.A2(n_1046),
.B1(n_1047),
.B2(n_1045),
.Y(n_5653)
);

INVx1_ASAP7_75t_L g5654 ( 
.A(n_5028),
.Y(n_5654)
);

AND2x4_ASAP7_75t_L g5655 ( 
.A(n_4985),
.B(n_1047),
.Y(n_5655)
);

INVx3_ASAP7_75t_L g5656 ( 
.A(n_5270),
.Y(n_5656)
);

OAI21x1_ASAP7_75t_L g5657 ( 
.A1(n_5336),
.A2(n_1048),
.B(n_1047),
.Y(n_5657)
);

OAI21x1_ASAP7_75t_L g5658 ( 
.A1(n_5198),
.A2(n_1049),
.B(n_1048),
.Y(n_5658)
);

NAND2x1p5_ASAP7_75t_L g5659 ( 
.A(n_4915),
.B(n_1049),
.Y(n_5659)
);

OAI21x1_ASAP7_75t_L g5660 ( 
.A1(n_5042),
.A2(n_1050),
.B(n_1049),
.Y(n_5660)
);

AOI21xp5_ASAP7_75t_L g5661 ( 
.A1(n_5161),
.A2(n_1051),
.B(n_1050),
.Y(n_5661)
);

OR2x2_ASAP7_75t_L g5662 ( 
.A(n_5466),
.B(n_5409),
.Y(n_5662)
);

NAND2xp5_ASAP7_75t_L g5663 ( 
.A(n_5399),
.B(n_5310),
.Y(n_5663)
);

OA21x2_ASAP7_75t_L g5664 ( 
.A1(n_5354),
.A2(n_5271),
.B(n_5304),
.Y(n_5664)
);

INVx1_ASAP7_75t_L g5665 ( 
.A(n_5346),
.Y(n_5665)
);

NAND2xp5_ASAP7_75t_L g5666 ( 
.A(n_5400),
.B(n_5314),
.Y(n_5666)
);

OAI21x1_ASAP7_75t_L g5667 ( 
.A1(n_5406),
.A2(n_5015),
.B(n_4994),
.Y(n_5667)
);

OAI21x1_ASAP7_75t_L g5668 ( 
.A1(n_5433),
.A2(n_5278),
.B(n_5115),
.Y(n_5668)
);

INVx1_ASAP7_75t_L g5669 ( 
.A(n_5352),
.Y(n_5669)
);

NAND2xp5_ASAP7_75t_L g5670 ( 
.A(n_5578),
.B(n_5262),
.Y(n_5670)
);

OAI21x1_ASAP7_75t_L g5671 ( 
.A1(n_5514),
.A2(n_5122),
.B(n_5112),
.Y(n_5671)
);

INVx2_ASAP7_75t_L g5672 ( 
.A(n_5447),
.Y(n_5672)
);

BUFx2_ASAP7_75t_L g5673 ( 
.A(n_5354),
.Y(n_5673)
);

INVx2_ASAP7_75t_SL g5674 ( 
.A(n_5483),
.Y(n_5674)
);

OAI21x1_ASAP7_75t_L g5675 ( 
.A1(n_5452),
.A2(n_5138),
.B(n_5131),
.Y(n_5675)
);

INVx1_ASAP7_75t_L g5676 ( 
.A(n_5358),
.Y(n_5676)
);

NAND2xp5_ASAP7_75t_L g5677 ( 
.A(n_5582),
.B(n_5186),
.Y(n_5677)
);

INVx1_ASAP7_75t_L g5678 ( 
.A(n_5362),
.Y(n_5678)
);

AOI21xp5_ASAP7_75t_L g5679 ( 
.A1(n_5404),
.A2(n_5369),
.B(n_5366),
.Y(n_5679)
);

INVx1_ASAP7_75t_L g5680 ( 
.A(n_5364),
.Y(n_5680)
);

INVx1_ASAP7_75t_L g5681 ( 
.A(n_5384),
.Y(n_5681)
);

INVx2_ASAP7_75t_L g5682 ( 
.A(n_5447),
.Y(n_5682)
);

INVx4_ASAP7_75t_SL g5683 ( 
.A(n_5387),
.Y(n_5683)
);

OR2x2_ASAP7_75t_L g5684 ( 
.A(n_5419),
.B(n_4893),
.Y(n_5684)
);

NAND2xp5_ASAP7_75t_L g5685 ( 
.A(n_5561),
.B(n_4942),
.Y(n_5685)
);

OAI21xp5_ASAP7_75t_L g5686 ( 
.A1(n_5457),
.A2(n_4903),
.B(n_4943),
.Y(n_5686)
);

INVx1_ASAP7_75t_L g5687 ( 
.A(n_5391),
.Y(n_5687)
);

OAI21xp33_ASAP7_75t_SL g5688 ( 
.A1(n_5387),
.A2(n_5030),
.B(n_5154),
.Y(n_5688)
);

AO21x2_ASAP7_75t_L g5689 ( 
.A1(n_5424),
.A2(n_5047),
.B(n_5039),
.Y(n_5689)
);

AO31x2_ASAP7_75t_L g5690 ( 
.A1(n_5645),
.A2(n_5534),
.A3(n_5448),
.B(n_5440),
.Y(n_5690)
);

AND2x4_ASAP7_75t_L g5691 ( 
.A(n_5382),
.B(n_5164),
.Y(n_5691)
);

AO31x2_ASAP7_75t_L g5692 ( 
.A1(n_5645),
.A2(n_4941),
.A3(n_5090),
.B(n_5212),
.Y(n_5692)
);

INVx1_ASAP7_75t_L g5693 ( 
.A(n_5401),
.Y(n_5693)
);

CKINVDCx11_ASAP7_75t_R g5694 ( 
.A(n_5446),
.Y(n_5694)
);

INVx2_ASAP7_75t_L g5695 ( 
.A(n_5378),
.Y(n_5695)
);

INVx2_ASAP7_75t_L g5696 ( 
.A(n_5385),
.Y(n_5696)
);

INVx1_ASAP7_75t_L g5697 ( 
.A(n_5417),
.Y(n_5697)
);

AOI21x1_ASAP7_75t_L g5698 ( 
.A1(n_5601),
.A2(n_5267),
.B(n_5196),
.Y(n_5698)
);

INVx1_ASAP7_75t_L g5699 ( 
.A(n_5422),
.Y(n_5699)
);

AOI21x1_ASAP7_75t_L g5700 ( 
.A1(n_5601),
.A2(n_5393),
.B(n_5355),
.Y(n_5700)
);

OR2x2_ASAP7_75t_L g5701 ( 
.A(n_5441),
.B(n_4897),
.Y(n_5701)
);

INVx2_ASAP7_75t_L g5702 ( 
.A(n_5395),
.Y(n_5702)
);

INVx1_ASAP7_75t_L g5703 ( 
.A(n_5585),
.Y(n_5703)
);

NOR2xp33_ASAP7_75t_L g5704 ( 
.A(n_5367),
.B(n_5199),
.Y(n_5704)
);

INVx1_ASAP7_75t_L g5705 ( 
.A(n_5588),
.Y(n_5705)
);

NAND2xp5_ASAP7_75t_SL g5706 ( 
.A(n_5507),
.B(n_5241),
.Y(n_5706)
);

INVx2_ASAP7_75t_L g5707 ( 
.A(n_5405),
.Y(n_5707)
);

INVx2_ASAP7_75t_L g5708 ( 
.A(n_5407),
.Y(n_5708)
);

INVx1_ASAP7_75t_L g5709 ( 
.A(n_5456),
.Y(n_5709)
);

INVx1_ASAP7_75t_L g5710 ( 
.A(n_5512),
.Y(n_5710)
);

AOI21xp5_ASAP7_75t_L g5711 ( 
.A1(n_5393),
.A2(n_4981),
.B(n_5157),
.Y(n_5711)
);

OAI21x1_ASAP7_75t_L g5712 ( 
.A1(n_5480),
.A2(n_5414),
.B(n_5499),
.Y(n_5712)
);

INVx1_ASAP7_75t_L g5713 ( 
.A(n_5437),
.Y(n_5713)
);

INVx2_ASAP7_75t_L g5714 ( 
.A(n_5408),
.Y(n_5714)
);

CKINVDCx20_ASAP7_75t_R g5715 ( 
.A(n_5463),
.Y(n_5715)
);

OAI21x1_ASAP7_75t_L g5716 ( 
.A1(n_5418),
.A2(n_4976),
.B(n_5009),
.Y(n_5716)
);

NAND2x1p5_ASAP7_75t_L g5717 ( 
.A(n_5524),
.B(n_5027),
.Y(n_5717)
);

AOI21xp5_ASAP7_75t_L g5718 ( 
.A1(n_5356),
.A2(n_5283),
.B(n_5096),
.Y(n_5718)
);

BUFx8_ASAP7_75t_L g5719 ( 
.A(n_5357),
.Y(n_5719)
);

OA21x2_ASAP7_75t_L g5720 ( 
.A1(n_5349),
.A2(n_5232),
.B(n_5059),
.Y(n_5720)
);

OAI21x1_ASAP7_75t_L g5721 ( 
.A1(n_5370),
.A2(n_5273),
.B(n_5057),
.Y(n_5721)
);

INVx2_ASAP7_75t_L g5722 ( 
.A(n_5415),
.Y(n_5722)
);

INVx1_ASAP7_75t_L g5723 ( 
.A(n_5425),
.Y(n_5723)
);

INVx1_ASAP7_75t_L g5724 ( 
.A(n_5434),
.Y(n_5724)
);

AO31x2_ASAP7_75t_L g5725 ( 
.A1(n_5501),
.A2(n_5204),
.A3(n_5317),
.B(n_5299),
.Y(n_5725)
);

NAND2xp5_ASAP7_75t_L g5726 ( 
.A(n_5487),
.B(n_5228),
.Y(n_5726)
);

OR2x2_ASAP7_75t_L g5727 ( 
.A(n_5350),
.B(n_5490),
.Y(n_5727)
);

INVx1_ASAP7_75t_L g5728 ( 
.A(n_5505),
.Y(n_5728)
);

NAND2xp5_ASAP7_75t_L g5729 ( 
.A(n_5613),
.B(n_4901),
.Y(n_5729)
);

AND2x4_ASAP7_75t_L g5730 ( 
.A(n_5555),
.B(n_5013),
.Y(n_5730)
);

INVx1_ASAP7_75t_L g5731 ( 
.A(n_5606),
.Y(n_5731)
);

AND2x2_ASAP7_75t_L g5732 ( 
.A(n_5359),
.B(n_5137),
.Y(n_5732)
);

AOI21xp5_ASAP7_75t_L g5733 ( 
.A1(n_5356),
.A2(n_5332),
.B(n_5040),
.Y(n_5733)
);

NAND2xp5_ASAP7_75t_SL g5734 ( 
.A(n_5555),
.B(n_5438),
.Y(n_5734)
);

AOI22xp5_ASAP7_75t_L g5735 ( 
.A1(n_5426),
.A2(n_4908),
.B1(n_5056),
.B2(n_5124),
.Y(n_5735)
);

BUFx3_ASAP7_75t_L g5736 ( 
.A(n_5413),
.Y(n_5736)
);

OA21x2_ASAP7_75t_L g5737 ( 
.A1(n_5523),
.A2(n_5105),
.B(n_5053),
.Y(n_5737)
);

OAI21x1_ASAP7_75t_L g5738 ( 
.A1(n_5353),
.A2(n_5143),
.B(n_4951),
.Y(n_5738)
);

AO21x2_ASAP7_75t_L g5739 ( 
.A1(n_5423),
.A2(n_5121),
.B(n_5113),
.Y(n_5739)
);

AOI21xp5_ASAP7_75t_L g5740 ( 
.A1(n_5577),
.A2(n_5486),
.B(n_5510),
.Y(n_5740)
);

AO31x2_ASAP7_75t_L g5741 ( 
.A1(n_5465),
.A2(n_5481),
.A3(n_5549),
.B(n_5541),
.Y(n_5741)
);

AOI22x1_ASAP7_75t_L g5742 ( 
.A1(n_5502),
.A2(n_5195),
.B1(n_4924),
.B2(n_5098),
.Y(n_5742)
);

BUFx3_ASAP7_75t_L g5743 ( 
.A(n_5475),
.Y(n_5743)
);

INVx4_ASAP7_75t_L g5744 ( 
.A(n_5586),
.Y(n_5744)
);

AO21x2_ASAP7_75t_L g5745 ( 
.A1(n_5361),
.A2(n_5128),
.B(n_5151),
.Y(n_5745)
);

OA21x2_ASAP7_75t_L g5746 ( 
.A1(n_5583),
.A2(n_5178),
.B(n_5224),
.Y(n_5746)
);

AO31x2_ASAP7_75t_L g5747 ( 
.A1(n_5465),
.A2(n_5254),
.A3(n_5252),
.B(n_5288),
.Y(n_5747)
);

NAND2xp5_ASAP7_75t_L g5748 ( 
.A(n_5516),
.B(n_5150),
.Y(n_5748)
);

INVx1_ASAP7_75t_L g5749 ( 
.A(n_5454),
.Y(n_5749)
);

AOI21x1_ASAP7_75t_L g5750 ( 
.A1(n_5563),
.A2(n_5085),
.B(n_5163),
.Y(n_5750)
);

OAI21x1_ASAP7_75t_SL g5751 ( 
.A1(n_5520),
.A2(n_5060),
.B(n_5136),
.Y(n_5751)
);

INVx1_ASAP7_75t_L g5752 ( 
.A(n_5474),
.Y(n_5752)
);

NAND2xp5_ASAP7_75t_SL g5753 ( 
.A(n_5511),
.B(n_5166),
.Y(n_5753)
);

AOI21xp5_ASAP7_75t_L g5754 ( 
.A1(n_5510),
.A2(n_5287),
.B(n_5279),
.Y(n_5754)
);

AO21x2_ASAP7_75t_L g5755 ( 
.A1(n_5376),
.A2(n_4894),
.B(n_5206),
.Y(n_5755)
);

INVx1_ASAP7_75t_L g5756 ( 
.A(n_5476),
.Y(n_5756)
);

OAI21x1_ASAP7_75t_L g5757 ( 
.A1(n_5347),
.A2(n_5380),
.B(n_5427),
.Y(n_5757)
);

BUFx6f_ASAP7_75t_L g5758 ( 
.A(n_5521),
.Y(n_5758)
);

INVx1_ASAP7_75t_L g5759 ( 
.A(n_5392),
.Y(n_5759)
);

INVx2_ASAP7_75t_L g5760 ( 
.A(n_5526),
.Y(n_5760)
);

CKINVDCx20_ASAP7_75t_R g5761 ( 
.A(n_5468),
.Y(n_5761)
);

NAND2x1_ASAP7_75t_L g5762 ( 
.A(n_5515),
.B(n_5085),
.Y(n_5762)
);

BUFx8_ASAP7_75t_L g5763 ( 
.A(n_5455),
.Y(n_5763)
);

OAI21x1_ASAP7_75t_SL g5764 ( 
.A1(n_5397),
.A2(n_5230),
.B(n_5125),
.Y(n_5764)
);

AOI21xp5_ASAP7_75t_L g5765 ( 
.A1(n_5412),
.A2(n_5132),
.B(n_5048),
.Y(n_5765)
);

INVx1_ASAP7_75t_L g5766 ( 
.A(n_5386),
.Y(n_5766)
);

INVx3_ASAP7_75t_L g5767 ( 
.A(n_5372),
.Y(n_5767)
);

A2O1A1Ixp33_ASAP7_75t_L g5768 ( 
.A1(n_5500),
.A2(n_5274),
.B(n_5234),
.C(n_4954),
.Y(n_5768)
);

INVx3_ASAP7_75t_L g5769 ( 
.A(n_5381),
.Y(n_5769)
);

AO21x1_ASAP7_75t_L g5770 ( 
.A1(n_5584),
.A2(n_5068),
.B(n_5019),
.Y(n_5770)
);

NAND2xp5_ASAP7_75t_L g5771 ( 
.A(n_5529),
.B(n_5239),
.Y(n_5771)
);

AO31x2_ASAP7_75t_L g5772 ( 
.A1(n_5481),
.A2(n_5200),
.A3(n_5202),
.B(n_5135),
.Y(n_5772)
);

OAI22xp5_ASAP7_75t_L g5773 ( 
.A1(n_5558),
.A2(n_5291),
.B1(n_4874),
.B2(n_5160),
.Y(n_5773)
);

BUFx2_ASAP7_75t_L g5774 ( 
.A(n_5537),
.Y(n_5774)
);

INVx2_ASAP7_75t_L g5775 ( 
.A(n_5573),
.Y(n_5775)
);

INVx1_ASAP7_75t_L g5776 ( 
.A(n_5616),
.Y(n_5776)
);

BUFx8_ASAP7_75t_L g5777 ( 
.A(n_5455),
.Y(n_5777)
);

INVx2_ASAP7_75t_L g5778 ( 
.A(n_5575),
.Y(n_5778)
);

NAND2xp5_ASAP7_75t_L g5779 ( 
.A(n_5547),
.B(n_5276),
.Y(n_5779)
);

AOI21xp5_ASAP7_75t_L g5780 ( 
.A1(n_5607),
.A2(n_5265),
.B(n_5259),
.Y(n_5780)
);

INVx2_ASAP7_75t_L g5781 ( 
.A(n_5403),
.Y(n_5781)
);

INVx2_ASAP7_75t_L g5782 ( 
.A(n_5402),
.Y(n_5782)
);

NAND2xp5_ASAP7_75t_L g5783 ( 
.A(n_5556),
.B(n_5297),
.Y(n_5783)
);

AO21x2_ASAP7_75t_L g5784 ( 
.A1(n_5545),
.A2(n_5315),
.B(n_5300),
.Y(n_5784)
);

AND2x4_ASAP7_75t_L g5785 ( 
.A(n_5388),
.B(n_5172),
.Y(n_5785)
);

INVx1_ASAP7_75t_L g5786 ( 
.A(n_5617),
.Y(n_5786)
);

INVx2_ASAP7_75t_L g5787 ( 
.A(n_5396),
.Y(n_5787)
);

NOR2xp33_ASAP7_75t_L g5788 ( 
.A(n_5470),
.B(n_5211),
.Y(n_5788)
);

HB1xp67_ASAP7_75t_L g5789 ( 
.A(n_5587),
.Y(n_5789)
);

INVx2_ASAP7_75t_L g5790 ( 
.A(n_5629),
.Y(n_5790)
);

OAI21x1_ASAP7_75t_L g5791 ( 
.A1(n_5628),
.A2(n_5086),
.B(n_5078),
.Y(n_5791)
);

BUFx12f_ASAP7_75t_L g5792 ( 
.A(n_5508),
.Y(n_5792)
);

OR2x2_ASAP7_75t_L g5793 ( 
.A(n_5656),
.B(n_5329),
.Y(n_5793)
);

AOI21xp5_ASAP7_75t_L g5794 ( 
.A1(n_5368),
.A2(n_5126),
.B(n_5255),
.Y(n_5794)
);

NOR2xp33_ASAP7_75t_L g5795 ( 
.A(n_5539),
.B(n_5331),
.Y(n_5795)
);

INVx1_ASAP7_75t_L g5796 ( 
.A(n_5618),
.Y(n_5796)
);

CKINVDCx20_ASAP7_75t_R g5797 ( 
.A(n_5527),
.Y(n_5797)
);

INVx2_ASAP7_75t_L g5798 ( 
.A(n_5626),
.Y(n_5798)
);

OAI21x1_ASAP7_75t_L g5799 ( 
.A1(n_5484),
.A2(n_5650),
.B(n_5525),
.Y(n_5799)
);

INVx1_ASAP7_75t_SL g5800 ( 
.A(n_5498),
.Y(n_5800)
);

AOI21xp5_ASAP7_75t_L g5801 ( 
.A1(n_5430),
.A2(n_5045),
.B(n_5139),
.Y(n_5801)
);

INVx1_ASAP7_75t_L g5802 ( 
.A(n_5622),
.Y(n_5802)
);

INVx2_ASAP7_75t_L g5803 ( 
.A(n_5596),
.Y(n_5803)
);

OR2x2_ASAP7_75t_L g5804 ( 
.A(n_5624),
.B(n_5348),
.Y(n_5804)
);

NAND3xp33_ASAP7_75t_L g5805 ( 
.A(n_5493),
.B(n_5302),
.C(n_5296),
.Y(n_5805)
);

BUFx12f_ASAP7_75t_L g5806 ( 
.A(n_5593),
.Y(n_5806)
);

AO222x2_ASAP7_75t_L g5807 ( 
.A1(n_5478),
.A2(n_65),
.B1(n_67),
.B2(n_63),
.C1(n_64),
.C2(n_66),
.Y(n_5807)
);

AND2x4_ASAP7_75t_L g5808 ( 
.A(n_5642),
.B(n_5243),
.Y(n_5808)
);

NAND2xp5_ASAP7_75t_L g5809 ( 
.A(n_5557),
.B(n_5560),
.Y(n_5809)
);

OAI21x1_ASAP7_75t_L g5810 ( 
.A1(n_5411),
.A2(n_5630),
.B(n_5491),
.Y(n_5810)
);

OAI21x1_ASAP7_75t_L g5811 ( 
.A1(n_5371),
.A2(n_5140),
.B(n_5114),
.Y(n_5811)
);

INVx4_ASAP7_75t_L g5812 ( 
.A(n_5511),
.Y(n_5812)
);

OAI21x1_ASAP7_75t_L g5813 ( 
.A1(n_5375),
.A2(n_5152),
.B(n_5146),
.Y(n_5813)
);

AO31x2_ASAP7_75t_L g5814 ( 
.A1(n_5598),
.A2(n_5343),
.A3(n_5171),
.B(n_5183),
.Y(n_5814)
);

NAND2xp5_ASAP7_75t_L g5815 ( 
.A(n_5635),
.B(n_5340),
.Y(n_5815)
);

BUFx4f_ASAP7_75t_L g5816 ( 
.A(n_5551),
.Y(n_5816)
);

INVx1_ASAP7_75t_L g5817 ( 
.A(n_5373),
.Y(n_5817)
);

INVx2_ASAP7_75t_L g5818 ( 
.A(n_5439),
.Y(n_5818)
);

AOI21xp5_ASAP7_75t_L g5819 ( 
.A1(n_5472),
.A2(n_5242),
.B(n_5076),
.Y(n_5819)
);

AOI21xp5_ASAP7_75t_L g5820 ( 
.A1(n_5410),
.A2(n_5067),
.B(n_4884),
.Y(n_5820)
);

AO31x2_ASAP7_75t_L g5821 ( 
.A1(n_5636),
.A2(n_5187),
.A3(n_5221),
.B(n_5156),
.Y(n_5821)
);

INVx2_ASAP7_75t_SL g5822 ( 
.A(n_5511),
.Y(n_5822)
);

AOI21xp5_ASAP7_75t_L g5823 ( 
.A1(n_5383),
.A2(n_5050),
.B(n_5044),
.Y(n_5823)
);

INVx1_ASAP7_75t_L g5824 ( 
.A(n_5637),
.Y(n_5824)
);

AOI21xp33_ASAP7_75t_SL g5825 ( 
.A1(n_5568),
.A2(n_64),
.B(n_65),
.Y(n_5825)
);

OAI21xp5_ASAP7_75t_L g5826 ( 
.A1(n_5428),
.A2(n_4963),
.B(n_5235),
.Y(n_5826)
);

NAND2xp5_ASAP7_75t_L g5827 ( 
.A(n_5654),
.B(n_5340),
.Y(n_5827)
);

BUFx2_ASAP7_75t_L g5828 ( 
.A(n_5439),
.Y(n_5828)
);

OA21x2_ASAP7_75t_L g5829 ( 
.A1(n_5679),
.A2(n_5351),
.B(n_5489),
.Y(n_5829)
);

CKINVDCx6p67_ASAP7_75t_R g5830 ( 
.A(n_5792),
.Y(n_5830)
);

INVx2_ASAP7_75t_L g5831 ( 
.A(n_5673),
.Y(n_5831)
);

INVx1_ASAP7_75t_L g5832 ( 
.A(n_5665),
.Y(n_5832)
);

INVx1_ASAP7_75t_L g5833 ( 
.A(n_5669),
.Y(n_5833)
);

INVx1_ASAP7_75t_L g5834 ( 
.A(n_5676),
.Y(n_5834)
);

CKINVDCx20_ASAP7_75t_R g5835 ( 
.A(n_5715),
.Y(n_5835)
);

INVx2_ASAP7_75t_L g5836 ( 
.A(n_5690),
.Y(n_5836)
);

INVx1_ASAP7_75t_SL g5837 ( 
.A(n_5694),
.Y(n_5837)
);

INVx2_ASAP7_75t_SL g5838 ( 
.A(n_5763),
.Y(n_5838)
);

INVx3_ASAP7_75t_L g5839 ( 
.A(n_5744),
.Y(n_5839)
);

INVx2_ASAP7_75t_L g5840 ( 
.A(n_5690),
.Y(n_5840)
);

INVx2_ASAP7_75t_SL g5841 ( 
.A(n_5777),
.Y(n_5841)
);

INVx2_ASAP7_75t_L g5842 ( 
.A(n_5789),
.Y(n_5842)
);

AND2x2_ASAP7_75t_L g5843 ( 
.A(n_5782),
.B(n_5631),
.Y(n_5843)
);

AND2x2_ASAP7_75t_L g5844 ( 
.A(n_5781),
.B(n_5625),
.Y(n_5844)
);

INVx1_ASAP7_75t_L g5845 ( 
.A(n_5678),
.Y(n_5845)
);

INVx1_ASAP7_75t_L g5846 ( 
.A(n_5680),
.Y(n_5846)
);

NAND2xp5_ASAP7_75t_L g5847 ( 
.A(n_5817),
.B(n_5649),
.Y(n_5847)
);

NAND2x1p5_ASAP7_75t_L g5848 ( 
.A(n_5816),
.B(n_5445),
.Y(n_5848)
);

BUFx2_ASAP7_75t_L g5849 ( 
.A(n_5683),
.Y(n_5849)
);

INVx2_ASAP7_75t_L g5850 ( 
.A(n_5695),
.Y(n_5850)
);

BUFx2_ASAP7_75t_L g5851 ( 
.A(n_5683),
.Y(n_5851)
);

INVx2_ASAP7_75t_L g5852 ( 
.A(n_5696),
.Y(n_5852)
);

INVx2_ASAP7_75t_SL g5853 ( 
.A(n_5719),
.Y(n_5853)
);

AO21x2_ASAP7_75t_L g5854 ( 
.A1(n_5712),
.A2(n_5421),
.B(n_5394),
.Y(n_5854)
);

OAI21x1_ASAP7_75t_L g5855 ( 
.A1(n_5700),
.A2(n_5540),
.B(n_5389),
.Y(n_5855)
);

INVx1_ASAP7_75t_L g5856 ( 
.A(n_5681),
.Y(n_5856)
);

INVx1_ASAP7_75t_SL g5857 ( 
.A(n_5736),
.Y(n_5857)
);

INVx1_ASAP7_75t_L g5858 ( 
.A(n_5687),
.Y(n_5858)
);

INVx1_ASAP7_75t_L g5859 ( 
.A(n_5693),
.Y(n_5859)
);

INVxp33_ASAP7_75t_L g5860 ( 
.A(n_5717),
.Y(n_5860)
);

INVx2_ASAP7_75t_L g5861 ( 
.A(n_5702),
.Y(n_5861)
);

BUFx3_ASAP7_75t_L g5862 ( 
.A(n_5806),
.Y(n_5862)
);

INVx2_ASAP7_75t_L g5863 ( 
.A(n_5707),
.Y(n_5863)
);

INVx1_ASAP7_75t_L g5864 ( 
.A(n_5697),
.Y(n_5864)
);

INVx2_ASAP7_75t_L g5865 ( 
.A(n_5708),
.Y(n_5865)
);

INVx1_ASAP7_75t_L g5866 ( 
.A(n_5699),
.Y(n_5866)
);

BUFx3_ASAP7_75t_L g5867 ( 
.A(n_5797),
.Y(n_5867)
);

INVx1_ASAP7_75t_SL g5868 ( 
.A(n_5743),
.Y(n_5868)
);

INVx1_ASAP7_75t_L g5869 ( 
.A(n_5713),
.Y(n_5869)
);

INVx1_ASAP7_75t_L g5870 ( 
.A(n_5703),
.Y(n_5870)
);

INVx1_ASAP7_75t_L g5871 ( 
.A(n_5705),
.Y(n_5871)
);

OAI21xp5_ASAP7_75t_L g5872 ( 
.A1(n_5688),
.A2(n_5444),
.B(n_5536),
.Y(n_5872)
);

INVx1_ASAP7_75t_L g5873 ( 
.A(n_5776),
.Y(n_5873)
);

NOR2xp33_ASAP7_75t_L g5874 ( 
.A(n_5800),
.B(n_5614),
.Y(n_5874)
);

INVx2_ASAP7_75t_L g5875 ( 
.A(n_5714),
.Y(n_5875)
);

INVx1_ASAP7_75t_L g5876 ( 
.A(n_5786),
.Y(n_5876)
);

INVx1_ASAP7_75t_L g5877 ( 
.A(n_5796),
.Y(n_5877)
);

INVx2_ASAP7_75t_L g5878 ( 
.A(n_5722),
.Y(n_5878)
);

INVx1_ASAP7_75t_L g5879 ( 
.A(n_5802),
.Y(n_5879)
);

OA21x2_ASAP7_75t_L g5880 ( 
.A1(n_5757),
.A2(n_5733),
.B(n_5815),
.Y(n_5880)
);

INVx3_ASAP7_75t_L g5881 ( 
.A(n_5812),
.Y(n_5881)
);

AND2x4_ASAP7_75t_L g5882 ( 
.A(n_5741),
.B(n_5453),
.Y(n_5882)
);

INVx2_ASAP7_75t_L g5883 ( 
.A(n_5672),
.Y(n_5883)
);

INVx2_ASAP7_75t_L g5884 ( 
.A(n_5682),
.Y(n_5884)
);

INVx2_ASAP7_75t_L g5885 ( 
.A(n_5775),
.Y(n_5885)
);

OR2x2_ASAP7_75t_L g5886 ( 
.A(n_5727),
.B(n_5503),
.Y(n_5886)
);

INVx2_ASAP7_75t_L g5887 ( 
.A(n_5778),
.Y(n_5887)
);

INVx2_ASAP7_75t_L g5888 ( 
.A(n_5760),
.Y(n_5888)
);

INVx2_ASAP7_75t_L g5889 ( 
.A(n_5803),
.Y(n_5889)
);

NAND2xp5_ASAP7_75t_L g5890 ( 
.A(n_5731),
.B(n_5443),
.Y(n_5890)
);

AO21x2_ASAP7_75t_L g5891 ( 
.A1(n_5734),
.A2(n_5597),
.B(n_5544),
.Y(n_5891)
);

BUFx2_ASAP7_75t_L g5892 ( 
.A(n_5774),
.Y(n_5892)
);

OR2x2_ASAP7_75t_L g5893 ( 
.A(n_5662),
.B(n_5766),
.Y(n_5893)
);

INVx1_ASAP7_75t_L g5894 ( 
.A(n_5824),
.Y(n_5894)
);

NAND2xp5_ASAP7_75t_L g5895 ( 
.A(n_5759),
.B(n_5494),
.Y(n_5895)
);

INVx1_ASAP7_75t_L g5896 ( 
.A(n_5709),
.Y(n_5896)
);

INVx2_ASAP7_75t_L g5897 ( 
.A(n_5749),
.Y(n_5897)
);

INVx1_ASAP7_75t_L g5898 ( 
.A(n_5723),
.Y(n_5898)
);

INVx1_ASAP7_75t_L g5899 ( 
.A(n_5724),
.Y(n_5899)
);

INVx1_ASAP7_75t_L g5900 ( 
.A(n_5710),
.Y(n_5900)
);

AND2x2_ASAP7_75t_L g5901 ( 
.A(n_5732),
.B(n_5634),
.Y(n_5901)
);

INVx1_ASAP7_75t_L g5902 ( 
.A(n_5752),
.Y(n_5902)
);

INVx1_ASAP7_75t_L g5903 ( 
.A(n_5756),
.Y(n_5903)
);

AO21x1_ASAP7_75t_SL g5904 ( 
.A1(n_5804),
.A2(n_5609),
.B(n_5374),
.Y(n_5904)
);

INVx3_ASAP7_75t_L g5905 ( 
.A(n_5730),
.Y(n_5905)
);

INVx1_ASAP7_75t_L g5906 ( 
.A(n_5728),
.Y(n_5906)
);

AND2x2_ASAP7_75t_L g5907 ( 
.A(n_5691),
.B(n_5432),
.Y(n_5907)
);

INVx2_ASAP7_75t_SL g5908 ( 
.A(n_5674),
.Y(n_5908)
);

NAND2xp5_ASAP7_75t_L g5909 ( 
.A(n_5827),
.B(n_5615),
.Y(n_5909)
);

INVx3_ASAP7_75t_L g5910 ( 
.A(n_5758),
.Y(n_5910)
);

INVx2_ASAP7_75t_SL g5911 ( 
.A(n_5758),
.Y(n_5911)
);

INVx1_ASAP7_75t_L g5912 ( 
.A(n_5809),
.Y(n_5912)
);

AND2x2_ASAP7_75t_L g5913 ( 
.A(n_5790),
.B(n_5565),
.Y(n_5913)
);

HB1xp67_ASAP7_75t_L g5914 ( 
.A(n_5747),
.Y(n_5914)
);

INVx1_ASAP7_75t_L g5915 ( 
.A(n_5670),
.Y(n_5915)
);

INVx1_ASAP7_75t_L g5916 ( 
.A(n_5663),
.Y(n_5916)
);

INVx1_ASAP7_75t_L g5917 ( 
.A(n_5666),
.Y(n_5917)
);

NAND2xp5_ASAP7_75t_L g5918 ( 
.A(n_5798),
.B(n_5469),
.Y(n_5918)
);

INVx2_ASAP7_75t_L g5919 ( 
.A(n_5787),
.Y(n_5919)
);

AND2x2_ASAP7_75t_L g5920 ( 
.A(n_5684),
.B(n_5554),
.Y(n_5920)
);

INVx2_ASAP7_75t_L g5921 ( 
.A(n_5737),
.Y(n_5921)
);

BUFx2_ASAP7_75t_L g5922 ( 
.A(n_5741),
.Y(n_5922)
);

HB1xp67_ASAP7_75t_L g5923 ( 
.A(n_5747),
.Y(n_5923)
);

AO21x1_ASAP7_75t_SL g5924 ( 
.A1(n_5677),
.A2(n_5519),
.B(n_5442),
.Y(n_5924)
);

INVx1_ASAP7_75t_L g5925 ( 
.A(n_5685),
.Y(n_5925)
);

OR2x6_ASAP7_75t_L g5926 ( 
.A(n_5762),
.B(n_5551),
.Y(n_5926)
);

INVx2_ASAP7_75t_L g5927 ( 
.A(n_5785),
.Y(n_5927)
);

AOI21x1_ASAP7_75t_L g5928 ( 
.A1(n_5750),
.A2(n_5473),
.B(n_5467),
.Y(n_5928)
);

AOI21x1_ASAP7_75t_L g5929 ( 
.A1(n_5698),
.A2(n_5473),
.B(n_5467),
.Y(n_5929)
);

INVx2_ASAP7_75t_SL g5930 ( 
.A(n_5822),
.Y(n_5930)
);

CKINVDCx5p33_ASAP7_75t_R g5931 ( 
.A(n_5761),
.Y(n_5931)
);

AND2x2_ASAP7_75t_L g5932 ( 
.A(n_5726),
.B(n_5360),
.Y(n_5932)
);

INVx2_ASAP7_75t_L g5933 ( 
.A(n_5808),
.Y(n_5933)
);

INVx1_ASAP7_75t_L g5934 ( 
.A(n_5701),
.Y(n_5934)
);

AND2x2_ASAP7_75t_L g5935 ( 
.A(n_5793),
.B(n_5506),
.Y(n_5935)
);

OAI21x1_ASAP7_75t_L g5936 ( 
.A1(n_5668),
.A2(n_5671),
.B(n_5740),
.Y(n_5936)
);

AND2x4_ASAP7_75t_L g5937 ( 
.A(n_5818),
.B(n_5453),
.Y(n_5937)
);

AND2x4_ASAP7_75t_L g5938 ( 
.A(n_5828),
.B(n_5521),
.Y(n_5938)
);

BUFx6f_ASAP7_75t_L g5939 ( 
.A(n_5767),
.Y(n_5939)
);

INVx2_ASAP7_75t_L g5940 ( 
.A(n_5746),
.Y(n_5940)
);

BUFx6f_ASAP7_75t_L g5941 ( 
.A(n_5769),
.Y(n_5941)
);

AO31x2_ASAP7_75t_L g5942 ( 
.A1(n_5770),
.A2(n_5531),
.A3(n_5592),
.B(n_5580),
.Y(n_5942)
);

INVx2_ASAP7_75t_L g5943 ( 
.A(n_5745),
.Y(n_5943)
);

OR2x6_ASAP7_75t_L g5944 ( 
.A(n_5753),
.B(n_5640),
.Y(n_5944)
);

INVx1_ASAP7_75t_L g5945 ( 
.A(n_5729),
.Y(n_5945)
);

INVx2_ASAP7_75t_L g5946 ( 
.A(n_5755),
.Y(n_5946)
);

BUFx3_ASAP7_75t_L g5947 ( 
.A(n_5795),
.Y(n_5947)
);

AND2x2_ASAP7_75t_L g5948 ( 
.A(n_5704),
.B(n_5589),
.Y(n_5948)
);

NOR2xp33_ASAP7_75t_L g5949 ( 
.A(n_5807),
.B(n_5533),
.Y(n_5949)
);

AND2x2_ASAP7_75t_L g5950 ( 
.A(n_5771),
.B(n_5655),
.Y(n_5950)
);

INVx1_ASAP7_75t_L g5951 ( 
.A(n_5779),
.Y(n_5951)
);

AOI221xp5_ASAP7_75t_L g5952 ( 
.A1(n_5949),
.A2(n_5872),
.B1(n_5923),
.B2(n_5914),
.C(n_5773),
.Y(n_5952)
);

AOI22xp33_ASAP7_75t_L g5953 ( 
.A1(n_5904),
.A2(n_5742),
.B1(n_5686),
.B2(n_5764),
.Y(n_5953)
);

AOI22xp5_ASAP7_75t_L g5954 ( 
.A1(n_5926),
.A2(n_5735),
.B1(n_5720),
.B2(n_5706),
.Y(n_5954)
);

INVx2_ASAP7_75t_L g5955 ( 
.A(n_5892),
.Y(n_5955)
);

OA21x2_ASAP7_75t_L g5956 ( 
.A1(n_5922),
.A2(n_5783),
.B(n_5718),
.Y(n_5956)
);

OAI22xp5_ASAP7_75t_L g5957 ( 
.A1(n_5944),
.A2(n_5711),
.B1(n_5431),
.B2(n_5640),
.Y(n_5957)
);

OR2x2_ASAP7_75t_L g5958 ( 
.A(n_5934),
.B(n_5748),
.Y(n_5958)
);

INVx1_ASAP7_75t_L g5959 ( 
.A(n_5897),
.Y(n_5959)
);

OAI22xp5_ASAP7_75t_L g5960 ( 
.A1(n_5944),
.A2(n_5819),
.B1(n_5496),
.B2(n_5754),
.Y(n_5960)
);

INVx1_ASAP7_75t_L g5961 ( 
.A(n_5898),
.Y(n_5961)
);

AND2x2_ASAP7_75t_L g5962 ( 
.A(n_5892),
.B(n_5788),
.Y(n_5962)
);

AND2x4_ASAP7_75t_L g5963 ( 
.A(n_5849),
.B(n_5689),
.Y(n_5963)
);

OAI222xp33_ASAP7_75t_L g5964 ( 
.A1(n_5926),
.A2(n_5471),
.B1(n_5659),
.B2(n_5509),
.C1(n_5794),
.C2(n_5780),
.Y(n_5964)
);

AOI22xp33_ASAP7_75t_L g5965 ( 
.A1(n_5904),
.A2(n_5751),
.B1(n_5805),
.B2(n_5784),
.Y(n_5965)
);

OR2x2_ASAP7_75t_L g5966 ( 
.A(n_5893),
.B(n_5725),
.Y(n_5966)
);

OR2x2_ASAP7_75t_L g5967 ( 
.A(n_5925),
.B(n_5725),
.Y(n_5967)
);

OR2x2_ASAP7_75t_L g5968 ( 
.A(n_5917),
.B(n_5692),
.Y(n_5968)
);

AOI222xp33_ASAP7_75t_L g5969 ( 
.A1(n_5849),
.A2(n_5603),
.B1(n_5464),
.B2(n_5462),
.C1(n_5647),
.C2(n_5390),
.Y(n_5969)
);

NAND2xp5_ASAP7_75t_L g5970 ( 
.A(n_5951),
.B(n_5692),
.Y(n_5970)
);

AOI22xp33_ASAP7_75t_L g5971 ( 
.A1(n_5851),
.A2(n_5820),
.B1(n_5826),
.B2(n_5823),
.Y(n_5971)
);

AO31x2_ASAP7_75t_L g5972 ( 
.A1(n_5851),
.A2(n_5768),
.A3(n_5801),
.B(n_5479),
.Y(n_5972)
);

AOI22xp33_ASAP7_75t_L g5973 ( 
.A1(n_5829),
.A2(n_5488),
.B1(n_5664),
.B2(n_5739),
.Y(n_5973)
);

OAI22xp33_ASAP7_75t_L g5974 ( 
.A1(n_5860),
.A2(n_5825),
.B1(n_5538),
.B2(n_5532),
.Y(n_5974)
);

OAI211xp5_ASAP7_75t_L g5975 ( 
.A1(n_5874),
.A2(n_5492),
.B(n_5429),
.C(n_5651),
.Y(n_5975)
);

OAI22xp33_ASAP7_75t_L g5976 ( 
.A1(n_5839),
.A2(n_5450),
.B1(n_5648),
.B2(n_5559),
.Y(n_5976)
);

NOR2x1_ASAP7_75t_SL g5977 ( 
.A(n_5930),
.B(n_5599),
.Y(n_5977)
);

INVx1_ASAP7_75t_L g5978 ( 
.A(n_5899),
.Y(n_5978)
);

OA21x2_ASAP7_75t_L g5979 ( 
.A1(n_5922),
.A2(n_5721),
.B(n_5716),
.Y(n_5979)
);

AOI22xp33_ASAP7_75t_L g5980 ( 
.A1(n_5829),
.A2(n_5528),
.B1(n_5522),
.B2(n_5363),
.Y(n_5980)
);

AND2x2_ASAP7_75t_L g5981 ( 
.A(n_5905),
.B(n_5572),
.Y(n_5981)
);

AOI22xp33_ASAP7_75t_L g5982 ( 
.A1(n_5947),
.A2(n_5569),
.B1(n_5416),
.B2(n_5765),
.Y(n_5982)
);

BUFx6f_ASAP7_75t_L g5983 ( 
.A(n_5830),
.Y(n_5983)
);

INVx3_ASAP7_75t_L g5984 ( 
.A(n_5838),
.Y(n_5984)
);

INVx5_ASAP7_75t_SL g5985 ( 
.A(n_5938),
.Y(n_5985)
);

INVx1_ASAP7_75t_L g5986 ( 
.A(n_5902),
.Y(n_5986)
);

AOI22xp33_ASAP7_75t_L g5987 ( 
.A1(n_5854),
.A2(n_5605),
.B1(n_5542),
.B2(n_5648),
.Y(n_5987)
);

NOR2xp33_ASAP7_75t_L g5988 ( 
.A(n_5837),
.B(n_5562),
.Y(n_5988)
);

AND2x2_ASAP7_75t_L g5989 ( 
.A(n_5933),
.B(n_5814),
.Y(n_5989)
);

AND2x2_ASAP7_75t_L g5990 ( 
.A(n_5927),
.B(n_5814),
.Y(n_5990)
);

AOI22xp33_ASAP7_75t_L g5991 ( 
.A1(n_5924),
.A2(n_5542),
.B1(n_5566),
.B2(n_5610),
.Y(n_5991)
);

CKINVDCx20_ASAP7_75t_R g5992 ( 
.A(n_5835),
.Y(n_5992)
);

INVx2_ASAP7_75t_SL g5993 ( 
.A(n_5841),
.Y(n_5993)
);

A2O1A1Ixp33_ASAP7_75t_L g5994 ( 
.A1(n_5853),
.A2(n_5581),
.B(n_5449),
.C(n_5639),
.Y(n_5994)
);

AOI22xp33_ASAP7_75t_L g5995 ( 
.A1(n_5924),
.A2(n_5610),
.B1(n_5574),
.B2(n_5638),
.Y(n_5995)
);

AOI221xp5_ASAP7_75t_L g5996 ( 
.A1(n_5946),
.A2(n_5398),
.B1(n_5543),
.B2(n_5458),
.C(n_5611),
.Y(n_5996)
);

OR2x2_ASAP7_75t_L g5997 ( 
.A(n_5915),
.B(n_5420),
.Y(n_5997)
);

AOI22xp33_ASAP7_75t_SL g5998 ( 
.A1(n_5901),
.A2(n_5550),
.B1(n_5517),
.B2(n_5644),
.Y(n_5998)
);

NAND2xp5_ASAP7_75t_L g5999 ( 
.A(n_5912),
.B(n_5772),
.Y(n_5999)
);

HB1xp67_ASAP7_75t_L g6000 ( 
.A(n_5889),
.Y(n_6000)
);

AOI221xp5_ASAP7_75t_L g6001 ( 
.A1(n_5909),
.A2(n_5945),
.B1(n_5940),
.B2(n_5916),
.C(n_5943),
.Y(n_6001)
);

OR2x2_ASAP7_75t_L g6002 ( 
.A(n_5919),
.B(n_5886),
.Y(n_6002)
);

AOI22xp5_ASAP7_75t_L g6003 ( 
.A1(n_5891),
.A2(n_5482),
.B1(n_5518),
.B2(n_5365),
.Y(n_6003)
);

INVx1_ASAP7_75t_L g6004 ( 
.A(n_5903),
.Y(n_6004)
);

OAI22xp5_ASAP7_75t_L g6005 ( 
.A1(n_5857),
.A2(n_5564),
.B1(n_5570),
.B2(n_5632),
.Y(n_6005)
);

NAND3xp33_ASAP7_75t_L g6006 ( 
.A(n_5880),
.B(n_5921),
.C(n_5840),
.Y(n_6006)
);

INVx1_ASAP7_75t_L g6007 ( 
.A(n_5832),
.Y(n_6007)
);

NAND2xp5_ASAP7_75t_L g6008 ( 
.A(n_5900),
.B(n_5772),
.Y(n_6008)
);

NAND2xp5_ASAP7_75t_L g6009 ( 
.A(n_5873),
.B(n_5497),
.Y(n_6009)
);

AOI22xp33_ASAP7_75t_L g6010 ( 
.A1(n_5842),
.A2(n_5811),
.B1(n_5813),
.B2(n_5604),
.Y(n_6010)
);

AOI221xp5_ASAP7_75t_L g6011 ( 
.A1(n_5918),
.A2(n_5461),
.B1(n_5653),
.B2(n_5612),
.C(n_5633),
.Y(n_6011)
);

INVx2_ASAP7_75t_L g6012 ( 
.A(n_5850),
.Y(n_6012)
);

NOR2x1_ASAP7_75t_L g6013 ( 
.A(n_5868),
.B(n_5517),
.Y(n_6013)
);

INVx1_ASAP7_75t_L g6014 ( 
.A(n_5833),
.Y(n_6014)
);

AOI22xp33_ASAP7_75t_SL g6015 ( 
.A1(n_5881),
.A2(n_5738),
.B1(n_5667),
.B2(n_5530),
.Y(n_6015)
);

AOI221xp5_ASAP7_75t_L g6016 ( 
.A1(n_5847),
.A2(n_5261),
.B1(n_5661),
.B2(n_5594),
.C(n_5600),
.Y(n_6016)
);

OAI221xp5_ASAP7_75t_L g6017 ( 
.A1(n_5848),
.A2(n_5293),
.B1(n_5308),
.B2(n_5290),
.C(n_5238),
.Y(n_6017)
);

AOI22xp33_ASAP7_75t_L g6018 ( 
.A1(n_5920),
.A2(n_5530),
.B1(n_5791),
.B2(n_5546),
.Y(n_6018)
);

AOI22xp33_ASAP7_75t_L g6019 ( 
.A1(n_5935),
.A2(n_5546),
.B1(n_5646),
.B2(n_5799),
.Y(n_6019)
);

AOI21xp5_ASAP7_75t_L g6020 ( 
.A1(n_5855),
.A2(n_5810),
.B(n_5675),
.Y(n_6020)
);

OAI33xp33_ASAP7_75t_L g6021 ( 
.A1(n_5890),
.A2(n_4984),
.A3(n_5608),
.B1(n_5192),
.B2(n_5203),
.B3(n_5321),
.Y(n_6021)
);

INVx2_ASAP7_75t_L g6022 ( 
.A(n_5852),
.Y(n_6022)
);

AND2x2_ASAP7_75t_L g6023 ( 
.A(n_5843),
.B(n_5821),
.Y(n_6023)
);

NAND2xp5_ASAP7_75t_L g6024 ( 
.A(n_5876),
.B(n_5379),
.Y(n_6024)
);

AOI221xp5_ASAP7_75t_L g6025 ( 
.A1(n_5877),
.A2(n_5326),
.B1(n_5337),
.B2(n_5334),
.C(n_5311),
.Y(n_6025)
);

NAND2xp5_ASAP7_75t_L g6026 ( 
.A(n_5879),
.B(n_5379),
.Y(n_6026)
);

OAI21x1_ASAP7_75t_L g6027 ( 
.A1(n_5936),
.A2(n_5436),
.B(n_5553),
.Y(n_6027)
);

OAI22xp33_ASAP7_75t_L g6028 ( 
.A1(n_5908),
.A2(n_4984),
.B1(n_5608),
.B2(n_5189),
.Y(n_6028)
);

AOI22xp5_ASAP7_75t_L g6029 ( 
.A1(n_5913),
.A2(n_5504),
.B1(n_5377),
.B2(n_5591),
.Y(n_6029)
);

INVx3_ASAP7_75t_SL g6030 ( 
.A(n_5931),
.Y(n_6030)
);

OR2x2_ASAP7_75t_L g6031 ( 
.A(n_5831),
.B(n_5451),
.Y(n_6031)
);

AOI222xp33_ASAP7_75t_L g6032 ( 
.A1(n_5895),
.A2(n_5485),
.B1(n_5619),
.B2(n_5620),
.C1(n_5595),
.C2(n_5657),
.Y(n_6032)
);

OR2x2_ASAP7_75t_L g6033 ( 
.A(n_5883),
.B(n_5451),
.Y(n_6033)
);

AOI22xp33_ASAP7_75t_L g6034 ( 
.A1(n_5932),
.A2(n_5590),
.B1(n_5641),
.B2(n_5643),
.Y(n_6034)
);

OAI221xp5_ASAP7_75t_L g6035 ( 
.A1(n_5867),
.A2(n_5192),
.B1(n_5203),
.B2(n_5321),
.C(n_5189),
.Y(n_6035)
);

OAI22xp5_ASAP7_75t_L g6036 ( 
.A1(n_5939),
.A2(n_5203),
.B1(n_5535),
.B2(n_5821),
.Y(n_6036)
);

OAI22xp5_ASAP7_75t_L g6037 ( 
.A1(n_5939),
.A2(n_5535),
.B1(n_5220),
.B2(n_5213),
.Y(n_6037)
);

OAI211xp5_ASAP7_75t_L g6038 ( 
.A1(n_5907),
.A2(n_5579),
.B(n_5660),
.C(n_5652),
.Y(n_6038)
);

OR2x2_ASAP7_75t_L g6039 ( 
.A(n_5884),
.B(n_5220),
.Y(n_6039)
);

INVx2_ASAP7_75t_L g6040 ( 
.A(n_5861),
.Y(n_6040)
);

NAND3xp33_ASAP7_75t_L g6041 ( 
.A(n_5880),
.B(n_5548),
.C(n_5658),
.Y(n_6041)
);

OAI221xp5_ASAP7_75t_L g6042 ( 
.A1(n_5906),
.A2(n_5213),
.B1(n_66),
.B2(n_64),
.C(n_65),
.Y(n_6042)
);

AOI221xp5_ASAP7_75t_L g6043 ( 
.A1(n_5894),
.A2(n_1052),
.B1(n_1053),
.B2(n_1051),
.C(n_1050),
.Y(n_6043)
);

INVxp67_ASAP7_75t_L g6044 ( 
.A(n_5948),
.Y(n_6044)
);

INVx1_ASAP7_75t_L g6045 ( 
.A(n_5834),
.Y(n_6045)
);

AOI22xp33_ASAP7_75t_L g6046 ( 
.A1(n_5844),
.A2(n_5571),
.B1(n_5576),
.B2(n_5552),
.Y(n_6046)
);

OAI22xp5_ASAP7_75t_L g6047 ( 
.A1(n_5941),
.A2(n_5459),
.B1(n_5460),
.B2(n_5513),
.Y(n_6047)
);

BUFx10_ASAP7_75t_L g6048 ( 
.A(n_5862),
.Y(n_6048)
);

AOI211xp5_ASAP7_75t_L g6049 ( 
.A1(n_5882),
.A2(n_5623),
.B(n_5621),
.C(n_5567),
.Y(n_6049)
);

OAI222xp33_ASAP7_75t_L g6050 ( 
.A1(n_5882),
.A2(n_5627),
.B1(n_5495),
.B2(n_5435),
.C1(n_5477),
.C2(n_1056),
.Y(n_6050)
);

NAND2xp5_ASAP7_75t_L g6051 ( 
.A(n_5970),
.B(n_5942),
.Y(n_6051)
);

INVx3_ASAP7_75t_L g6052 ( 
.A(n_5985),
.Y(n_6052)
);

AND2x2_ASAP7_75t_L g6053 ( 
.A(n_6023),
.B(n_5941),
.Y(n_6053)
);

AND2x2_ASAP7_75t_L g6054 ( 
.A(n_5962),
.B(n_5938),
.Y(n_6054)
);

XNOR2xp5_ASAP7_75t_L g6055 ( 
.A(n_5992),
.B(n_5957),
.Y(n_6055)
);

INVxp67_ASAP7_75t_L g6056 ( 
.A(n_5983),
.Y(n_6056)
);

AND2x2_ASAP7_75t_L g6057 ( 
.A(n_5981),
.B(n_5911),
.Y(n_6057)
);

INVx2_ASAP7_75t_L g6058 ( 
.A(n_6000),
.Y(n_6058)
);

INVx1_ASAP7_75t_L g6059 ( 
.A(n_6031),
.Y(n_6059)
);

BUFx3_ASAP7_75t_L g6060 ( 
.A(n_6048),
.Y(n_6060)
);

INVx1_ASAP7_75t_L g6061 ( 
.A(n_5968),
.Y(n_6061)
);

OR2x2_ASAP7_75t_L g6062 ( 
.A(n_6002),
.B(n_5885),
.Y(n_6062)
);

AOI22xp33_ASAP7_75t_L g6063 ( 
.A1(n_5952),
.A2(n_5950),
.B1(n_5910),
.B2(n_5937),
.Y(n_6063)
);

OR2x2_ASAP7_75t_L g6064 ( 
.A(n_5958),
.B(n_5887),
.Y(n_6064)
);

NOR3xp33_ASAP7_75t_L g6065 ( 
.A(n_5960),
.B(n_5929),
.C(n_5928),
.Y(n_6065)
);

NAND2xp5_ASAP7_75t_L g6066 ( 
.A(n_6001),
.B(n_5973),
.Y(n_6066)
);

NAND2xp5_ASAP7_75t_L g6067 ( 
.A(n_5999),
.B(n_5942),
.Y(n_6067)
);

INVx1_ASAP7_75t_L g6068 ( 
.A(n_5961),
.Y(n_6068)
);

OR2x2_ASAP7_75t_L g6069 ( 
.A(n_5966),
.B(n_6039),
.Y(n_6069)
);

INVx2_ASAP7_75t_L g6070 ( 
.A(n_6012),
.Y(n_6070)
);

NAND2xp5_ASAP7_75t_L g6071 ( 
.A(n_5967),
.B(n_5942),
.Y(n_6071)
);

NAND2xp5_ASAP7_75t_L g6072 ( 
.A(n_5971),
.B(n_5845),
.Y(n_6072)
);

INVx1_ASAP7_75t_L g6073 ( 
.A(n_5978),
.Y(n_6073)
);

AND2x2_ASAP7_75t_L g6074 ( 
.A(n_5963),
.B(n_5937),
.Y(n_6074)
);

OR2x2_ASAP7_75t_L g6075 ( 
.A(n_5955),
.B(n_5863),
.Y(n_6075)
);

AND2x4_ASAP7_75t_L g6076 ( 
.A(n_5990),
.B(n_5846),
.Y(n_6076)
);

OR2x2_ASAP7_75t_L g6077 ( 
.A(n_6009),
.B(n_6024),
.Y(n_6077)
);

NAND2xp5_ASAP7_75t_L g6078 ( 
.A(n_6026),
.B(n_5856),
.Y(n_6078)
);

INVx1_ASAP7_75t_L g6079 ( 
.A(n_5986),
.Y(n_6079)
);

INVx1_ASAP7_75t_L g6080 ( 
.A(n_6004),
.Y(n_6080)
);

AOI22xp33_ASAP7_75t_L g6081 ( 
.A1(n_5953),
.A2(n_5896),
.B1(n_5859),
.B2(n_5864),
.Y(n_6081)
);

AND2x2_ASAP7_75t_L g6082 ( 
.A(n_5989),
.B(n_5858),
.Y(n_6082)
);

INVx2_ASAP7_75t_L g6083 ( 
.A(n_6022),
.Y(n_6083)
);

INVx1_ASAP7_75t_L g6084 ( 
.A(n_6007),
.Y(n_6084)
);

AOI22xp33_ASAP7_75t_SL g6085 ( 
.A1(n_5977),
.A2(n_5869),
.B1(n_5870),
.B2(n_5866),
.Y(n_6085)
);

INVx1_ASAP7_75t_SL g6086 ( 
.A(n_5984),
.Y(n_6086)
);

AOI22xp33_ASAP7_75t_L g6087 ( 
.A1(n_5965),
.A2(n_5871),
.B1(n_5836),
.B2(n_5888),
.Y(n_6087)
);

INVx1_ASAP7_75t_L g6088 ( 
.A(n_6033),
.Y(n_6088)
);

INVx1_ASAP7_75t_L g6089 ( 
.A(n_6014),
.Y(n_6089)
);

AND2x2_ASAP7_75t_L g6090 ( 
.A(n_5985),
.B(n_5865),
.Y(n_6090)
);

INVx1_ASAP7_75t_L g6091 ( 
.A(n_6045),
.Y(n_6091)
);

OR2x2_ASAP7_75t_L g6092 ( 
.A(n_5997),
.B(n_5875),
.Y(n_6092)
);

OR2x2_ASAP7_75t_L g6093 ( 
.A(n_6008),
.B(n_5878),
.Y(n_6093)
);

AND2x2_ASAP7_75t_L g6094 ( 
.A(n_6044),
.B(n_5928),
.Y(n_6094)
);

INVx1_ASAP7_75t_L g6095 ( 
.A(n_5959),
.Y(n_6095)
);

AND2x2_ASAP7_75t_L g6096 ( 
.A(n_5954),
.B(n_5929),
.Y(n_6096)
);

AND2x4_ASAP7_75t_L g6097 ( 
.A(n_6006),
.B(n_5602),
.Y(n_6097)
);

OAI222xp33_ASAP7_75t_L g6098 ( 
.A1(n_6035),
.A2(n_67),
.B1(n_69),
.B2(n_65),
.C1(n_66),
.C2(n_68),
.Y(n_6098)
);

AND2x2_ASAP7_75t_L g6099 ( 
.A(n_5956),
.B(n_66),
.Y(n_6099)
);

INVx1_ASAP7_75t_L g6100 ( 
.A(n_6040),
.Y(n_6100)
);

AND2x2_ASAP7_75t_L g6101 ( 
.A(n_5956),
.B(n_67),
.Y(n_6101)
);

INVx2_ASAP7_75t_L g6102 ( 
.A(n_5979),
.Y(n_6102)
);

INVx1_ASAP7_75t_L g6103 ( 
.A(n_6041),
.Y(n_6103)
);

BUFx2_ASAP7_75t_L g6104 ( 
.A(n_5993),
.Y(n_6104)
);

AOI22xp33_ASAP7_75t_L g6105 ( 
.A1(n_5969),
.A2(n_1148),
.B1(n_1054),
.B2(n_1055),
.Y(n_6105)
);

AND2x2_ASAP7_75t_L g6106 ( 
.A(n_5979),
.B(n_5988),
.Y(n_6106)
);

INVx2_ASAP7_75t_L g6107 ( 
.A(n_6013),
.Y(n_6107)
);

NAND2xp5_ASAP7_75t_L g6108 ( 
.A(n_5972),
.B(n_6028),
.Y(n_6108)
);

INVx2_ASAP7_75t_L g6109 ( 
.A(n_6027),
.Y(n_6109)
);

NAND2xp5_ASAP7_75t_L g6110 ( 
.A(n_5972),
.B(n_1052),
.Y(n_6110)
);

OR2x2_ASAP7_75t_L g6111 ( 
.A(n_6036),
.B(n_67),
.Y(n_6111)
);

AND2x2_ASAP7_75t_L g6112 ( 
.A(n_6020),
.B(n_68),
.Y(n_6112)
);

INVx2_ASAP7_75t_L g6113 ( 
.A(n_6029),
.Y(n_6113)
);

CKINVDCx14_ASAP7_75t_R g6114 ( 
.A(n_5983),
.Y(n_6114)
);

AND2x2_ASAP7_75t_L g6115 ( 
.A(n_6010),
.B(n_68),
.Y(n_6115)
);

NAND2xp5_ASAP7_75t_L g6116 ( 
.A(n_6003),
.B(n_1054),
.Y(n_6116)
);

INVxp67_ASAP7_75t_L g6117 ( 
.A(n_5994),
.Y(n_6117)
);

AND2x2_ASAP7_75t_L g6118 ( 
.A(n_6030),
.B(n_69),
.Y(n_6118)
);

INVx1_ASAP7_75t_L g6119 ( 
.A(n_6037),
.Y(n_6119)
);

INVx1_ASAP7_75t_L g6120 ( 
.A(n_6049),
.Y(n_6120)
);

INVx4_ASAP7_75t_L g6121 ( 
.A(n_5964),
.Y(n_6121)
);

INVx2_ASAP7_75t_L g6122 ( 
.A(n_6047),
.Y(n_6122)
);

NAND2xp5_ASAP7_75t_L g6123 ( 
.A(n_5982),
.B(n_1054),
.Y(n_6123)
);

NAND2xp5_ASAP7_75t_L g6124 ( 
.A(n_5987),
.B(n_1055),
.Y(n_6124)
);

NAND2xp5_ASAP7_75t_L g6125 ( 
.A(n_6120),
.B(n_5980),
.Y(n_6125)
);

INVx1_ASAP7_75t_L g6126 ( 
.A(n_6095),
.Y(n_6126)
);

NAND2xp5_ASAP7_75t_L g6127 ( 
.A(n_6120),
.B(n_5991),
.Y(n_6127)
);

NAND4xp25_ASAP7_75t_L g6128 ( 
.A(n_6121),
.B(n_5996),
.C(n_5975),
.D(n_5995),
.Y(n_6128)
);

AND2x2_ASAP7_75t_L g6129 ( 
.A(n_6074),
.B(n_6015),
.Y(n_6129)
);

NAND3xp33_ASAP7_75t_L g6130 ( 
.A(n_6065),
.B(n_5998),
.C(n_6038),
.Y(n_6130)
);

HB1xp67_ASAP7_75t_L g6131 ( 
.A(n_6058),
.Y(n_6131)
);

INVx1_ASAP7_75t_L g6132 ( 
.A(n_6092),
.Y(n_6132)
);

AND2x2_ASAP7_75t_L g6133 ( 
.A(n_6104),
.B(n_6053),
.Y(n_6133)
);

AND2x2_ASAP7_75t_L g6134 ( 
.A(n_6052),
.B(n_6019),
.Y(n_6134)
);

INVx1_ASAP7_75t_SL g6135 ( 
.A(n_6060),
.Y(n_6135)
);

OR2x6_ASAP7_75t_SL g6136 ( 
.A(n_6108),
.B(n_6005),
.Y(n_6136)
);

INVx2_ASAP7_75t_L g6137 ( 
.A(n_6062),
.Y(n_6137)
);

INVx2_ASAP7_75t_L g6138 ( 
.A(n_6064),
.Y(n_6138)
);

HB1xp67_ASAP7_75t_L g6139 ( 
.A(n_6061),
.Y(n_6139)
);

AND2x4_ASAP7_75t_SL g6140 ( 
.A(n_6052),
.B(n_6046),
.Y(n_6140)
);

INVx4_ASAP7_75t_L g6141 ( 
.A(n_6114),
.Y(n_6141)
);

AND2x2_ASAP7_75t_L g6142 ( 
.A(n_6106),
.B(n_6018),
.Y(n_6142)
);

NAND2xp5_ASAP7_75t_L g6143 ( 
.A(n_6099),
.B(n_6032),
.Y(n_6143)
);

NAND2xp5_ASAP7_75t_L g6144 ( 
.A(n_6101),
.B(n_5976),
.Y(n_6144)
);

AND2x2_ASAP7_75t_L g6145 ( 
.A(n_6086),
.B(n_6034),
.Y(n_6145)
);

NOR2xp33_ASAP7_75t_L g6146 ( 
.A(n_6056),
.B(n_5974),
.Y(n_6146)
);

AND2x2_ASAP7_75t_L g6147 ( 
.A(n_6094),
.B(n_6025),
.Y(n_6147)
);

AND2x2_ASAP7_75t_L g6148 ( 
.A(n_6082),
.B(n_6011),
.Y(n_6148)
);

AND2x4_ASAP7_75t_L g6149 ( 
.A(n_6122),
.B(n_1055),
.Y(n_6149)
);

NOR2xp33_ASAP7_75t_L g6150 ( 
.A(n_6055),
.B(n_6021),
.Y(n_6150)
);

AND2x2_ASAP7_75t_L g6151 ( 
.A(n_6121),
.B(n_6016),
.Y(n_6151)
);

AND2x2_ASAP7_75t_L g6152 ( 
.A(n_6076),
.B(n_6043),
.Y(n_6152)
);

NAND2xp5_ASAP7_75t_L g6153 ( 
.A(n_6112),
.B(n_6042),
.Y(n_6153)
);

INVx1_ASAP7_75t_L g6154 ( 
.A(n_6078),
.Y(n_6154)
);

AND2x2_ASAP7_75t_L g6155 ( 
.A(n_6076),
.B(n_69),
.Y(n_6155)
);

NOR2xp33_ASAP7_75t_L g6156 ( 
.A(n_6117),
.B(n_6050),
.Y(n_6156)
);

NAND2xp5_ASAP7_75t_SL g6157 ( 
.A(n_6085),
.B(n_6017),
.Y(n_6157)
);

AOI21xp33_ASAP7_75t_L g6158 ( 
.A1(n_6066),
.A2(n_70),
.B(n_71),
.Y(n_6158)
);

INVx1_ASAP7_75t_L g6159 ( 
.A(n_6068),
.Y(n_6159)
);

INVx1_ASAP7_75t_L g6160 ( 
.A(n_6073),
.Y(n_6160)
);

NAND2xp5_ASAP7_75t_L g6161 ( 
.A(n_6051),
.B(n_70),
.Y(n_6161)
);

INVx1_ASAP7_75t_L g6162 ( 
.A(n_6079),
.Y(n_6162)
);

NOR2xp67_ASAP7_75t_L g6163 ( 
.A(n_6107),
.B(n_70),
.Y(n_6163)
);

OAI221xp5_ASAP7_75t_SL g6164 ( 
.A1(n_6063),
.A2(n_1058),
.B1(n_1059),
.B2(n_1057),
.C(n_1056),
.Y(n_6164)
);

AND2x2_ASAP7_75t_L g6165 ( 
.A(n_6054),
.B(n_70),
.Y(n_6165)
);

AND2x2_ASAP7_75t_L g6166 ( 
.A(n_6090),
.B(n_71),
.Y(n_6166)
);

BUFx2_ASAP7_75t_L g6167 ( 
.A(n_6057),
.Y(n_6167)
);

AND2x2_ASAP7_75t_L g6168 ( 
.A(n_6119),
.B(n_72),
.Y(n_6168)
);

INVx1_ASAP7_75t_L g6169 ( 
.A(n_6080),
.Y(n_6169)
);

NAND2xp5_ASAP7_75t_L g6170 ( 
.A(n_6067),
.B(n_72),
.Y(n_6170)
);

NAND2xp5_ASAP7_75t_L g6171 ( 
.A(n_6113),
.B(n_73),
.Y(n_6171)
);

NOR2xp33_ASAP7_75t_L g6172 ( 
.A(n_6072),
.B(n_6098),
.Y(n_6172)
);

INVx1_ASAP7_75t_L g6173 ( 
.A(n_6084),
.Y(n_6173)
);

AND2x2_ASAP7_75t_L g6174 ( 
.A(n_6119),
.B(n_73),
.Y(n_6174)
);

NAND2xp5_ASAP7_75t_L g6175 ( 
.A(n_6071),
.B(n_73),
.Y(n_6175)
);

CKINVDCx20_ASAP7_75t_R g6176 ( 
.A(n_6118),
.Y(n_6176)
);

INVx1_ASAP7_75t_L g6177 ( 
.A(n_6089),
.Y(n_6177)
);

OR2x2_ASAP7_75t_L g6178 ( 
.A(n_6077),
.B(n_73),
.Y(n_6178)
);

INVx2_ASAP7_75t_SL g6179 ( 
.A(n_6075),
.Y(n_6179)
);

NAND2xp5_ASAP7_75t_L g6180 ( 
.A(n_6096),
.B(n_74),
.Y(n_6180)
);

AND2x2_ASAP7_75t_L g6181 ( 
.A(n_6059),
.B(n_74),
.Y(n_6181)
);

INVx1_ASAP7_75t_L g6182 ( 
.A(n_6091),
.Y(n_6182)
);

NAND2xp5_ASAP7_75t_L g6183 ( 
.A(n_6110),
.B(n_74),
.Y(n_6183)
);

AND2x4_ASAP7_75t_L g6184 ( 
.A(n_6109),
.B(n_1056),
.Y(n_6184)
);

INVx2_ASAP7_75t_L g6185 ( 
.A(n_6070),
.Y(n_6185)
);

NAND2xp5_ASAP7_75t_L g6186 ( 
.A(n_6081),
.B(n_75),
.Y(n_6186)
);

AND2x4_ASAP7_75t_L g6187 ( 
.A(n_6088),
.B(n_1057),
.Y(n_6187)
);

NAND2xp5_ASAP7_75t_L g6188 ( 
.A(n_6103),
.B(n_75),
.Y(n_6188)
);

INVxp67_ASAP7_75t_SL g6189 ( 
.A(n_6111),
.Y(n_6189)
);

INVx2_ASAP7_75t_L g6190 ( 
.A(n_6083),
.Y(n_6190)
);

INVx2_ASAP7_75t_SL g6191 ( 
.A(n_6093),
.Y(n_6191)
);

AND2x2_ASAP7_75t_L g6192 ( 
.A(n_6088),
.B(n_75),
.Y(n_6192)
);

AND2x2_ASAP7_75t_L g6193 ( 
.A(n_6133),
.B(n_6087),
.Y(n_6193)
);

AND2x2_ASAP7_75t_L g6194 ( 
.A(n_6167),
.B(n_6069),
.Y(n_6194)
);

AOI22xp33_ASAP7_75t_L g6195 ( 
.A1(n_6128),
.A2(n_6105),
.B1(n_6097),
.B2(n_6115),
.Y(n_6195)
);

AND2x2_ASAP7_75t_L g6196 ( 
.A(n_6134),
.B(n_6102),
.Y(n_6196)
);

INVx1_ASAP7_75t_L g6197 ( 
.A(n_6139),
.Y(n_6197)
);

INVx1_ASAP7_75t_L g6198 ( 
.A(n_6126),
.Y(n_6198)
);

INVx1_ASAP7_75t_L g6199 ( 
.A(n_6187),
.Y(n_6199)
);

INVx1_ASAP7_75t_L g6200 ( 
.A(n_6187),
.Y(n_6200)
);

INVx1_ASAP7_75t_L g6201 ( 
.A(n_6192),
.Y(n_6201)
);

AND2x2_ASAP7_75t_L g6202 ( 
.A(n_6146),
.B(n_6168),
.Y(n_6202)
);

AND2x2_ASAP7_75t_L g6203 ( 
.A(n_6174),
.B(n_6097),
.Y(n_6203)
);

BUFx3_ASAP7_75t_L g6204 ( 
.A(n_6141),
.Y(n_6204)
);

INVx1_ASAP7_75t_L g6205 ( 
.A(n_6132),
.Y(n_6205)
);

AND2x4_ASAP7_75t_L g6206 ( 
.A(n_6135),
.B(n_6124),
.Y(n_6206)
);

OAI211xp5_ASAP7_75t_SL g6207 ( 
.A1(n_6125),
.A2(n_6116),
.B(n_6123),
.C(n_6100),
.Y(n_6207)
);

AND2x2_ASAP7_75t_SL g6208 ( 
.A(n_6141),
.B(n_1057),
.Y(n_6208)
);

INVxp67_ASAP7_75t_SL g6209 ( 
.A(n_6163),
.Y(n_6209)
);

BUFx3_ASAP7_75t_L g6210 ( 
.A(n_6166),
.Y(n_6210)
);

HB1xp67_ASAP7_75t_L g6211 ( 
.A(n_6131),
.Y(n_6211)
);

INVx1_ASAP7_75t_L g6212 ( 
.A(n_6126),
.Y(n_6212)
);

AND2x2_ASAP7_75t_L g6213 ( 
.A(n_6129),
.B(n_75),
.Y(n_6213)
);

AOI221xp5_ASAP7_75t_L g6214 ( 
.A1(n_6151),
.A2(n_1061),
.B1(n_1062),
.B2(n_1060),
.C(n_1059),
.Y(n_6214)
);

INVx1_ASAP7_75t_L g6215 ( 
.A(n_6159),
.Y(n_6215)
);

AND2x2_ASAP7_75t_L g6216 ( 
.A(n_6140),
.B(n_76),
.Y(n_6216)
);

INVx3_ASAP7_75t_L g6217 ( 
.A(n_6184),
.Y(n_6217)
);

INVx2_ASAP7_75t_L g6218 ( 
.A(n_6137),
.Y(n_6218)
);

AND2x2_ASAP7_75t_L g6219 ( 
.A(n_6145),
.B(n_76),
.Y(n_6219)
);

AND2x2_ASAP7_75t_L g6220 ( 
.A(n_6189),
.B(n_6149),
.Y(n_6220)
);

AOI22xp5_ASAP7_75t_L g6221 ( 
.A1(n_6150),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_6221)
);

INVx2_ASAP7_75t_L g6222 ( 
.A(n_6179),
.Y(n_6222)
);

BUFx2_ASAP7_75t_L g6223 ( 
.A(n_6184),
.Y(n_6223)
);

INVx2_ASAP7_75t_L g6224 ( 
.A(n_6138),
.Y(n_6224)
);

HB1xp67_ASAP7_75t_L g6225 ( 
.A(n_6180),
.Y(n_6225)
);

INVx1_ASAP7_75t_L g6226 ( 
.A(n_6181),
.Y(n_6226)
);

AND2x4_ASAP7_75t_L g6227 ( 
.A(n_6149),
.B(n_1059),
.Y(n_6227)
);

NAND2xp5_ASAP7_75t_L g6228 ( 
.A(n_6148),
.B(n_76),
.Y(n_6228)
);

INVx1_ASAP7_75t_L g6229 ( 
.A(n_6159),
.Y(n_6229)
);

INVx1_ASAP7_75t_L g6230 ( 
.A(n_6160),
.Y(n_6230)
);

AND2x2_ASAP7_75t_L g6231 ( 
.A(n_6152),
.B(n_6147),
.Y(n_6231)
);

AND2x4_ASAP7_75t_SL g6232 ( 
.A(n_6165),
.B(n_77),
.Y(n_6232)
);

AOI22xp5_ASAP7_75t_L g6233 ( 
.A1(n_6156),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_6233)
);

INVx2_ASAP7_75t_L g6234 ( 
.A(n_6191),
.Y(n_6234)
);

INVx1_ASAP7_75t_L g6235 ( 
.A(n_6162),
.Y(n_6235)
);

NAND2xp5_ASAP7_75t_L g6236 ( 
.A(n_6172),
.B(n_78),
.Y(n_6236)
);

AND2x2_ASAP7_75t_L g6237 ( 
.A(n_6204),
.B(n_6142),
.Y(n_6237)
);

AND2x2_ASAP7_75t_L g6238 ( 
.A(n_6220),
.B(n_6154),
.Y(n_6238)
);

AND2x2_ASAP7_75t_L g6239 ( 
.A(n_6196),
.B(n_6157),
.Y(n_6239)
);

AND2x2_ASAP7_75t_L g6240 ( 
.A(n_6206),
.B(n_6136),
.Y(n_6240)
);

INVx1_ASAP7_75t_SL g6241 ( 
.A(n_6216),
.Y(n_6241)
);

AND2x2_ASAP7_75t_L g6242 ( 
.A(n_6206),
.B(n_6209),
.Y(n_6242)
);

INVx1_ASAP7_75t_L g6243 ( 
.A(n_6211),
.Y(n_6243)
);

AND2x4_ASAP7_75t_L g6244 ( 
.A(n_6234),
.B(n_6176),
.Y(n_6244)
);

AND2x2_ASAP7_75t_L g6245 ( 
.A(n_6203),
.B(n_6194),
.Y(n_6245)
);

INVx2_ASAP7_75t_L g6246 ( 
.A(n_6222),
.Y(n_6246)
);

AND2x2_ASAP7_75t_L g6247 ( 
.A(n_6223),
.B(n_6144),
.Y(n_6247)
);

NAND2x1_ASAP7_75t_L g6248 ( 
.A(n_6217),
.B(n_6130),
.Y(n_6248)
);

NAND2xp5_ASAP7_75t_L g6249 ( 
.A(n_6231),
.B(n_6127),
.Y(n_6249)
);

INVx1_ASAP7_75t_L g6250 ( 
.A(n_6197),
.Y(n_6250)
);

AND2x2_ASAP7_75t_L g6251 ( 
.A(n_6202),
.B(n_6171),
.Y(n_6251)
);

INVx1_ASAP7_75t_L g6252 ( 
.A(n_6197),
.Y(n_6252)
);

AND2x2_ASAP7_75t_L g6253 ( 
.A(n_6219),
.B(n_6155),
.Y(n_6253)
);

BUFx2_ASAP7_75t_L g6254 ( 
.A(n_6217),
.Y(n_6254)
);

AND2x2_ASAP7_75t_L g6255 ( 
.A(n_6210),
.B(n_6143),
.Y(n_6255)
);

INVx2_ASAP7_75t_L g6256 ( 
.A(n_6218),
.Y(n_6256)
);

AND2x2_ASAP7_75t_L g6257 ( 
.A(n_6193),
.B(n_6188),
.Y(n_6257)
);

NOR2x1_ASAP7_75t_L g6258 ( 
.A(n_6236),
.B(n_6175),
.Y(n_6258)
);

AND2x2_ASAP7_75t_L g6259 ( 
.A(n_6199),
.B(n_6178),
.Y(n_6259)
);

INVx1_ASAP7_75t_L g6260 ( 
.A(n_6224),
.Y(n_6260)
);

AND2x2_ASAP7_75t_L g6261 ( 
.A(n_6200),
.B(n_6161),
.Y(n_6261)
);

INVx1_ASAP7_75t_L g6262 ( 
.A(n_6226),
.Y(n_6262)
);

NAND2xp5_ASAP7_75t_L g6263 ( 
.A(n_6221),
.B(n_6169),
.Y(n_6263)
);

NOR2xp67_ASAP7_75t_L g6264 ( 
.A(n_6230),
.B(n_6235),
.Y(n_6264)
);

INVx1_ASAP7_75t_L g6265 ( 
.A(n_6201),
.Y(n_6265)
);

OR2x2_ASAP7_75t_L g6266 ( 
.A(n_6228),
.B(n_6170),
.Y(n_6266)
);

INVx2_ASAP7_75t_L g6267 ( 
.A(n_6227),
.Y(n_6267)
);

BUFx2_ASAP7_75t_L g6268 ( 
.A(n_6227),
.Y(n_6268)
);

A2O1A1Ixp33_ASAP7_75t_L g6269 ( 
.A1(n_6213),
.A2(n_6158),
.B(n_6164),
.C(n_6153),
.Y(n_6269)
);

INVx2_ASAP7_75t_SL g6270 ( 
.A(n_6208),
.Y(n_6270)
);

AOI22xp33_ASAP7_75t_L g6271 ( 
.A1(n_6207),
.A2(n_6177),
.B1(n_6182),
.B2(n_6173),
.Y(n_6271)
);

INVx1_ASAP7_75t_L g6272 ( 
.A(n_6205),
.Y(n_6272)
);

NAND3xp33_ASAP7_75t_L g6273 ( 
.A(n_6233),
.B(n_6186),
.C(n_6183),
.Y(n_6273)
);

INVx1_ASAP7_75t_L g6274 ( 
.A(n_6243),
.Y(n_6274)
);

AND2x2_ASAP7_75t_L g6275 ( 
.A(n_6237),
.B(n_6225),
.Y(n_6275)
);

INVx1_ASAP7_75t_SL g6276 ( 
.A(n_6244),
.Y(n_6276)
);

INVx1_ASAP7_75t_SL g6277 ( 
.A(n_6244),
.Y(n_6277)
);

INVx2_ASAP7_75t_L g6278 ( 
.A(n_6254),
.Y(n_6278)
);

NAND2xp5_ASAP7_75t_L g6279 ( 
.A(n_6241),
.B(n_6195),
.Y(n_6279)
);

INVx1_ASAP7_75t_L g6280 ( 
.A(n_6260),
.Y(n_6280)
);

NAND2xp5_ASAP7_75t_L g6281 ( 
.A(n_6241),
.B(n_6230),
.Y(n_6281)
);

INVx1_ASAP7_75t_L g6282 ( 
.A(n_6256),
.Y(n_6282)
);

AOI22xp5_ASAP7_75t_L g6283 ( 
.A1(n_6239),
.A2(n_6232),
.B1(n_6214),
.B2(n_6235),
.Y(n_6283)
);

NAND2xp5_ASAP7_75t_L g6284 ( 
.A(n_6247),
.B(n_6251),
.Y(n_6284)
);

INVx2_ASAP7_75t_L g6285 ( 
.A(n_6246),
.Y(n_6285)
);

NAND2xp5_ASAP7_75t_L g6286 ( 
.A(n_6257),
.B(n_6229),
.Y(n_6286)
);

INVx1_ASAP7_75t_L g6287 ( 
.A(n_6259),
.Y(n_6287)
);

OR2x2_ASAP7_75t_L g6288 ( 
.A(n_6263),
.B(n_6185),
.Y(n_6288)
);

AND2x4_ASAP7_75t_L g6289 ( 
.A(n_6267),
.B(n_6190),
.Y(n_6289)
);

NAND2xp5_ASAP7_75t_L g6290 ( 
.A(n_6269),
.B(n_6198),
.Y(n_6290)
);

INVx2_ASAP7_75t_SL g6291 ( 
.A(n_6242),
.Y(n_6291)
);

INVx1_ASAP7_75t_L g6292 ( 
.A(n_6268),
.Y(n_6292)
);

NAND2xp5_ASAP7_75t_L g6293 ( 
.A(n_6255),
.B(n_6198),
.Y(n_6293)
);

OR2x2_ASAP7_75t_L g6294 ( 
.A(n_6263),
.B(n_6212),
.Y(n_6294)
);

INVx1_ASAP7_75t_L g6295 ( 
.A(n_6238),
.Y(n_6295)
);

INVx2_ASAP7_75t_L g6296 ( 
.A(n_6245),
.Y(n_6296)
);

NAND2xp5_ASAP7_75t_L g6297 ( 
.A(n_6270),
.B(n_6212),
.Y(n_6297)
);

NAND2xp5_ASAP7_75t_SL g6298 ( 
.A(n_6240),
.B(n_6215),
.Y(n_6298)
);

INVx1_ASAP7_75t_L g6299 ( 
.A(n_6264),
.Y(n_6299)
);

AND2x2_ASAP7_75t_L g6300 ( 
.A(n_6253),
.B(n_6215),
.Y(n_6300)
);

AND2x2_ASAP7_75t_L g6301 ( 
.A(n_6261),
.B(n_6258),
.Y(n_6301)
);

AND2x2_ASAP7_75t_L g6302 ( 
.A(n_6258),
.B(n_6262),
.Y(n_6302)
);

BUFx2_ASAP7_75t_L g6303 ( 
.A(n_6250),
.Y(n_6303)
);

INVx1_ASAP7_75t_SL g6304 ( 
.A(n_6265),
.Y(n_6304)
);

INVx1_ASAP7_75t_L g6305 ( 
.A(n_6264),
.Y(n_6305)
);

INVx2_ASAP7_75t_L g6306 ( 
.A(n_6252),
.Y(n_6306)
);

INVx3_ASAP7_75t_SL g6307 ( 
.A(n_6266),
.Y(n_6307)
);

NAND2xp5_ASAP7_75t_L g6308 ( 
.A(n_6249),
.B(n_78),
.Y(n_6308)
);

AND2x2_ASAP7_75t_L g6309 ( 
.A(n_6248),
.B(n_79),
.Y(n_6309)
);

AND2x2_ASAP7_75t_L g6310 ( 
.A(n_6249),
.B(n_79),
.Y(n_6310)
);

NAND2xp5_ASAP7_75t_L g6311 ( 
.A(n_6271),
.B(n_79),
.Y(n_6311)
);

NAND2xp5_ASAP7_75t_L g6312 ( 
.A(n_6273),
.B(n_6272),
.Y(n_6312)
);

INVx1_ASAP7_75t_L g6313 ( 
.A(n_6273),
.Y(n_6313)
);

NOR2xp33_ASAP7_75t_L g6314 ( 
.A(n_6237),
.B(n_80),
.Y(n_6314)
);

INVx1_ASAP7_75t_L g6315 ( 
.A(n_6288),
.Y(n_6315)
);

INVx1_ASAP7_75t_L g6316 ( 
.A(n_6291),
.Y(n_6316)
);

INVxp67_ASAP7_75t_L g6317 ( 
.A(n_6309),
.Y(n_6317)
);

NAND4xp25_ASAP7_75t_L g6318 ( 
.A(n_6279),
.B(n_82),
.C(n_80),
.D(n_81),
.Y(n_6318)
);

INVx1_ASAP7_75t_L g6319 ( 
.A(n_6292),
.Y(n_6319)
);

AOI22xp5_ASAP7_75t_L g6320 ( 
.A1(n_6276),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_6320)
);

AOI32xp33_ASAP7_75t_L g6321 ( 
.A1(n_6277),
.A2(n_83),
.A3(n_81),
.B1(n_82),
.B2(n_84),
.Y(n_6321)
);

AOI22xp5_ASAP7_75t_L g6322 ( 
.A1(n_6314),
.A2(n_84),
.B1(n_81),
.B2(n_83),
.Y(n_6322)
);

AND2x2_ASAP7_75t_L g6323 ( 
.A(n_6275),
.B(n_83),
.Y(n_6323)
);

NAND2xp5_ASAP7_75t_L g6324 ( 
.A(n_6310),
.B(n_83),
.Y(n_6324)
);

BUFx2_ASAP7_75t_L g6325 ( 
.A(n_6278),
.Y(n_6325)
);

OAI321xp33_ASAP7_75t_L g6326 ( 
.A1(n_6313),
.A2(n_86),
.A3(n_88),
.B1(n_84),
.B2(n_85),
.C(n_87),
.Y(n_6326)
);

AND2x2_ASAP7_75t_L g6327 ( 
.A(n_6307),
.B(n_85),
.Y(n_6327)
);

INVx1_ASAP7_75t_L g6328 ( 
.A(n_6285),
.Y(n_6328)
);

OR2x2_ASAP7_75t_L g6329 ( 
.A(n_6308),
.B(n_85),
.Y(n_6329)
);

INVx2_ASAP7_75t_L g6330 ( 
.A(n_6289),
.Y(n_6330)
);

OAI21xp5_ASAP7_75t_L g6331 ( 
.A1(n_6313),
.A2(n_86),
.B(n_87),
.Y(n_6331)
);

OR2x2_ASAP7_75t_L g6332 ( 
.A(n_6287),
.B(n_86),
.Y(n_6332)
);

INVx1_ASAP7_75t_L g6333 ( 
.A(n_6282),
.Y(n_6333)
);

OR2x2_ASAP7_75t_L g6334 ( 
.A(n_6281),
.B(n_86),
.Y(n_6334)
);

O2A1O1Ixp33_ASAP7_75t_L g6335 ( 
.A1(n_6311),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_6335)
);

AO22x1_ASAP7_75t_L g6336 ( 
.A1(n_6274),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_6336)
);

NAND2xp5_ASAP7_75t_L g6337 ( 
.A(n_6296),
.B(n_88),
.Y(n_6337)
);

AND2x2_ASAP7_75t_L g6338 ( 
.A(n_6301),
.B(n_6295),
.Y(n_6338)
);

O2A1O1Ixp33_ASAP7_75t_L g6339 ( 
.A1(n_6274),
.A2(n_91),
.B(n_89),
.C(n_90),
.Y(n_6339)
);

OAI22xp33_ASAP7_75t_SL g6340 ( 
.A1(n_6284),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_6340)
);

NAND2x1p5_ASAP7_75t_L g6341 ( 
.A(n_6298),
.B(n_90),
.Y(n_6341)
);

INVx1_ASAP7_75t_SL g6342 ( 
.A(n_6304),
.Y(n_6342)
);

HB1xp67_ASAP7_75t_L g6343 ( 
.A(n_6280),
.Y(n_6343)
);

AND2x2_ASAP7_75t_L g6344 ( 
.A(n_6300),
.B(n_6289),
.Y(n_6344)
);

INVx1_ASAP7_75t_L g6345 ( 
.A(n_6297),
.Y(n_6345)
);

INVx1_ASAP7_75t_L g6346 ( 
.A(n_6303),
.Y(n_6346)
);

OAI32xp33_ASAP7_75t_L g6347 ( 
.A1(n_6290),
.A2(n_93),
.A3(n_91),
.B1(n_92),
.B2(n_94),
.Y(n_6347)
);

OR2x6_ASAP7_75t_L g6348 ( 
.A(n_6312),
.B(n_1147),
.Y(n_6348)
);

NOR2xp33_ASAP7_75t_L g6349 ( 
.A(n_6283),
.B(n_91),
.Y(n_6349)
);

INVx1_ASAP7_75t_L g6350 ( 
.A(n_6293),
.Y(n_6350)
);

INVx2_ASAP7_75t_SL g6351 ( 
.A(n_6302),
.Y(n_6351)
);

INVx1_ASAP7_75t_SL g6352 ( 
.A(n_6294),
.Y(n_6352)
);

INVx2_ASAP7_75t_L g6353 ( 
.A(n_6306),
.Y(n_6353)
);

AOI32xp33_ASAP7_75t_L g6354 ( 
.A1(n_6299),
.A2(n_94),
.A3(n_92),
.B1(n_93),
.B2(n_95),
.Y(n_6354)
);

OAI31xp33_ASAP7_75t_L g6355 ( 
.A1(n_6341),
.A2(n_6305),
.A3(n_6286),
.B(n_95),
.Y(n_6355)
);

INVxp67_ASAP7_75t_L g6356 ( 
.A(n_6323),
.Y(n_6356)
);

NAND2xp5_ASAP7_75t_L g6357 ( 
.A(n_6336),
.B(n_93),
.Y(n_6357)
);

AOI21xp33_ASAP7_75t_L g6358 ( 
.A1(n_6316),
.A2(n_93),
.B(n_94),
.Y(n_6358)
);

AOI221xp5_ASAP7_75t_L g6359 ( 
.A1(n_6315),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.C(n_98),
.Y(n_6359)
);

INVx1_ASAP7_75t_L g6360 ( 
.A(n_6327),
.Y(n_6360)
);

INVx1_ASAP7_75t_L g6361 ( 
.A(n_6325),
.Y(n_6361)
);

AND4x1_ASAP7_75t_L g6362 ( 
.A(n_6349),
.B(n_98),
.C(n_96),
.D(n_97),
.Y(n_6362)
);

INVx1_ASAP7_75t_L g6363 ( 
.A(n_6328),
.Y(n_6363)
);

INVx2_ASAP7_75t_SL g6364 ( 
.A(n_6330),
.Y(n_6364)
);

INVx2_ASAP7_75t_SL g6365 ( 
.A(n_6344),
.Y(n_6365)
);

AOI22xp5_ASAP7_75t_L g6366 ( 
.A1(n_6351),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_6366)
);

INVx1_ASAP7_75t_SL g6367 ( 
.A(n_6342),
.Y(n_6367)
);

XOR2x2_ASAP7_75t_L g6368 ( 
.A(n_6320),
.B(n_97),
.Y(n_6368)
);

AOI22xp5_ASAP7_75t_L g6369 ( 
.A1(n_6318),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_6369)
);

AND2x2_ASAP7_75t_L g6370 ( 
.A(n_6338),
.B(n_99),
.Y(n_6370)
);

AOI22xp5_ASAP7_75t_L g6371 ( 
.A1(n_6317),
.A2(n_6352),
.B1(n_6350),
.B2(n_6319),
.Y(n_6371)
);

NAND2xp5_ASAP7_75t_L g6372 ( 
.A(n_6321),
.B(n_99),
.Y(n_6372)
);

INVx1_ASAP7_75t_L g6373 ( 
.A(n_6337),
.Y(n_6373)
);

OAI21xp5_ASAP7_75t_SL g6374 ( 
.A1(n_6346),
.A2(n_100),
.B(n_101),
.Y(n_6374)
);

INVx2_ASAP7_75t_SL g6375 ( 
.A(n_6353),
.Y(n_6375)
);

OAI22xp5_ASAP7_75t_L g6376 ( 
.A1(n_6332),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_6376)
);

AOI211xp5_ASAP7_75t_SL g6377 ( 
.A1(n_6340),
.A2(n_103),
.B(n_101),
.C(n_102),
.Y(n_6377)
);

AND2x2_ASAP7_75t_L g6378 ( 
.A(n_6348),
.B(n_101),
.Y(n_6378)
);

NAND2xp5_ASAP7_75t_L g6379 ( 
.A(n_6354),
.B(n_102),
.Y(n_6379)
);

AND2x2_ASAP7_75t_L g6380 ( 
.A(n_6348),
.B(n_6345),
.Y(n_6380)
);

INVx1_ASAP7_75t_L g6381 ( 
.A(n_6324),
.Y(n_6381)
);

INVx1_ASAP7_75t_L g6382 ( 
.A(n_6343),
.Y(n_6382)
);

INVx1_ASAP7_75t_L g6383 ( 
.A(n_6329),
.Y(n_6383)
);

OAI21xp33_ASAP7_75t_L g6384 ( 
.A1(n_6333),
.A2(n_102),
.B(n_103),
.Y(n_6384)
);

AND2x2_ASAP7_75t_L g6385 ( 
.A(n_6322),
.B(n_103),
.Y(n_6385)
);

AOI221xp5_ASAP7_75t_L g6386 ( 
.A1(n_6347),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.C(n_107),
.Y(n_6386)
);

INVx1_ASAP7_75t_SL g6387 ( 
.A(n_6334),
.Y(n_6387)
);

NAND2xp5_ASAP7_75t_SL g6388 ( 
.A(n_6335),
.B(n_104),
.Y(n_6388)
);

INVx1_ASAP7_75t_L g6389 ( 
.A(n_6339),
.Y(n_6389)
);

NOR4xp25_ASAP7_75t_L g6390 ( 
.A(n_6331),
.B(n_106),
.C(n_104),
.D(n_105),
.Y(n_6390)
);

NAND2x1p5_ASAP7_75t_L g6391 ( 
.A(n_6326),
.B(n_1060),
.Y(n_6391)
);

OAI22xp5_ASAP7_75t_L g6392 ( 
.A1(n_6316),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_6392)
);

INVx2_ASAP7_75t_L g6393 ( 
.A(n_6330),
.Y(n_6393)
);

INVxp33_ASAP7_75t_L g6394 ( 
.A(n_6327),
.Y(n_6394)
);

INVx2_ASAP7_75t_L g6395 ( 
.A(n_6330),
.Y(n_6395)
);

AND3x1_ASAP7_75t_L g6396 ( 
.A(n_6349),
.B(n_106),
.C(n_107),
.Y(n_6396)
);

XNOR2xp5_ASAP7_75t_L g6397 ( 
.A(n_6318),
.B(n_107),
.Y(n_6397)
);

AND2x2_ASAP7_75t_L g6398 ( 
.A(n_6323),
.B(n_108),
.Y(n_6398)
);

INVx1_ASAP7_75t_L g6399 ( 
.A(n_6327),
.Y(n_6399)
);

OAI22xp5_ASAP7_75t_L g6400 ( 
.A1(n_6316),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_6400)
);

AND2x2_ASAP7_75t_L g6401 ( 
.A(n_6323),
.B(n_108),
.Y(n_6401)
);

INVx1_ASAP7_75t_L g6402 ( 
.A(n_6327),
.Y(n_6402)
);

OAI21xp33_ASAP7_75t_L g6403 ( 
.A1(n_6316),
.A2(n_109),
.B(n_110),
.Y(n_6403)
);

INVx1_ASAP7_75t_L g6404 ( 
.A(n_6327),
.Y(n_6404)
);

INVx1_ASAP7_75t_L g6405 ( 
.A(n_6327),
.Y(n_6405)
);

INVx1_ASAP7_75t_L g6406 ( 
.A(n_6327),
.Y(n_6406)
);

AOI31xp33_ASAP7_75t_L g6407 ( 
.A1(n_6342),
.A2(n_112),
.A3(n_110),
.B(n_111),
.Y(n_6407)
);

NAND2xp5_ASAP7_75t_L g6408 ( 
.A(n_6336),
.B(n_110),
.Y(n_6408)
);

AOI21xp5_ASAP7_75t_L g6409 ( 
.A1(n_6357),
.A2(n_6408),
.B(n_6388),
.Y(n_6409)
);

NOR2xp33_ASAP7_75t_SL g6410 ( 
.A(n_6367),
.B(n_111),
.Y(n_6410)
);

OAI32xp33_ASAP7_75t_L g6411 ( 
.A1(n_6394),
.A2(n_113),
.A3(n_111),
.B1(n_112),
.B2(n_114),
.Y(n_6411)
);

OAI221xp5_ASAP7_75t_SL g6412 ( 
.A1(n_6371),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.C(n_114),
.Y(n_6412)
);

INVx2_ASAP7_75t_L g6413 ( 
.A(n_6364),
.Y(n_6413)
);

NOR2xp33_ASAP7_75t_L g6414 ( 
.A(n_6407),
.B(n_113),
.Y(n_6414)
);

AOI32xp33_ASAP7_75t_L g6415 ( 
.A1(n_6396),
.A2(n_115),
.A3(n_113),
.B1(n_114),
.B2(n_116),
.Y(n_6415)
);

AO211x2_ASAP7_75t_L g6416 ( 
.A1(n_6361),
.A2(n_6389),
.B(n_6363),
.C(n_6360),
.Y(n_6416)
);

AOI21xp5_ASAP7_75t_L g6417 ( 
.A1(n_6372),
.A2(n_114),
.B(n_115),
.Y(n_6417)
);

OAI22xp33_ASAP7_75t_L g6418 ( 
.A1(n_6377),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_6418)
);

AOI22xp33_ASAP7_75t_L g6419 ( 
.A1(n_6365),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_6419)
);

AND2x2_ASAP7_75t_L g6420 ( 
.A(n_6370),
.B(n_117),
.Y(n_6420)
);

O2A1O1Ixp5_ASAP7_75t_L g6421 ( 
.A1(n_6393),
.A2(n_120),
.B(n_118),
.C(n_119),
.Y(n_6421)
);

INVx1_ASAP7_75t_L g6422 ( 
.A(n_6378),
.Y(n_6422)
);

NAND2xp5_ASAP7_75t_L g6423 ( 
.A(n_6398),
.B(n_118),
.Y(n_6423)
);

AOI211xp5_ASAP7_75t_L g6424 ( 
.A1(n_6374),
.A2(n_120),
.B(n_118),
.C(n_119),
.Y(n_6424)
);

OAI32xp33_ASAP7_75t_L g6425 ( 
.A1(n_6395),
.A2(n_120),
.A3(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_6425)
);

INVx1_ASAP7_75t_L g6426 ( 
.A(n_6375),
.Y(n_6426)
);

INVx1_ASAP7_75t_L g6427 ( 
.A(n_6368),
.Y(n_6427)
);

NAND2xp5_ASAP7_75t_L g6428 ( 
.A(n_6401),
.B(n_119),
.Y(n_6428)
);

NAND2xp5_ASAP7_75t_L g6429 ( 
.A(n_6397),
.B(n_120),
.Y(n_6429)
);

INVx1_ASAP7_75t_L g6430 ( 
.A(n_6380),
.Y(n_6430)
);

INVx1_ASAP7_75t_L g6431 ( 
.A(n_6392),
.Y(n_6431)
);

NAND2xp5_ASAP7_75t_L g6432 ( 
.A(n_6369),
.B(n_121),
.Y(n_6432)
);

INVx1_ASAP7_75t_L g6433 ( 
.A(n_6400),
.Y(n_6433)
);

BUFx6f_ASAP7_75t_L g6434 ( 
.A(n_6391),
.Y(n_6434)
);

INVx1_ASAP7_75t_L g6435 ( 
.A(n_6403),
.Y(n_6435)
);

AOI22xp5_ASAP7_75t_L g6436 ( 
.A1(n_6379),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_6436)
);

AND2x2_ASAP7_75t_L g6437 ( 
.A(n_6385),
.B(n_121),
.Y(n_6437)
);

OAI221xp5_ASAP7_75t_L g6438 ( 
.A1(n_6355),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.C(n_125),
.Y(n_6438)
);

OR2x2_ASAP7_75t_L g6439 ( 
.A(n_6390),
.B(n_122),
.Y(n_6439)
);

AND2x2_ASAP7_75t_L g6440 ( 
.A(n_6356),
.B(n_122),
.Y(n_6440)
);

OAI21xp33_ASAP7_75t_L g6441 ( 
.A1(n_6399),
.A2(n_124),
.B(n_125),
.Y(n_6441)
);

INVx1_ASAP7_75t_L g6442 ( 
.A(n_6366),
.Y(n_6442)
);

INVx1_ASAP7_75t_L g6443 ( 
.A(n_6402),
.Y(n_6443)
);

AOI21xp5_ASAP7_75t_L g6444 ( 
.A1(n_6358),
.A2(n_6376),
.B(n_6384),
.Y(n_6444)
);

AND2x4_ASAP7_75t_SL g6445 ( 
.A(n_6383),
.B(n_124),
.Y(n_6445)
);

INVx2_ASAP7_75t_L g6446 ( 
.A(n_6382),
.Y(n_6446)
);

AOI211xp5_ASAP7_75t_L g6447 ( 
.A1(n_6387),
.A2(n_126),
.B(n_124),
.C(n_125),
.Y(n_6447)
);

NAND2xp5_ASAP7_75t_L g6448 ( 
.A(n_6359),
.B(n_125),
.Y(n_6448)
);

INVx1_ASAP7_75t_SL g6449 ( 
.A(n_6382),
.Y(n_6449)
);

AOI221xp5_ASAP7_75t_L g6450 ( 
.A1(n_6404),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.C(n_129),
.Y(n_6450)
);

INVx2_ASAP7_75t_L g6451 ( 
.A(n_6405),
.Y(n_6451)
);

AOI21xp33_ASAP7_75t_SL g6452 ( 
.A1(n_6406),
.A2(n_126),
.B(n_127),
.Y(n_6452)
);

OAI221xp5_ASAP7_75t_SL g6453 ( 
.A1(n_6415),
.A2(n_6373),
.B1(n_6381),
.B2(n_6386),
.C(n_6362),
.Y(n_6453)
);

AOI322xp5_ASAP7_75t_L g6454 ( 
.A1(n_6426),
.A2(n_127),
.A3(n_128),
.B1(n_129),
.B2(n_130),
.C1(n_131),
.C2(n_132),
.Y(n_6454)
);

NAND2xp33_ASAP7_75t_L g6455 ( 
.A(n_6434),
.B(n_130),
.Y(n_6455)
);

A2O1A1Ixp33_ASAP7_75t_L g6456 ( 
.A1(n_6414),
.A2(n_132),
.B(n_130),
.C(n_131),
.Y(n_6456)
);

OAI221xp5_ASAP7_75t_L g6457 ( 
.A1(n_6419),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.C(n_133),
.Y(n_6457)
);

AOI221xp5_ASAP7_75t_L g6458 ( 
.A1(n_6418),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.C(n_134),
.Y(n_6458)
);

NOR4xp25_ASAP7_75t_L g6459 ( 
.A(n_6449),
.B(n_6427),
.C(n_6413),
.D(n_6446),
.Y(n_6459)
);

AND2x2_ASAP7_75t_L g6460 ( 
.A(n_6420),
.B(n_133),
.Y(n_6460)
);

NAND3xp33_ASAP7_75t_L g6461 ( 
.A(n_6447),
.B(n_6450),
.C(n_6412),
.Y(n_6461)
);

INVxp67_ASAP7_75t_SL g6462 ( 
.A(n_6434),
.Y(n_6462)
);

NAND2xp5_ASAP7_75t_SL g6463 ( 
.A(n_6452),
.B(n_134),
.Y(n_6463)
);

INVx1_ASAP7_75t_L g6464 ( 
.A(n_6445),
.Y(n_6464)
);

OAI21xp33_ASAP7_75t_SL g6465 ( 
.A1(n_6431),
.A2(n_134),
.B(n_135),
.Y(n_6465)
);

NAND2xp5_ASAP7_75t_L g6466 ( 
.A(n_6440),
.B(n_134),
.Y(n_6466)
);

AOI221xp5_ASAP7_75t_SL g6467 ( 
.A1(n_6444),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.C(n_138),
.Y(n_6467)
);

OAI21xp33_ASAP7_75t_SL g6468 ( 
.A1(n_6433),
.A2(n_135),
.B(n_136),
.Y(n_6468)
);

NOR2xp33_ASAP7_75t_L g6469 ( 
.A(n_6410),
.B(n_135),
.Y(n_6469)
);

NAND2xp5_ASAP7_75t_L g6470 ( 
.A(n_6437),
.B(n_136),
.Y(n_6470)
);

AOI22xp5_ASAP7_75t_L g6471 ( 
.A1(n_6435),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_6471)
);

AOI21xp5_ASAP7_75t_L g6472 ( 
.A1(n_6423),
.A2(n_137),
.B(n_138),
.Y(n_6472)
);

AOI221xp5_ASAP7_75t_L g6473 ( 
.A1(n_6438),
.A2(n_140),
.B1(n_137),
.B2(n_139),
.C(n_141),
.Y(n_6473)
);

AOI21xp5_ASAP7_75t_L g6474 ( 
.A1(n_6428),
.A2(n_139),
.B(n_140),
.Y(n_6474)
);

O2A1O1Ixp33_ASAP7_75t_L g6475 ( 
.A1(n_6411),
.A2(n_141),
.B(n_139),
.C(n_140),
.Y(n_6475)
);

AOI21xp5_ASAP7_75t_L g6476 ( 
.A1(n_6429),
.A2(n_139),
.B(n_142),
.Y(n_6476)
);

AOI221xp5_ASAP7_75t_L g6477 ( 
.A1(n_6430),
.A2(n_6417),
.B1(n_6442),
.B2(n_6409),
.C(n_6421),
.Y(n_6477)
);

INVxp67_ASAP7_75t_SL g6478 ( 
.A(n_6432),
.Y(n_6478)
);

AND2x2_ASAP7_75t_L g6479 ( 
.A(n_6451),
.B(n_142),
.Y(n_6479)
);

OAI211xp5_ASAP7_75t_L g6480 ( 
.A1(n_6436),
.A2(n_144),
.B(n_142),
.C(n_143),
.Y(n_6480)
);

OAI211xp5_ASAP7_75t_SL g6481 ( 
.A1(n_6443),
.A2(n_145),
.B(n_143),
.C(n_144),
.Y(n_6481)
);

NOR3xp33_ASAP7_75t_L g6482 ( 
.A(n_6441),
.B(n_143),
.C(n_144),
.Y(n_6482)
);

NOR2xp67_ASAP7_75t_L g6483 ( 
.A(n_6439),
.B(n_144),
.Y(n_6483)
);

OAI221xp5_ASAP7_75t_L g6484 ( 
.A1(n_6424),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.C(n_148),
.Y(n_6484)
);

NOR4xp25_ASAP7_75t_SL g6485 ( 
.A(n_6422),
.B(n_147),
.C(n_145),
.D(n_146),
.Y(n_6485)
);

O2A1O1Ixp33_ASAP7_75t_L g6486 ( 
.A1(n_6448),
.A2(n_148),
.B(n_146),
.C(n_147),
.Y(n_6486)
);

INVx1_ASAP7_75t_L g6487 ( 
.A(n_6425),
.Y(n_6487)
);

AOI221xp5_ASAP7_75t_L g6488 ( 
.A1(n_6416),
.A2(n_149),
.B1(n_146),
.B2(n_147),
.C(n_150),
.Y(n_6488)
);

XNOR2xp5_ASAP7_75t_L g6489 ( 
.A(n_6416),
.B(n_149),
.Y(n_6489)
);

NOR3xp33_ASAP7_75t_L g6490 ( 
.A(n_6412),
.B(n_149),
.C(n_150),
.Y(n_6490)
);

OAI321xp33_ASAP7_75t_L g6491 ( 
.A1(n_6426),
.A2(n_150),
.A3(n_151),
.B1(n_152),
.B2(n_153),
.C(n_154),
.Y(n_6491)
);

OAI221xp5_ASAP7_75t_L g6492 ( 
.A1(n_6415),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.C(n_153),
.Y(n_6492)
);

AND2x2_ASAP7_75t_L g6493 ( 
.A(n_6420),
.B(n_151),
.Y(n_6493)
);

NAND3xp33_ASAP7_75t_SL g6494 ( 
.A(n_6424),
.B(n_152),
.C(n_153),
.Y(n_6494)
);

AOI222xp33_ASAP7_75t_L g6495 ( 
.A1(n_6426),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.C1(n_156),
.C2(n_157),
.Y(n_6495)
);

AOI31xp33_ASAP7_75t_L g6496 ( 
.A1(n_6439),
.A2(n_156),
.A3(n_154),
.B(n_155),
.Y(n_6496)
);

INVx1_ASAP7_75t_L g6497 ( 
.A(n_6413),
.Y(n_6497)
);

XOR2x2_ASAP7_75t_L g6498 ( 
.A(n_6438),
.B(n_155),
.Y(n_6498)
);

INVx2_ASAP7_75t_SL g6499 ( 
.A(n_6497),
.Y(n_6499)
);

NAND2xp5_ASAP7_75t_L g6500 ( 
.A(n_6454),
.B(n_155),
.Y(n_6500)
);

INVx1_ASAP7_75t_L g6501 ( 
.A(n_6479),
.Y(n_6501)
);

AOI22xp5_ASAP7_75t_L g6502 ( 
.A1(n_6490),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_6502)
);

NAND3xp33_ASAP7_75t_L g6503 ( 
.A(n_6495),
.B(n_156),
.C(n_157),
.Y(n_6503)
);

OAI22xp5_ASAP7_75t_L g6504 ( 
.A1(n_6461),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_6504)
);

NOR2xp67_ASAP7_75t_L g6505 ( 
.A(n_6464),
.B(n_158),
.Y(n_6505)
);

AOI22xp33_ASAP7_75t_L g6506 ( 
.A1(n_6482),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.Y(n_6506)
);

A2O1A1Ixp33_ASAP7_75t_L g6507 ( 
.A1(n_6475),
.A2(n_161),
.B(n_159),
.C(n_160),
.Y(n_6507)
);

AOI21xp33_ASAP7_75t_L g6508 ( 
.A1(n_6465),
.A2(n_159),
.B(n_160),
.Y(n_6508)
);

INVx1_ASAP7_75t_L g6509 ( 
.A(n_6462),
.Y(n_6509)
);

NOR3xp33_ASAP7_75t_L g6510 ( 
.A(n_6491),
.B(n_161),
.C(n_162),
.Y(n_6510)
);

AND4x1_ASAP7_75t_L g6511 ( 
.A(n_6459),
.B(n_163),
.C(n_161),
.D(n_162),
.Y(n_6511)
);

NOR2x1_ASAP7_75t_L g6512 ( 
.A(n_6494),
.B(n_162),
.Y(n_6512)
);

AOI21xp5_ASAP7_75t_L g6513 ( 
.A1(n_6463),
.A2(n_162),
.B(n_163),
.Y(n_6513)
);

OAI322xp33_ASAP7_75t_L g6514 ( 
.A1(n_6487),
.A2(n_163),
.A3(n_164),
.B1(n_165),
.B2(n_166),
.C1(n_167),
.C2(n_168),
.Y(n_6514)
);

AOI21xp5_ASAP7_75t_SL g6515 ( 
.A1(n_6456),
.A2(n_163),
.B(n_164),
.Y(n_6515)
);

NAND2xp5_ASAP7_75t_SL g6516 ( 
.A(n_6488),
.B(n_165),
.Y(n_6516)
);

O2A1O1Ixp33_ASAP7_75t_L g6517 ( 
.A1(n_6496),
.A2(n_168),
.B(n_166),
.C(n_167),
.Y(n_6517)
);

A2O1A1Ixp33_ASAP7_75t_L g6518 ( 
.A1(n_6469),
.A2(n_169),
.B(n_166),
.C(n_168),
.Y(n_6518)
);

AOI21xp5_ASAP7_75t_SL g6519 ( 
.A1(n_6486),
.A2(n_168),
.B(n_169),
.Y(n_6519)
);

O2A1O1Ixp33_ASAP7_75t_SL g6520 ( 
.A1(n_6466),
.A2(n_6470),
.B(n_6489),
.C(n_6477),
.Y(n_6520)
);

AOI21xp33_ASAP7_75t_SL g6521 ( 
.A1(n_6492),
.A2(n_169),
.B(n_170),
.Y(n_6521)
);

OAI211xp5_ASAP7_75t_L g6522 ( 
.A1(n_6468),
.A2(n_171),
.B(n_169),
.C(n_170),
.Y(n_6522)
);

OAI22xp5_ASAP7_75t_L g6523 ( 
.A1(n_6483),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_6523)
);

AOI322xp5_ASAP7_75t_L g6524 ( 
.A1(n_6478),
.A2(n_6467),
.A3(n_6455),
.B1(n_6473),
.B2(n_6460),
.C1(n_6493),
.C2(n_6458),
.Y(n_6524)
);

INVxp67_ASAP7_75t_L g6525 ( 
.A(n_6484),
.Y(n_6525)
);

AOI322xp5_ASAP7_75t_L g6526 ( 
.A1(n_6471),
.A2(n_170),
.A3(n_171),
.B1(n_172),
.B2(n_173),
.C1(n_174),
.C2(n_175),
.Y(n_6526)
);

AOI21xp33_ASAP7_75t_L g6527 ( 
.A1(n_6457),
.A2(n_171),
.B(n_172),
.Y(n_6527)
);

NAND2xp5_ASAP7_75t_L g6528 ( 
.A(n_6485),
.B(n_172),
.Y(n_6528)
);

AOI21xp5_ASAP7_75t_L g6529 ( 
.A1(n_6472),
.A2(n_173),
.B(n_174),
.Y(n_6529)
);

OAI32xp33_ASAP7_75t_L g6530 ( 
.A1(n_6481),
.A2(n_176),
.A3(n_173),
.B1(n_175),
.B2(n_177),
.Y(n_6530)
);

OAI21xp33_ASAP7_75t_L g6531 ( 
.A1(n_6498),
.A2(n_175),
.B(n_176),
.Y(n_6531)
);

AOI222xp33_ASAP7_75t_L g6532 ( 
.A1(n_6480),
.A2(n_175),
.B1(n_176),
.B2(n_178),
.C1(n_179),
.C2(n_180),
.Y(n_6532)
);

NOR2xp33_ASAP7_75t_L g6533 ( 
.A(n_6453),
.B(n_6474),
.Y(n_6533)
);

AOI211xp5_ASAP7_75t_L g6534 ( 
.A1(n_6476),
.A2(n_179),
.B(n_176),
.C(n_178),
.Y(n_6534)
);

NAND2x1_ASAP7_75t_SL g6535 ( 
.A(n_6479),
.B(n_178),
.Y(n_6535)
);

AOI211xp5_ASAP7_75t_L g6536 ( 
.A1(n_6459),
.A2(n_181),
.B(n_178),
.C(n_180),
.Y(n_6536)
);

OR2x2_ASAP7_75t_L g6537 ( 
.A(n_6459),
.B(n_180),
.Y(n_6537)
);

AND2x2_ASAP7_75t_L g6538 ( 
.A(n_6460),
.B(n_181),
.Y(n_6538)
);

INVx2_ASAP7_75t_SL g6539 ( 
.A(n_6509),
.Y(n_6539)
);

INVx1_ASAP7_75t_L g6540 ( 
.A(n_6537),
.Y(n_6540)
);

OAI22xp5_ASAP7_75t_L g6541 ( 
.A1(n_6502),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_6541)
);

INVx1_ASAP7_75t_L g6542 ( 
.A(n_6528),
.Y(n_6542)
);

A2O1A1Ixp33_ASAP7_75t_L g6543 ( 
.A1(n_6533),
.A2(n_185),
.B(n_182),
.C(n_184),
.Y(n_6543)
);

OAI21xp5_ASAP7_75t_L g6544 ( 
.A1(n_6503),
.A2(n_182),
.B(n_185),
.Y(n_6544)
);

INVx2_ASAP7_75t_SL g6545 ( 
.A(n_6499),
.Y(n_6545)
);

OAI21xp33_ASAP7_75t_L g6546 ( 
.A1(n_6531),
.A2(n_182),
.B(n_185),
.Y(n_6546)
);

OAI22xp5_ASAP7_75t_L g6547 ( 
.A1(n_6525),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.Y(n_6547)
);

INVxp67_ASAP7_75t_L g6548 ( 
.A(n_6512),
.Y(n_6548)
);

NAND2xp5_ASAP7_75t_L g6549 ( 
.A(n_6510),
.B(n_186),
.Y(n_6549)
);

AOI221xp5_ASAP7_75t_L g6550 ( 
.A1(n_6530),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.C(n_189),
.Y(n_6550)
);

O2A1O1Ixp33_ASAP7_75t_L g6551 ( 
.A1(n_6508),
.A2(n_189),
.B(n_187),
.C(n_188),
.Y(n_6551)
);

NOR2xp67_ASAP7_75t_L g6552 ( 
.A(n_6522),
.B(n_187),
.Y(n_6552)
);

OAI22xp5_ASAP7_75t_L g6553 ( 
.A1(n_6500),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.Y(n_6553)
);

INVxp67_ASAP7_75t_SL g6554 ( 
.A(n_6505),
.Y(n_6554)
);

CKINVDCx5p33_ASAP7_75t_R g6555 ( 
.A(n_6504),
.Y(n_6555)
);

CKINVDCx16_ASAP7_75t_R g6556 ( 
.A(n_6538),
.Y(n_6556)
);

INVx1_ASAP7_75t_L g6557 ( 
.A(n_6511),
.Y(n_6557)
);

INVx1_ASAP7_75t_L g6558 ( 
.A(n_6535),
.Y(n_6558)
);

AO22x2_ASAP7_75t_L g6559 ( 
.A1(n_6523),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.Y(n_6559)
);

NAND5xp2_ASAP7_75t_L g6560 ( 
.A(n_6524),
.B(n_190),
.C(n_191),
.D(n_192),
.E(n_193),
.Y(n_6560)
);

INVx1_ASAP7_75t_SL g6561 ( 
.A(n_6501),
.Y(n_6561)
);

OAI221xp5_ASAP7_75t_SL g6562 ( 
.A1(n_6517),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.C(n_193),
.Y(n_6562)
);

HB1xp67_ASAP7_75t_L g6563 ( 
.A(n_6516),
.Y(n_6563)
);

AOI221xp5_ASAP7_75t_L g6564 ( 
.A1(n_6514),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.C(n_194),
.Y(n_6564)
);

OA22x2_ASAP7_75t_L g6565 ( 
.A1(n_6519),
.A2(n_193),
.B1(n_191),
.B2(n_192),
.Y(n_6565)
);

OAI211xp5_ASAP7_75t_L g6566 ( 
.A1(n_6527),
.A2(n_196),
.B(n_194),
.C(n_195),
.Y(n_6566)
);

AOI221xp5_ASAP7_75t_L g6567 ( 
.A1(n_6521),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.C(n_197),
.Y(n_6567)
);

INVx1_ASAP7_75t_L g6568 ( 
.A(n_6507),
.Y(n_6568)
);

INVx2_ASAP7_75t_SL g6569 ( 
.A(n_6536),
.Y(n_6569)
);

AOI221xp5_ASAP7_75t_L g6570 ( 
.A1(n_6520),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.C(n_199),
.Y(n_6570)
);

AOI22xp5_ASAP7_75t_L g6571 ( 
.A1(n_6532),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_6571)
);

O2A1O1Ixp33_ASAP7_75t_L g6572 ( 
.A1(n_6518),
.A2(n_200),
.B(n_198),
.C(n_199),
.Y(n_6572)
);

NAND2xp5_ASAP7_75t_L g6573 ( 
.A(n_6540),
.B(n_6526),
.Y(n_6573)
);

OAI21xp33_ASAP7_75t_L g6574 ( 
.A1(n_6560),
.A2(n_6506),
.B(n_6515),
.Y(n_6574)
);

NAND3xp33_ASAP7_75t_L g6575 ( 
.A(n_6570),
.B(n_6534),
.C(n_6513),
.Y(n_6575)
);

NAND2xp5_ASAP7_75t_L g6576 ( 
.A(n_6552),
.B(n_6529),
.Y(n_6576)
);

AOI22xp5_ASAP7_75t_L g6577 ( 
.A1(n_6539),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.Y(n_6577)
);

XOR2x2_ASAP7_75t_L g6578 ( 
.A(n_6562),
.B(n_200),
.Y(n_6578)
);

INVx1_ASAP7_75t_L g6579 ( 
.A(n_6565),
.Y(n_6579)
);

NAND4xp25_ASAP7_75t_L g6580 ( 
.A(n_6564),
.B(n_203),
.C(n_201),
.D(n_202),
.Y(n_6580)
);

INVx1_ASAP7_75t_L g6581 ( 
.A(n_6557),
.Y(n_6581)
);

HB1xp67_ASAP7_75t_L g6582 ( 
.A(n_6545),
.Y(n_6582)
);

OA33x2_ASAP7_75t_L g6583 ( 
.A1(n_6553),
.A2(n_201),
.A3(n_202),
.B1(n_203),
.B2(n_204),
.B3(n_205),
.Y(n_6583)
);

AOI21xp5_ASAP7_75t_L g6584 ( 
.A1(n_6549),
.A2(n_6543),
.B(n_6551),
.Y(n_6584)
);

OAI221xp5_ASAP7_75t_L g6585 ( 
.A1(n_6567),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.C(n_204),
.Y(n_6585)
);

AOI21xp5_ASAP7_75t_L g6586 ( 
.A1(n_6547),
.A2(n_6572),
.B(n_6544),
.Y(n_6586)
);

OAI21xp5_ASAP7_75t_L g6587 ( 
.A1(n_6571),
.A2(n_6566),
.B(n_6548),
.Y(n_6587)
);

OAI211xp5_ASAP7_75t_L g6588 ( 
.A1(n_6546),
.A2(n_203),
.B(n_201),
.C(n_202),
.Y(n_6588)
);

XNOR2x1_ASAP7_75t_L g6589 ( 
.A(n_6559),
.B(n_204),
.Y(n_6589)
);

NOR3xp33_ASAP7_75t_SL g6590 ( 
.A(n_6555),
.B(n_205),
.C(n_206),
.Y(n_6590)
);

OAI21xp33_ASAP7_75t_SL g6591 ( 
.A1(n_6569),
.A2(n_6554),
.B(n_6568),
.Y(n_6591)
);

OAI31xp33_ASAP7_75t_L g6592 ( 
.A1(n_6541),
.A2(n_207),
.A3(n_205),
.B(n_206),
.Y(n_6592)
);

XOR2xp5_ASAP7_75t_L g6593 ( 
.A(n_6556),
.B(n_205),
.Y(n_6593)
);

AND2x2_ASAP7_75t_SL g6594 ( 
.A(n_6550),
.B(n_6558),
.Y(n_6594)
);

O2A1O1Ixp33_ASAP7_75t_L g6595 ( 
.A1(n_6563),
.A2(n_209),
.B(n_207),
.C(n_208),
.Y(n_6595)
);

INVx1_ASAP7_75t_L g6596 ( 
.A(n_6582),
.Y(n_6596)
);

INVx1_ASAP7_75t_SL g6597 ( 
.A(n_6581),
.Y(n_6597)
);

INVxp33_ASAP7_75t_SL g6598 ( 
.A(n_6593),
.Y(n_6598)
);

NOR2x1_ASAP7_75t_L g6599 ( 
.A(n_6580),
.B(n_6542),
.Y(n_6599)
);

INVx2_ASAP7_75t_L g6600 ( 
.A(n_6579),
.Y(n_6600)
);

AOI22xp5_ASAP7_75t_L g6601 ( 
.A1(n_6574),
.A2(n_6561),
.B1(n_6559),
.B2(n_210),
.Y(n_6601)
);

OA22x2_ASAP7_75t_L g6602 ( 
.A1(n_6577),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.Y(n_6602)
);

INVx1_ASAP7_75t_L g6603 ( 
.A(n_6578),
.Y(n_6603)
);

NOR2x1_ASAP7_75t_L g6604 ( 
.A(n_6575),
.B(n_208),
.Y(n_6604)
);

NOR2x1_ASAP7_75t_L g6605 ( 
.A(n_6589),
.B(n_209),
.Y(n_6605)
);

INVx1_ASAP7_75t_L g6606 ( 
.A(n_6595),
.Y(n_6606)
);

NAND2xp5_ASAP7_75t_L g6607 ( 
.A(n_6594),
.B(n_6590),
.Y(n_6607)
);

NOR2x1_ASAP7_75t_L g6608 ( 
.A(n_6573),
.B(n_210),
.Y(n_6608)
);

AND2x4_ASAP7_75t_L g6609 ( 
.A(n_6587),
.B(n_211),
.Y(n_6609)
);

INVx1_ASAP7_75t_SL g6610 ( 
.A(n_6576),
.Y(n_6610)
);

INVx1_ASAP7_75t_L g6611 ( 
.A(n_6588),
.Y(n_6611)
);

NOR2x1_ASAP7_75t_L g6612 ( 
.A(n_6584),
.B(n_211),
.Y(n_6612)
);

AOI22xp5_ASAP7_75t_L g6613 ( 
.A1(n_6591),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.Y(n_6613)
);

INVx1_ASAP7_75t_L g6614 ( 
.A(n_6585),
.Y(n_6614)
);

INVx2_ASAP7_75t_SL g6615 ( 
.A(n_6583),
.Y(n_6615)
);

INVx1_ASAP7_75t_L g6616 ( 
.A(n_6586),
.Y(n_6616)
);

OR2x2_ASAP7_75t_L g6617 ( 
.A(n_6592),
.B(n_211),
.Y(n_6617)
);

NOR4xp75_ASAP7_75t_L g6618 ( 
.A(n_6607),
.B(n_214),
.C(n_212),
.D(n_213),
.Y(n_6618)
);

NOR2x1_ASAP7_75t_SL g6619 ( 
.A(n_6596),
.B(n_6600),
.Y(n_6619)
);

INVx1_ASAP7_75t_L g6620 ( 
.A(n_6617),
.Y(n_6620)
);

AND2x4_ASAP7_75t_L g6621 ( 
.A(n_6597),
.B(n_212),
.Y(n_6621)
);

NOR2x1_ASAP7_75t_L g6622 ( 
.A(n_6604),
.B(n_212),
.Y(n_6622)
);

NOR2x1_ASAP7_75t_L g6623 ( 
.A(n_6612),
.B(n_213),
.Y(n_6623)
);

NAND4xp75_ASAP7_75t_L g6624 ( 
.A(n_6608),
.B(n_6599),
.C(n_6605),
.D(n_6616),
.Y(n_6624)
);

NOR2xp33_ASAP7_75t_L g6625 ( 
.A(n_6598),
.B(n_214),
.Y(n_6625)
);

INVx2_ASAP7_75t_L g6626 ( 
.A(n_6609),
.Y(n_6626)
);

INVx1_ASAP7_75t_L g6627 ( 
.A(n_6613),
.Y(n_6627)
);

AOI22xp5_ASAP7_75t_L g6628 ( 
.A1(n_6614),
.A2(n_6611),
.B1(n_6615),
.B2(n_6603),
.Y(n_6628)
);

NOR2x1_ASAP7_75t_L g6629 ( 
.A(n_6606),
.B(n_214),
.Y(n_6629)
);

INVx1_ASAP7_75t_L g6630 ( 
.A(n_6602),
.Y(n_6630)
);

NAND2xp5_ASAP7_75t_L g6631 ( 
.A(n_6601),
.B(n_214),
.Y(n_6631)
);

O2A1O1Ixp33_ASAP7_75t_L g6632 ( 
.A1(n_6610),
.A2(n_217),
.B(n_215),
.C(n_216),
.Y(n_6632)
);

XNOR2x1_ASAP7_75t_L g6633 ( 
.A(n_6604),
.B(n_215),
.Y(n_6633)
);

XNOR2xp5_ASAP7_75t_L g6634 ( 
.A(n_6596),
.B(n_215),
.Y(n_6634)
);

NAND4xp75_ASAP7_75t_L g6635 ( 
.A(n_6604),
.B(n_217),
.C(n_215),
.D(n_216),
.Y(n_6635)
);

AOI311xp33_ASAP7_75t_L g6636 ( 
.A1(n_6620),
.A2(n_216),
.A3(n_217),
.B(n_218),
.C(n_219),
.Y(n_6636)
);

AOI32xp33_ASAP7_75t_L g6637 ( 
.A1(n_6625),
.A2(n_217),
.A3(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_6637)
);

OAI22xp5_ASAP7_75t_L g6638 ( 
.A1(n_6628),
.A2(n_220),
.B1(n_218),
.B2(n_219),
.Y(n_6638)
);

OAI211xp5_ASAP7_75t_SL g6639 ( 
.A1(n_6631),
.A2(n_221),
.B(n_218),
.C(n_219),
.Y(n_6639)
);

NAND4xp25_ASAP7_75t_L g6640 ( 
.A(n_6627),
.B(n_223),
.C(n_221),
.D(n_222),
.Y(n_6640)
);

O2A1O1Ixp33_ASAP7_75t_L g6641 ( 
.A1(n_6632),
.A2(n_223),
.B(n_221),
.C(n_222),
.Y(n_6641)
);

OAI22xp5_ASAP7_75t_SL g6642 ( 
.A1(n_6634),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_6642)
);

NAND4xp25_ASAP7_75t_SL g6643 ( 
.A(n_6630),
.B(n_227),
.C(n_224),
.D(n_226),
.Y(n_6643)
);

NOR3xp33_ASAP7_75t_L g6644 ( 
.A(n_6624),
.B(n_224),
.C(n_226),
.Y(n_6644)
);

OAI21xp33_ASAP7_75t_SL g6645 ( 
.A1(n_6629),
.A2(n_6622),
.B(n_6623),
.Y(n_6645)
);

AOI22xp5_ASAP7_75t_L g6646 ( 
.A1(n_6644),
.A2(n_6626),
.B1(n_6621),
.B2(n_6633),
.Y(n_6646)
);

INVx2_ASAP7_75t_L g6647 ( 
.A(n_6638),
.Y(n_6647)
);

AND2x4_ASAP7_75t_L g6648 ( 
.A(n_6645),
.B(n_6619),
.Y(n_6648)
);

XOR2x2_ASAP7_75t_L g6649 ( 
.A(n_6642),
.B(n_6618),
.Y(n_6649)
);

INVx2_ASAP7_75t_SL g6650 ( 
.A(n_6636),
.Y(n_6650)
);

OAI21xp5_ASAP7_75t_L g6651 ( 
.A1(n_6641),
.A2(n_6621),
.B(n_6639),
.Y(n_6651)
);

NOR2x1_ASAP7_75t_L g6652 ( 
.A(n_6643),
.B(n_6635),
.Y(n_6652)
);

XOR2xp5_ASAP7_75t_L g6653 ( 
.A(n_6640),
.B(n_224),
.Y(n_6653)
);

OAI21xp33_ASAP7_75t_L g6654 ( 
.A1(n_6648),
.A2(n_6637),
.B(n_226),
.Y(n_6654)
);

INVx1_ASAP7_75t_L g6655 ( 
.A(n_6653),
.Y(n_6655)
);

INVx1_ASAP7_75t_L g6656 ( 
.A(n_6650),
.Y(n_6656)
);

INVx2_ASAP7_75t_L g6657 ( 
.A(n_6649),
.Y(n_6657)
);

INVx1_ASAP7_75t_L g6658 ( 
.A(n_6646),
.Y(n_6658)
);

INVx1_ASAP7_75t_L g6659 ( 
.A(n_6656),
.Y(n_6659)
);

INVx2_ASAP7_75t_SL g6660 ( 
.A(n_6659),
.Y(n_6660)
);

AOI21xp5_ASAP7_75t_L g6661 ( 
.A1(n_6660),
.A2(n_6651),
.B(n_6658),
.Y(n_6661)
);

AOI22xp5_ASAP7_75t_L g6662 ( 
.A1(n_6660),
.A2(n_6657),
.B1(n_6655),
.B2(n_6647),
.Y(n_6662)
);

INVx1_ASAP7_75t_L g6663 ( 
.A(n_6661),
.Y(n_6663)
);

INVx2_ASAP7_75t_L g6664 ( 
.A(n_6663),
.Y(n_6664)
);

AOI222xp33_ASAP7_75t_L g6665 ( 
.A1(n_6664),
.A2(n_6662),
.B1(n_6654),
.B2(n_6652),
.C1(n_229),
.C2(n_230),
.Y(n_6665)
);

AOI21xp5_ASAP7_75t_L g6666 ( 
.A1(n_6664),
.A2(n_226),
.B(n_227),
.Y(n_6666)
);

AOI222xp33_ASAP7_75t_L g6667 ( 
.A1(n_6665),
.A2(n_6666),
.B1(n_228),
.B2(n_229),
.C1(n_230),
.C2(n_232),
.Y(n_6667)
);

AOI22xp33_ASAP7_75t_L g6668 ( 
.A1(n_6665),
.A2(n_229),
.B1(n_227),
.B2(n_228),
.Y(n_6668)
);

OR2x6_ASAP7_75t_L g6669 ( 
.A(n_6668),
.B(n_1060),
.Y(n_6669)
);

AO21x2_ASAP7_75t_L g6670 ( 
.A1(n_6667),
.A2(n_227),
.B(n_230),
.Y(n_6670)
);

AOI21xp33_ASAP7_75t_SL g6671 ( 
.A1(n_6669),
.A2(n_1062),
.B(n_1061),
.Y(n_6671)
);

AOI211xp5_ASAP7_75t_L g6672 ( 
.A1(n_6671),
.A2(n_6670),
.B(n_234),
.C(n_230),
.Y(n_6672)
);


endmodule