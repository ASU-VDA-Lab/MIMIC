module fake_netlist_6_4109_n_1249 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1249);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1249;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_245;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_836;
wire n_375;
wire n_522;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_224;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_530;
wire n_277;
wire n_618;
wire n_199;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_210;
wire n_1069;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_1052;
wire n_462;
wire n_1033;
wire n_304;
wire n_694;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_615;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1035;
wire n_294;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_272;
wire n_526;
wire n_1183;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_552;
wire n_216;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_292;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_211;
wire n_231;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_259;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1187;
wire n_610;
wire n_1024;
wire n_198;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_218;
wire n_1213;
wire n_239;
wire n_782;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_258;
wire n_456;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_273;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1241;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_306;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_502;
wire n_672;
wire n_285;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_855;
wire n_591;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_214;
wire n_246;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1147;
wire n_763;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_911;
wire n_236;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_709;
wire n_366;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_192;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_148),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_84),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_180),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_16),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_59),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_13),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_177),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_33),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_32),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_117),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_94),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_2),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_130),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_111),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_169),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_81),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_35),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_133),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_138),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_48),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_121),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_5),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_70),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_64),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_12),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_15),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_112),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_28),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_147),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_104),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_19),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_131),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_118),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_141),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_137),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_18),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_102),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_183),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_64),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_135),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_184),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_165),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_59),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_146),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_120),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_13),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_145),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_170),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_127),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_175),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_154),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_107),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_38),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_71),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_125),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_73),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_67),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_20),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_51),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_35),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_166),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_78),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_62),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_53),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_6),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_11),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_181),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_60),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_17),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_50),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_149),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_106),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_82),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_55),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_153),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_119),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_132),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_128),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_34),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_173),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_151),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_159),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_182),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_12),
.Y(n_275)
);

HB1xp67_ASAP7_75t_SL g276 ( 
.A(n_24),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_122),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_105),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_30),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_25),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_26),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_14),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_51),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_86),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_168),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_5),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_63),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_42),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_50),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_172),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_142),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_18),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_174),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_83),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_114),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_69),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_41),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_60),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_34),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_171),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_3),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_72),
.Y(n_302)
);

BUFx10_ASAP7_75t_L g303 ( 
.A(n_80),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_109),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_32),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_196),
.Y(n_306)
);

INVxp33_ASAP7_75t_SL g307 ( 
.A(n_190),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_185),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_192),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_196),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_191),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_215),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_194),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_197),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_238),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_266),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_300),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_276),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_196),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_218),
.B(n_0),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_196),
.Y(n_321)
);

NOR2xp67_ASAP7_75t_L g322 ( 
.A(n_236),
.B(n_0),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_236),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_199),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_272),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_281),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_248),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_273),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_189),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_205),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_281),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_294),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_298),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_207),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_206),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_208),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_212),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_213),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_298),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_305),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_305),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_188),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_223),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_188),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_193),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_248),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_224),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_227),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_193),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_292),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_228),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_204),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_L g353 ( 
.A(n_204),
.B(n_1),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_209),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_209),
.Y(n_355)
);

INVxp33_ASAP7_75t_L g356 ( 
.A(n_216),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_303),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_303),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_292),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_218),
.B(n_201),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_216),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_195),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_230),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_231),
.Y(n_364)
);

NOR2xp67_ASAP7_75t_L g365 ( 
.A(n_244),
.B(n_1),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_244),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_254),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_232),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_201),
.B(n_2),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_235),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_254),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_237),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_186),
.B(n_3),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_239),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_240),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_255),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_186),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_241),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_187),
.B(n_4),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_245),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_252),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_255),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_265),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_253),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_258),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_303),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_187),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_265),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_283),
.B(n_4),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_263),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_283),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_222),
.B(n_6),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_287),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_269),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_287),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_214),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_342),
.Y(n_397)
);

OAI21x1_ASAP7_75t_L g398 ( 
.A1(n_360),
.A2(n_242),
.B(n_222),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_321),
.B(n_304),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_306),
.B(n_242),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_377),
.B(n_271),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_308),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_342),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_387),
.B(n_274),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_344),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_344),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_306),
.B(n_198),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_350),
.B(n_198),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_346),
.B(n_277),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_362),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_345),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_362),
.Y(n_412)
);

AND2x2_ASAP7_75t_R g413 ( 
.A(n_386),
.B(n_297),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_345),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_329),
.B(n_260),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_362),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_311),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_352),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_352),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_329),
.A2(n_286),
.B1(n_275),
.B2(n_373),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_362),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_318),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_362),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_320),
.B(n_278),
.Y(n_424)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_369),
.A2(n_202),
.B(n_200),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_318),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_354),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_362),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_310),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_310),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_L g431 ( 
.A(n_309),
.B(n_219),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_354),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_386),
.B(n_303),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_319),
.B(n_200),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_357),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_307),
.B(n_225),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_319),
.B(n_202),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_355),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_334),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_323),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_355),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_337),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_361),
.Y(n_443)
);

BUFx8_ASAP7_75t_L g444 ( 
.A(n_357),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_312),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_323),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_389),
.B(n_203),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_357),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_326),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_338),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_359),
.B(n_304),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_389),
.B(n_203),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_326),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_331),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_331),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_333),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_327),
.B(n_210),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_327),
.B(n_302),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_361),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_327),
.B(n_284),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_366),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_358),
.B(n_226),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_353),
.B(n_210),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_315),
.B(n_211),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_353),
.B(n_211),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_379),
.B(n_285),
.Y(n_466)
);

CKINVDCx6p67_ASAP7_75t_R g467 ( 
.A(n_426),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_410),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_447),
.A2(n_369),
.B1(n_392),
.B2(n_317),
.Y(n_469)
);

INVx4_ASAP7_75t_SL g470 ( 
.A(n_423),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_436),
.B(n_313),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_458),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_423),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_429),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_397),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_409),
.B(n_314),
.Y(n_476)
);

BUFx10_ASAP7_75t_L g477 ( 
.A(n_436),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_433),
.B(n_435),
.Y(n_478)
);

AOI21x1_ASAP7_75t_L g479 ( 
.A1(n_407),
.A2(n_392),
.B(n_365),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_397),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_429),
.Y(n_481)
);

AND2x2_ASAP7_75t_SL g482 ( 
.A(n_433),
.B(n_195),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_324),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_457),
.B(n_358),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_458),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_423),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_423),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_409),
.B(n_330),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_424),
.B(n_335),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_L g490 ( 
.A1(n_447),
.A2(n_365),
.B1(n_322),
.B2(n_301),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_348),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_403),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_403),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_457),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_429),
.Y(n_495)
);

INVxp33_ASAP7_75t_L g496 ( 
.A(n_415),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_424),
.B(n_363),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_435),
.B(n_364),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_422),
.Y(n_499)
);

NOR2x1p5_ASAP7_75t_L g500 ( 
.A(n_402),
.B(n_358),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_423),
.Y(n_501)
);

AND2x6_ASAP7_75t_L g502 ( 
.A(n_447),
.B(n_195),
.Y(n_502)
);

OAI22xp33_ASAP7_75t_L g503 ( 
.A1(n_415),
.A2(n_356),
.B1(n_229),
.B2(n_233),
.Y(n_503)
);

NAND3xp33_ASAP7_75t_L g504 ( 
.A(n_464),
.B(n_399),
.C(n_408),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_430),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_405),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_423),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_430),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_405),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_SL g510 ( 
.A1(n_444),
.A2(n_325),
.B1(n_332),
.B2(n_328),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_406),
.Y(n_511)
);

AND2x6_ASAP7_75t_L g512 ( 
.A(n_447),
.B(n_195),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_430),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_454),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_448),
.B(n_368),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_457),
.B(n_333),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_406),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_460),
.B(n_372),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_417),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_411),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_423),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_425),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_454),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_448),
.B(n_374),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_444),
.B(n_380),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_420),
.A2(n_299),
.B1(n_249),
.B2(n_270),
.Y(n_526)
);

INVx5_ASAP7_75t_L g527 ( 
.A(n_410),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_422),
.Y(n_528)
);

INVx8_ASAP7_75t_L g529 ( 
.A(n_447),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_444),
.B(n_384),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_411),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_445),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_445),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_410),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_460),
.B(n_385),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_414),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_414),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_472),
.B(n_485),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_472),
.B(n_401),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_474),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_474),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_485),
.B(n_483),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_510),
.A2(n_420),
.B1(n_496),
.B2(n_316),
.Y(n_543)
);

OAI22xp33_ASAP7_75t_L g544 ( 
.A1(n_504),
.A2(n_426),
.B1(n_442),
.B2(n_439),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_475),
.Y(n_545)
);

NAND3xp33_ASAP7_75t_L g546 ( 
.A(n_504),
.B(n_464),
.C(n_399),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_482),
.B(n_401),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_482),
.B(n_404),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_475),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_491),
.B(n_404),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_471),
.B(n_489),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_497),
.B(n_336),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_L g553 ( 
.A(n_469),
.B(n_399),
.C(n_408),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_484),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_476),
.B(n_343),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_482),
.A2(n_452),
.B1(n_465),
.B2(n_463),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_480),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_474),
.Y(n_558)
);

OAI221xp5_ASAP7_75t_L g559 ( 
.A1(n_490),
.A2(n_322),
.B1(n_408),
.B2(n_451),
.C(n_349),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_494),
.B(n_452),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_481),
.Y(n_561)
);

OAI22x1_ASAP7_75t_L g562 ( 
.A1(n_526),
.A2(n_442),
.B1(n_450),
.B2(n_439),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_494),
.B(n_452),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_494),
.B(n_452),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_477),
.B(n_444),
.Y(n_565)
);

NAND2xp33_ASAP7_75t_L g566 ( 
.A(n_502),
.B(n_195),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_480),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_484),
.B(n_451),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_481),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_492),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_488),
.B(n_347),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_529),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_481),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_518),
.B(n_452),
.Y(n_574)
);

AO22x2_ASAP7_75t_L g575 ( 
.A1(n_478),
.A2(n_522),
.B1(n_463),
.B2(n_465),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_477),
.B(n_535),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_492),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_493),
.B(n_506),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_493),
.B(n_390),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_506),
.B(n_463),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_SL g581 ( 
.A1(n_477),
.A2(n_444),
.B1(n_450),
.B2(n_431),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_477),
.B(n_451),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_509),
.B(n_463),
.Y(n_583)
);

AOI221xp5_ASAP7_75t_L g584 ( 
.A1(n_503),
.A2(n_301),
.B1(n_297),
.B2(n_250),
.C(n_280),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_509),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_522),
.A2(n_465),
.B1(n_463),
.B2(n_425),
.Y(n_586)
);

AOI22x1_ASAP7_75t_L g587 ( 
.A1(n_511),
.A2(n_465),
.B1(n_407),
.B2(n_434),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_511),
.B(n_465),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_516),
.B(n_407),
.Y(n_589)
);

INVx8_ASAP7_75t_L g590 ( 
.A(n_529),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_516),
.B(n_407),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_517),
.B(n_407),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_495),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_525),
.B(n_351),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_498),
.B(n_370),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_495),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_515),
.B(n_375),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_495),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_534),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_534),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_517),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_520),
.B(n_434),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_520),
.B(n_434),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_529),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_531),
.B(n_434),
.Y(n_605)
);

AOI221xp5_ASAP7_75t_L g606 ( 
.A1(n_526),
.A2(n_261),
.B1(n_251),
.B2(n_256),
.C(n_257),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_530),
.B(n_378),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_505),
.Y(n_608)
);

INVx8_ASAP7_75t_L g609 ( 
.A(n_529),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_524),
.B(n_381),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_531),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_536),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_536),
.B(n_394),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_537),
.A2(n_434),
.B1(n_437),
.B2(n_400),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_537),
.B(n_437),
.Y(n_615)
);

NAND2x1_ASAP7_75t_L g616 ( 
.A(n_473),
.B(n_410),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_468),
.B(n_437),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_534),
.B(n_437),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_534),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_529),
.B(n_437),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_505),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_505),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_507),
.B(n_462),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_508),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_508),
.Y(n_625)
);

O2A1O1Ixp5_ASAP7_75t_L g626 ( 
.A1(n_479),
.A2(n_462),
.B(n_400),
.C(n_296),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_508),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_513),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_499),
.B(n_396),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_528),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_507),
.B(n_400),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_507),
.B(n_400),
.Y(n_632)
);

NOR3xp33_ASAP7_75t_L g633 ( 
.A(n_528),
.B(n_279),
.C(n_259),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_507),
.B(n_400),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_519),
.B(n_290),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_502),
.B(n_512),
.Y(n_636)
);

O2A1O1Ixp33_ASAP7_75t_L g637 ( 
.A1(n_550),
.A2(n_522),
.B(n_513),
.C(n_268),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_574),
.A2(n_620),
.B(n_563),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_546),
.A2(n_425),
.B1(n_502),
.B2(n_512),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_542),
.B(n_479),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g641 ( 
.A1(n_626),
.A2(n_398),
.B(n_513),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_551),
.B(n_500),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_604),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_560),
.A2(n_486),
.B(n_473),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_552),
.Y(n_645)
);

NOR3xp33_ASAP7_75t_L g646 ( 
.A(n_555),
.B(n_532),
.C(n_533),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_586),
.A2(n_500),
.B1(n_296),
.B2(n_247),
.Y(n_647)
);

O2A1O1Ixp33_ASAP7_75t_L g648 ( 
.A1(n_547),
.A2(n_264),
.B(n_262),
.C(n_247),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_556),
.B(n_514),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_564),
.A2(n_486),
.B(n_473),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_540),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_540),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_541),
.Y(n_653)
);

A2O1A1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_546),
.A2(n_398),
.B(n_293),
.C(n_217),
.Y(n_654)
);

AND2x2_ASAP7_75t_SL g655 ( 
.A(n_565),
.B(n_217),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_630),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_541),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_580),
.A2(n_588),
.B(n_583),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_539),
.B(n_502),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_568),
.B(n_538),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_545),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_604),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_617),
.A2(n_486),
.B(n_473),
.Y(n_663)
);

AOI21x1_ASAP7_75t_L g664 ( 
.A1(n_548),
.A2(n_523),
.B(n_514),
.Y(n_664)
);

A2O1A1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_553),
.A2(n_398),
.B(n_293),
.C(n_220),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_599),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_631),
.A2(n_487),
.B(n_486),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_630),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_604),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_568),
.B(n_502),
.Y(n_670)
);

CKINVDCx10_ASAP7_75t_R g671 ( 
.A(n_543),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_554),
.B(n_502),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_632),
.A2(n_487),
.B(n_501),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_554),
.B(n_502),
.Y(n_674)
);

A2O1A1Ixp33_ASAP7_75t_L g675 ( 
.A1(n_553),
.A2(n_246),
.B(n_268),
.C(n_220),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_592),
.A2(n_523),
.B(n_514),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_634),
.A2(n_487),
.B(n_501),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_SL g678 ( 
.A(n_571),
.B(n_467),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_545),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_618),
.A2(n_487),
.B(n_501),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_543),
.Y(n_681)
);

NOR2x1_ASAP7_75t_L g682 ( 
.A(n_576),
.B(n_221),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_604),
.B(n_523),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_575),
.A2(n_264),
.B1(n_262),
.B2(n_221),
.Y(n_684)
);

A2O1A1Ixp33_ASAP7_75t_L g685 ( 
.A1(n_584),
.A2(n_246),
.B(n_234),
.C(n_243),
.Y(n_685)
);

AO21x1_ASAP7_75t_L g686 ( 
.A1(n_623),
.A2(n_243),
.B(n_234),
.Y(n_686)
);

O2A1O1Ixp5_ASAP7_75t_L g687 ( 
.A1(n_578),
.A2(n_453),
.B(n_455),
.C(n_438),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_582),
.B(n_467),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_589),
.A2(n_512),
.B1(n_502),
.B2(n_295),
.Y(n_689)
);

A2O1A1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_559),
.A2(n_427),
.B(n_418),
.C(n_419),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_589),
.B(n_512),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_602),
.A2(n_521),
.B(n_501),
.Y(n_692)
);

OAI321xp33_ASAP7_75t_L g693 ( 
.A1(n_606),
.A2(n_544),
.A3(n_629),
.B1(n_610),
.B2(n_597),
.C(n_595),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_603),
.A2(n_521),
.B(n_501),
.Y(n_694)
);

O2A1O1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_549),
.A2(n_443),
.B(n_461),
.C(n_459),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_591),
.B(n_512),
.Y(n_696)
);

A2O1A1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_549),
.A2(n_427),
.B(n_418),
.C(n_419),
.Y(n_697)
);

AOI33xp33_ASAP7_75t_L g698 ( 
.A1(n_581),
.A2(n_371),
.A3(n_366),
.B1(n_395),
.B2(n_393),
.B3(n_391),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_613),
.B(n_432),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_591),
.B(n_512),
.Y(n_700)
);

OR2x6_ASAP7_75t_SL g701 ( 
.A(n_579),
.B(n_282),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_599),
.Y(n_702)
);

O2A1O1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_557),
.A2(n_441),
.B(n_461),
.C(n_459),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_L g704 ( 
.A1(n_605),
.A2(n_512),
.B(n_421),
.Y(n_704)
);

NOR2xp67_ASAP7_75t_L g705 ( 
.A(n_635),
.B(n_432),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_615),
.A2(n_521),
.B(n_501),
.Y(n_706)
);

OAI21xp5_ASAP7_75t_L g707 ( 
.A1(n_614),
.A2(n_512),
.B(n_421),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_599),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_557),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_567),
.B(n_521),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_567),
.B(n_521),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_590),
.A2(n_521),
.B(n_416),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_570),
.B(n_453),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_570),
.B(n_453),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_590),
.A2(n_416),
.B(n_410),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_577),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_633),
.B(n_438),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_577),
.Y(n_718)
);

OAI21xp5_ASAP7_75t_L g719 ( 
.A1(n_614),
.A2(n_421),
.B(n_412),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_590),
.A2(n_416),
.B(n_412),
.Y(n_720)
);

OAI21xp5_ASAP7_75t_L g721 ( 
.A1(n_585),
.A2(n_428),
.B(n_412),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_585),
.B(n_453),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_590),
.A2(n_416),
.B(n_428),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_601),
.B(n_453),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_604),
.B(n_470),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_590),
.A2(n_416),
.B(n_428),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_601),
.B(n_455),
.Y(n_727)
);

O2A1O1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_611),
.A2(n_441),
.B(n_443),
.C(n_455),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_611),
.B(n_455),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_612),
.B(n_455),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_612),
.A2(n_527),
.B(n_456),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_562),
.Y(n_732)
);

AO21x1_ASAP7_75t_L g733 ( 
.A1(n_565),
.A2(n_383),
.B(n_395),
.Y(n_733)
);

O2A1O1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_693),
.A2(n_594),
.B(n_607),
.C(n_566),
.Y(n_734)
);

OAI21xp33_ASAP7_75t_L g735 ( 
.A1(n_645),
.A2(n_562),
.B(n_289),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_699),
.B(n_575),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_R g737 ( 
.A(n_678),
.B(n_600),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_660),
.B(n_600),
.Y(n_738)
);

BUFx8_ASAP7_75t_L g739 ( 
.A(n_656),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_651),
.Y(n_740)
);

NOR2x1_ASAP7_75t_L g741 ( 
.A(n_642),
.B(n_572),
.Y(n_741)
);

INVx4_ASAP7_75t_L g742 ( 
.A(n_643),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_661),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_SL g744 ( 
.A1(n_637),
.A2(n_600),
.B(n_619),
.C(n_627),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_668),
.B(n_572),
.Y(n_745)
);

O2A1O1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_685),
.A2(n_675),
.B(n_690),
.C(n_732),
.Y(n_746)
);

O2A1O1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_685),
.A2(n_566),
.B(n_621),
.C(n_624),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_681),
.B(n_619),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_679),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_643),
.Y(n_750)
);

OR2x6_ASAP7_75t_L g751 ( 
.A(n_643),
.B(n_609),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_709),
.B(n_619),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_717),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_688),
.B(n_609),
.Y(n_754)
);

BUFx2_ASAP7_75t_L g755 ( 
.A(n_701),
.Y(n_755)
);

NAND2x1p5_ASAP7_75t_L g756 ( 
.A(n_643),
.B(n_616),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_716),
.B(n_575),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_651),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_688),
.B(n_621),
.Y(n_759)
);

AO32x1_ASAP7_75t_L g760 ( 
.A1(n_684),
.A2(n_624),
.A3(n_625),
.B1(n_627),
.B2(n_622),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_718),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_638),
.A2(n_609),
.B(n_636),
.Y(n_762)
);

O2A1O1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_675),
.A2(n_625),
.B(n_628),
.C(n_622),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_671),
.B(n_558),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_658),
.B(n_575),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_652),
.Y(n_766)
);

OAI21x1_ASAP7_75t_L g767 ( 
.A1(n_664),
.A2(n_587),
.B(n_616),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_SL g768 ( 
.A(n_662),
.B(n_609),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_646),
.B(n_705),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_682),
.B(n_367),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_640),
.A2(n_609),
.B(n_587),
.Y(n_771)
);

BUFx2_ASAP7_75t_L g772 ( 
.A(n_662),
.Y(n_772)
);

NAND2xp33_ASAP7_75t_SL g773 ( 
.A(n_662),
.B(n_291),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_702),
.B(n_708),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_R g775 ( 
.A(n_662),
.B(n_413),
.Y(n_775)
);

AO21x1_ASAP7_75t_L g776 ( 
.A1(n_647),
.A2(n_561),
.B(n_558),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_690),
.B(n_561),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_669),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_702),
.B(n_569),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_640),
.A2(n_573),
.B(n_569),
.Y(n_780)
);

INVx5_ASAP7_75t_L g781 ( 
.A(n_669),
.Y(n_781)
);

AO21x1_ASAP7_75t_L g782 ( 
.A1(n_648),
.A2(n_593),
.B(n_573),
.Y(n_782)
);

AOI21x1_ASAP7_75t_L g783 ( 
.A1(n_683),
.A2(n_628),
.B(n_596),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_698),
.A2(n_608),
.B(n_598),
.C(n_596),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_708),
.B(n_593),
.Y(n_785)
);

A2O1A1Ixp33_ASAP7_75t_SL g786 ( 
.A1(n_731),
.A2(n_608),
.B(n_598),
.C(n_391),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_655),
.A2(n_288),
.B1(n_382),
.B2(n_367),
.Y(n_787)
);

OR2x6_ASAP7_75t_L g788 ( 
.A(n_669),
.B(n_413),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_663),
.A2(n_527),
.B(n_470),
.Y(n_789)
);

BUFx3_ASAP7_75t_L g790 ( 
.A(n_669),
.Y(n_790)
);

BUFx2_ASAP7_75t_L g791 ( 
.A(n_697),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_641),
.A2(n_527),
.B(n_195),
.Y(n_792)
);

O2A1O1Ixp5_ASAP7_75t_L g793 ( 
.A1(n_733),
.A2(n_446),
.B(n_440),
.C(n_456),
.Y(n_793)
);

O2A1O1Ixp33_ASAP7_75t_SL g794 ( 
.A1(n_665),
.A2(n_383),
.B(n_371),
.C(n_376),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_652),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_670),
.A2(n_440),
.B1(n_456),
.B2(n_449),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_655),
.B(n_470),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_639),
.A2(n_388),
.B1(n_376),
.B2(n_382),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_753),
.B(n_659),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_743),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_751),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_740),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_749),
.Y(n_803)
);

BUFx4_ASAP7_75t_SL g804 ( 
.A(n_788),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_748),
.B(n_698),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_765),
.A2(n_649),
.B(n_691),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_761),
.Y(n_807)
);

AO31x2_ASAP7_75t_L g808 ( 
.A1(n_776),
.A2(n_654),
.A3(n_686),
.B(n_665),
.Y(n_808)
);

O2A1O1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_734),
.A2(n_735),
.B(n_787),
.C(n_746),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_758),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_762),
.A2(n_650),
.B(n_644),
.Y(n_811)
);

NOR2x1_ASAP7_75t_L g812 ( 
.A(n_790),
.B(n_666),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_759),
.B(n_695),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_764),
.B(n_697),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_771),
.A2(n_649),
.B(n_680),
.Y(n_815)
);

OAI21x1_ASAP7_75t_L g816 ( 
.A1(n_767),
.A2(n_676),
.B(n_692),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_739),
.Y(n_817)
);

OAI21x1_ASAP7_75t_L g818 ( 
.A1(n_780),
.A2(n_706),
.B(n_694),
.Y(n_818)
);

OAI21x1_ASAP7_75t_L g819 ( 
.A1(n_783),
.A2(n_677),
.B(n_673),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_765),
.A2(n_667),
.B(n_721),
.Y(n_820)
);

INVx5_ASAP7_75t_L g821 ( 
.A(n_751),
.Y(n_821)
);

AO31x2_ASAP7_75t_L g822 ( 
.A1(n_782),
.A2(n_654),
.A3(n_711),
.B(n_710),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_739),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_769),
.A2(n_696),
.B1(n_700),
.B2(n_672),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_738),
.B(n_703),
.Y(n_825)
);

OAI21x1_ASAP7_75t_L g826 ( 
.A1(n_792),
.A2(n_712),
.B(n_720),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_738),
.A2(n_687),
.B(n_707),
.Y(n_827)
);

NAND3xp33_ASAP7_75t_L g828 ( 
.A(n_787),
.B(n_728),
.C(n_689),
.Y(n_828)
);

INVx5_ASAP7_75t_L g829 ( 
.A(n_751),
.Y(n_829)
);

AOI211x1_ASAP7_75t_L g830 ( 
.A1(n_757),
.A2(n_719),
.B(n_674),
.C(n_727),
.Y(n_830)
);

OAI21x1_ASAP7_75t_L g831 ( 
.A1(n_792),
.A2(n_683),
.B(n_723),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_SL g832 ( 
.A1(n_754),
.A2(n_704),
.B(n_715),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_755),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_770),
.B(n_653),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_SL g835 ( 
.A1(n_757),
.A2(n_730),
.B(n_729),
.C(n_713),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_SL g836 ( 
.A1(n_744),
.A2(n_724),
.B(n_722),
.C(n_714),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_745),
.B(n_725),
.Y(n_837)
);

OAI21x1_ASAP7_75t_L g838 ( 
.A1(n_793),
.A2(n_726),
.B(n_639),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_745),
.B(n_725),
.Y(n_839)
);

AOI211x1_ASAP7_75t_L g840 ( 
.A1(n_736),
.A2(n_388),
.B(n_393),
.C(n_341),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_777),
.A2(n_657),
.B(n_653),
.Y(n_841)
);

OAI21x1_ASAP7_75t_L g842 ( 
.A1(n_789),
.A2(n_657),
.B(n_440),
.Y(n_842)
);

OAI21x1_ASAP7_75t_L g843 ( 
.A1(n_763),
.A2(n_449),
.B(n_446),
.Y(n_843)
);

OR2x6_ASAP7_75t_L g844 ( 
.A(n_788),
.B(n_267),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_L g845 ( 
.A1(n_777),
.A2(n_446),
.B(n_449),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_788),
.B(n_339),
.Y(n_846)
);

AO31x2_ASAP7_75t_L g847 ( 
.A1(n_791),
.A2(n_339),
.A3(n_340),
.B(n_341),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_786),
.A2(n_470),
.B(n_267),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_752),
.A2(n_267),
.B1(n_340),
.B2(n_527),
.Y(n_849)
);

AOI31xp67_ASAP7_75t_L g850 ( 
.A1(n_796),
.A2(n_470),
.A3(n_267),
.B(n_454),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_752),
.B(n_454),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_SL g852 ( 
.A(n_742),
.B(n_267),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_747),
.A2(n_527),
.B(n_267),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_741),
.B(n_454),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_800),
.Y(n_855)
);

NAND2x1p5_ASAP7_75t_L g856 ( 
.A(n_821),
.B(n_781),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_821),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_803),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_814),
.A2(n_773),
.B1(n_797),
.B2(n_768),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_813),
.A2(n_798),
.B1(n_775),
.B2(n_737),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_811),
.A2(n_760),
.B(n_781),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_SL g862 ( 
.A1(n_805),
.A2(n_798),
.B1(n_781),
.B2(n_774),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_799),
.B(n_795),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_833),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_824),
.A2(n_781),
.B1(n_785),
.B2(n_766),
.Y(n_865)
);

BUFx10_ASAP7_75t_L g866 ( 
.A(n_807),
.Y(n_866)
);

INVx6_ASAP7_75t_L g867 ( 
.A(n_821),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_821),
.Y(n_868)
);

OAI22xp33_ASAP7_75t_L g869 ( 
.A1(n_844),
.A2(n_779),
.B1(n_772),
.B2(n_742),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_828),
.A2(n_779),
.B1(n_454),
.B2(n_778),
.Y(n_870)
);

BUFx2_ASAP7_75t_SL g871 ( 
.A(n_823),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_846),
.B(n_750),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_802),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_844),
.A2(n_784),
.B1(n_756),
.B2(n_778),
.Y(n_874)
);

CKINVDCx16_ASAP7_75t_R g875 ( 
.A(n_823),
.Y(n_875)
);

BUFx2_ASAP7_75t_L g876 ( 
.A(n_837),
.Y(n_876)
);

OAI22xp33_ASAP7_75t_L g877 ( 
.A1(n_844),
.A2(n_778),
.B1(n_750),
.B2(n_756),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_810),
.Y(n_878)
);

INVx6_ASAP7_75t_L g879 ( 
.A(n_829),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_825),
.A2(n_454),
.B1(n_750),
.B2(n_794),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_SL g881 ( 
.A1(n_852),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_829),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_802),
.Y(n_883)
);

INVx6_ASAP7_75t_L g884 ( 
.A(n_829),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_806),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_847),
.Y(n_886)
);

BUFx12f_ASAP7_75t_L g887 ( 
.A(n_817),
.Y(n_887)
);

BUFx8_ASAP7_75t_L g888 ( 
.A(n_837),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_829),
.Y(n_889)
);

CKINVDCx11_ASAP7_75t_R g890 ( 
.A(n_833),
.Y(n_890)
);

CKINVDCx6p67_ASAP7_75t_R g891 ( 
.A(n_837),
.Y(n_891)
);

INVxp67_ASAP7_75t_SL g892 ( 
.A(n_841),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_SL g893 ( 
.A1(n_804),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.Y(n_893)
);

INVx4_ASAP7_75t_SL g894 ( 
.A(n_847),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_SL g895 ( 
.A1(n_804),
.A2(n_10),
.B1(n_15),
.B2(n_16),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_847),
.Y(n_896)
);

OAI22x1_ASAP7_75t_L g897 ( 
.A1(n_801),
.A2(n_760),
.B1(n_19),
.B2(n_20),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_847),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_834),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_839),
.B(n_17),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_839),
.B(n_801),
.Y(n_901)
);

AND2x4_ASAP7_75t_SL g902 ( 
.A(n_839),
.B(n_812),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_840),
.Y(n_903)
);

INVx4_ASAP7_75t_L g904 ( 
.A(n_809),
.Y(n_904)
);

CKINVDCx14_ASAP7_75t_R g905 ( 
.A(n_854),
.Y(n_905)
);

INVx5_ASAP7_75t_L g906 ( 
.A(n_832),
.Y(n_906)
);

CKINVDCx6p67_ASAP7_75t_R g907 ( 
.A(n_851),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_822),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_820),
.A2(n_760),
.B(n_527),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_843),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_827),
.A2(n_835),
.B1(n_815),
.B2(n_849),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_835),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_886),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_896),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_898),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_908),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_906),
.Y(n_917)
);

OAI21x1_ASAP7_75t_L g918 ( 
.A1(n_861),
.A2(n_826),
.B(n_818),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_910),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_894),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_894),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_894),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_883),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_873),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_890),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_892),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_906),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_904),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_904),
.B(n_808),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_892),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_855),
.Y(n_931)
);

OR2x6_ASAP7_75t_L g932 ( 
.A(n_868),
.B(n_826),
.Y(n_932)
);

OAI21x1_ASAP7_75t_L g933 ( 
.A1(n_909),
.A2(n_818),
.B(n_819),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_858),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_878),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_903),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_906),
.Y(n_937)
);

OAI21x1_ASAP7_75t_L g938 ( 
.A1(n_911),
.A2(n_819),
.B(n_816),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_906),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_860),
.B(n_830),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_876),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_897),
.Y(n_942)
);

O2A1O1Ixp5_ASAP7_75t_L g943 ( 
.A1(n_865),
.A2(n_853),
.B(n_845),
.C(n_848),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_899),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_901),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_907),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_912),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_866),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_866),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_863),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_921),
.B(n_857),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_940),
.A2(n_860),
.B1(n_905),
.B2(n_885),
.Y(n_952)
);

OA21x2_ASAP7_75t_L g953 ( 
.A1(n_918),
.A2(n_933),
.B(n_938),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_943),
.A2(n_877),
.B(n_885),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_923),
.Y(n_955)
);

OR2x6_ASAP7_75t_L g956 ( 
.A(n_927),
.B(n_867),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_928),
.B(n_905),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_947),
.A2(n_881),
.B(n_859),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_947),
.A2(n_881),
.B(n_895),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_SL g960 ( 
.A1(n_940),
.A2(n_877),
.B(n_869),
.C(n_874),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_945),
.B(n_872),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_925),
.Y(n_962)
);

AOI221xp5_ASAP7_75t_L g963 ( 
.A1(n_947),
.A2(n_895),
.B1(n_893),
.B2(n_900),
.C(n_862),
.Y(n_963)
);

INVxp67_ASAP7_75t_SL g964 ( 
.A(n_928),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_943),
.A2(n_893),
.B(n_862),
.C(n_880),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_943),
.A2(n_880),
.B(n_870),
.C(n_831),
.Y(n_966)
);

NOR2x1_ASAP7_75t_SL g967 ( 
.A(n_928),
.B(n_882),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_945),
.B(n_864),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_946),
.A2(n_875),
.B1(n_891),
.B2(n_871),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_921),
.B(n_922),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_928),
.A2(n_869),
.B(n_870),
.Y(n_971)
);

OAI211xp5_ASAP7_75t_SL g972 ( 
.A1(n_942),
.A2(n_890),
.B(n_836),
.C(n_887),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_942),
.A2(n_838),
.B(n_889),
.C(n_857),
.Y(n_973)
);

AO21x2_ASAP7_75t_L g974 ( 
.A1(n_918),
.A2(n_838),
.B(n_842),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_931),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_945),
.B(n_950),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_921),
.B(n_889),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_941),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_946),
.A2(n_888),
.B1(n_884),
.B2(n_867),
.Y(n_979)
);

OR2x6_ASAP7_75t_L g980 ( 
.A(n_920),
.B(n_867),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_945),
.B(n_902),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_950),
.B(n_926),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_921),
.B(n_922),
.Y(n_983)
);

AOI21x1_ASAP7_75t_L g984 ( 
.A1(n_946),
.A2(n_843),
.B(n_850),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_948),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_948),
.A2(n_856),
.B(n_868),
.Y(n_986)
);

AO32x2_ASAP7_75t_L g987 ( 
.A1(n_917),
.A2(n_808),
.A3(n_822),
.B1(n_836),
.B2(n_902),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_931),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_948),
.A2(n_856),
.B(n_884),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_975),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_970),
.B(n_922),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_976),
.B(n_926),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_982),
.B(n_926),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_985),
.B(n_930),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_978),
.B(n_950),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_955),
.B(n_916),
.Y(n_996)
);

OR2x2_ASAP7_75t_L g997 ( 
.A(n_955),
.B(n_916),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_985),
.B(n_930),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_988),
.B(n_930),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_952),
.A2(n_942),
.B1(n_929),
.B2(n_925),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_970),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_964),
.B(n_950),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_970),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_983),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_979),
.B(n_948),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_983),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_983),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_956),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_953),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_961),
.B(n_919),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_R g1011 ( 
.A(n_962),
.B(n_888),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_987),
.Y(n_1012)
);

INVx2_ASAP7_75t_SL g1013 ( 
.A(n_980),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_973),
.B(n_919),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_1005),
.B(n_962),
.Y(n_1015)
);

OAI221xp5_ASAP7_75t_L g1016 ( 
.A1(n_1000),
.A2(n_959),
.B1(n_958),
.B2(n_963),
.C(n_965),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_992),
.B(n_929),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_990),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_1008),
.B(n_1011),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_1003),
.B(n_973),
.Y(n_1020)
);

NOR2x1p5_ASAP7_75t_L g1021 ( 
.A(n_1008),
.B(n_949),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_996),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_1003),
.B(n_953),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_1008),
.Y(n_1024)
);

INVx2_ASAP7_75t_SL g1025 ( 
.A(n_991),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1001),
.B(n_981),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_992),
.B(n_929),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_1004),
.B(n_953),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_1000),
.A2(n_965),
.B1(n_954),
.B2(n_929),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_1004),
.B(n_919),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1006),
.B(n_1007),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1006),
.B(n_920),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_990),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_996),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_1014),
.A2(n_971),
.B1(n_957),
.B2(n_980),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_1022),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_1024),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_1025),
.B(n_1001),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1025),
.B(n_1023),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1025),
.B(n_1012),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1024),
.B(n_1021),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1023),
.B(n_1012),
.Y(n_1042)
);

OR2x2_ASAP7_75t_L g1043 ( 
.A(n_1034),
.B(n_1014),
.Y(n_1043)
);

NOR2x1p5_ASAP7_75t_L g1044 ( 
.A(n_1024),
.B(n_1008),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_1021),
.B(n_1007),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1018),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1018),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_1036),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1046),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_1044),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_1039),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1036),
.B(n_1034),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1044),
.B(n_1020),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_1043),
.B(n_1017),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_1041),
.B(n_1020),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_1054),
.B(n_1043),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1050),
.B(n_1041),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1050),
.Y(n_1058)
);

OR2x2_ASAP7_75t_L g1059 ( 
.A(n_1054),
.B(n_1037),
.Y(n_1059)
);

INVx4_ASAP7_75t_L g1060 ( 
.A(n_1048),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_1060),
.A2(n_1016),
.B(n_1029),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_1057),
.A2(n_1016),
.B(n_1019),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1060),
.B(n_1055),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1056),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_1058),
.A2(n_1015),
.B(n_1029),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1059),
.Y(n_1066)
);

OAI221xp5_ASAP7_75t_L g1067 ( 
.A1(n_1057),
.A2(n_1053),
.B1(n_1052),
.B2(n_1051),
.C(n_1055),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1060),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1060),
.B(n_1053),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1060),
.Y(n_1070)
);

AO221x1_ASAP7_75t_L g1071 ( 
.A1(n_1058),
.A2(n_1037),
.B1(n_1051),
.B2(n_1049),
.C(n_1035),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1068),
.B(n_1037),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1070),
.B(n_1037),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1063),
.Y(n_1074)
);

OAI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_1061),
.A2(n_1035),
.B1(n_1008),
.B2(n_969),
.Y(n_1075)
);

OAI21xp33_ASAP7_75t_SL g1076 ( 
.A1(n_1071),
.A2(n_1039),
.B(n_1049),
.Y(n_1076)
);

AOI32xp33_ASAP7_75t_L g1077 ( 
.A1(n_1069),
.A2(n_1045),
.A3(n_1039),
.B1(n_1020),
.B2(n_1038),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_1061),
.A2(n_1008),
.B1(n_972),
.B2(n_957),
.Y(n_1078)
);

NAND3xp33_ASAP7_75t_L g1079 ( 
.A(n_1066),
.B(n_949),
.C(n_960),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1064),
.Y(n_1080)
);

AOI21xp33_ASAP7_75t_L g1081 ( 
.A1(n_1067),
.A2(n_1047),
.B(n_1046),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1062),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_1065),
.B(n_1047),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_1061),
.B(n_1045),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_1063),
.Y(n_1085)
);

OAI221xp5_ASAP7_75t_SL g1086 ( 
.A1(n_1061),
.A2(n_966),
.B1(n_1042),
.B2(n_956),
.C(n_1040),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1064),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_1076),
.A2(n_1042),
.B(n_1038),
.C(n_1040),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1085),
.B(n_1042),
.Y(n_1089)
);

XNOR2xp5_ASAP7_75t_L g1090 ( 
.A(n_1082),
.B(n_21),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1074),
.Y(n_1091)
);

NAND2x1p5_ASAP7_75t_L g1092 ( 
.A(n_1080),
.B(n_882),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1087),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1083),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_1084),
.B(n_1038),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1072),
.Y(n_1096)
);

INVxp33_ASAP7_75t_L g1097 ( 
.A(n_1073),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1078),
.B(n_1040),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_1079),
.Y(n_1099)
);

AO22x2_ASAP7_75t_L g1100 ( 
.A1(n_1075),
.A2(n_1033),
.B1(n_949),
.B2(n_1009),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1081),
.Y(n_1101)
);

INVxp67_ASAP7_75t_SL g1102 ( 
.A(n_1075),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_1086),
.B(n_1031),
.Y(n_1103)
);

XNOR2xp5_ASAP7_75t_L g1104 ( 
.A(n_1077),
.B(n_22),
.Y(n_1104)
);

AOI21xp33_ASAP7_75t_L g1105 ( 
.A1(n_1086),
.A2(n_949),
.B(n_986),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1085),
.B(n_1031),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_1089),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1089),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_1091),
.Y(n_1109)
);

NAND4xp25_ASAP7_75t_L g1110 ( 
.A(n_1101),
.B(n_960),
.C(n_989),
.D(n_968),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_1088),
.B(n_1013),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_1097),
.B(n_1033),
.Y(n_1112)
);

AND2x2_ASAP7_75t_SL g1113 ( 
.A(n_1094),
.B(n_1091),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_1097),
.B(n_1031),
.Y(n_1114)
);

NAND3xp33_ASAP7_75t_L g1115 ( 
.A(n_1104),
.B(n_944),
.C(n_995),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1102),
.B(n_1023),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_1096),
.B(n_1026),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1094),
.A2(n_966),
.B(n_956),
.C(n_1013),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1095),
.B(n_1026),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_1099),
.A2(n_944),
.B(n_24),
.C(n_25),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1090),
.B(n_1032),
.Y(n_1121)
);

NAND3xp33_ASAP7_75t_L g1122 ( 
.A(n_1104),
.B(n_944),
.C(n_950),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1090),
.B(n_1028),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1107),
.B(n_1093),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1113),
.A2(n_1100),
.B(n_1092),
.Y(n_1125)
);

AOI221xp5_ASAP7_75t_L g1126 ( 
.A1(n_1115),
.A2(n_1100),
.B1(n_1098),
.B2(n_1103),
.C(n_1105),
.Y(n_1126)
);

AOI221xp5_ASAP7_75t_L g1127 ( 
.A1(n_1122),
.A2(n_1100),
.B1(n_1098),
.B2(n_1106),
.C(n_1092),
.Y(n_1127)
);

OAI32xp33_ASAP7_75t_L g1128 ( 
.A1(n_1116),
.A2(n_1106),
.A3(n_1100),
.B1(n_1017),
.B2(n_1027),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1108),
.Y(n_1129)
);

NAND4xp25_ASAP7_75t_L g1130 ( 
.A(n_1109),
.B(n_1032),
.C(n_937),
.D(n_1027),
.Y(n_1130)
);

AOI211xp5_ASAP7_75t_L g1131 ( 
.A1(n_1120),
.A2(n_882),
.B(n_1032),
.C(n_27),
.Y(n_1131)
);

NOR3xp33_ASAP7_75t_SL g1132 ( 
.A(n_1121),
.B(n_23),
.C(n_26),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1117),
.A2(n_951),
.B1(n_977),
.B2(n_1028),
.Y(n_1133)
);

AOI221xp5_ASAP7_75t_SL g1134 ( 
.A1(n_1123),
.A2(n_1028),
.B1(n_28),
.B2(n_29),
.C(n_30),
.Y(n_1134)
);

NAND3xp33_ASAP7_75t_L g1135 ( 
.A(n_1111),
.B(n_935),
.C(n_931),
.Y(n_1135)
);

NAND4xp75_ASAP7_75t_L g1136 ( 
.A(n_1114),
.B(n_27),
.C(n_29),
.D(n_31),
.Y(n_1136)
);

OAI221xp5_ASAP7_75t_L g1137 ( 
.A1(n_1110),
.A2(n_980),
.B1(n_937),
.B2(n_884),
.C(n_879),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1112),
.A2(n_1002),
.B(n_999),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1119),
.B(n_1030),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1118),
.A2(n_980),
.B1(n_1030),
.B2(n_1009),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_L g1141 ( 
.A(n_1110),
.B(n_935),
.C(n_934),
.Y(n_1141)
);

NOR4xp25_ASAP7_75t_L g1142 ( 
.A(n_1107),
.B(n_31),
.C(n_33),
.D(n_36),
.Y(n_1142)
);

NAND4xp25_ASAP7_75t_L g1143 ( 
.A(n_1107),
.B(n_937),
.C(n_1002),
.D(n_951),
.Y(n_1143)
);

AOI211xp5_ASAP7_75t_SL g1144 ( 
.A1(n_1108),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1107),
.B(n_1010),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_1107),
.B(n_37),
.Y(n_1146)
);

OAI211xp5_ASAP7_75t_SL g1147 ( 
.A1(n_1107),
.A2(n_39),
.B(n_40),
.C(n_41),
.Y(n_1147)
);

AOI211xp5_ASAP7_75t_L g1148 ( 
.A1(n_1147),
.A2(n_1142),
.B(n_1126),
.C(n_1124),
.Y(n_1148)
);

NOR2x1_ASAP7_75t_L g1149 ( 
.A(n_1136),
.B(n_39),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1146),
.A2(n_951),
.B1(n_977),
.B2(n_991),
.Y(n_1150)
);

AOI221xp5_ASAP7_75t_L g1151 ( 
.A1(n_1127),
.A2(n_935),
.B1(n_934),
.B2(n_1009),
.C(n_993),
.Y(n_1151)
);

OAI321xp33_ASAP7_75t_L g1152 ( 
.A1(n_1129),
.A2(n_882),
.A3(n_927),
.B1(n_917),
.B2(n_934),
.C(n_920),
.Y(n_1152)
);

NOR3xp33_ASAP7_75t_L g1153 ( 
.A(n_1131),
.B(n_40),
.C(n_42),
.Y(n_1153)
);

OAI211xp5_ASAP7_75t_SL g1154 ( 
.A1(n_1132),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1145),
.Y(n_1155)
);

OAI211xp5_ASAP7_75t_L g1156 ( 
.A1(n_1134),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_1156)
);

OAI311xp33_ASAP7_75t_L g1157 ( 
.A1(n_1130),
.A2(n_46),
.A3(n_47),
.B1(n_48),
.C1(n_49),
.Y(n_1157)
);

NAND3xp33_ASAP7_75t_L g1158 ( 
.A(n_1144),
.B(n_46),
.C(n_47),
.Y(n_1158)
);

AOI311xp33_ASAP7_75t_L g1159 ( 
.A1(n_1125),
.A2(n_49),
.A3(n_52),
.B(n_53),
.C(n_54),
.Y(n_1159)
);

NOR2x1_ASAP7_75t_L g1160 ( 
.A(n_1135),
.B(n_52),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1141),
.Y(n_1161)
);

AOI211xp5_ASAP7_75t_L g1162 ( 
.A1(n_1137),
.A2(n_54),
.B(n_55),
.C(n_56),
.Y(n_1162)
);

INVx2_ASAP7_75t_SL g1163 ( 
.A(n_1139),
.Y(n_1163)
);

AOI221x1_ASAP7_75t_L g1164 ( 
.A1(n_1140),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.C(n_61),
.Y(n_1164)
);

NOR2x1_ASAP7_75t_L g1165 ( 
.A(n_1143),
.B(n_57),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1133),
.B(n_1138),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1128),
.A2(n_999),
.B(n_967),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1125),
.A2(n_993),
.B(n_932),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1147),
.A2(n_917),
.B(n_937),
.C(n_62),
.Y(n_1169)
);

AOI221xp5_ASAP7_75t_L g1170 ( 
.A1(n_1126),
.A2(n_58),
.B1(n_61),
.B2(n_63),
.C(n_941),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1142),
.A2(n_977),
.B(n_917),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1148),
.B(n_927),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1149),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1155),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1163),
.Y(n_1175)
);

NOR2x1_ASAP7_75t_L g1176 ( 
.A(n_1158),
.B(n_937),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1160),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1153),
.B(n_991),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1165),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_1156),
.B(n_879),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1161),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1154),
.B(n_879),
.Y(n_1182)
);

NAND4xp25_ASAP7_75t_L g1183 ( 
.A(n_1170),
.B(n_991),
.C(n_939),
.D(n_998),
.Y(n_1183)
);

XOR2x1_ASAP7_75t_L g1184 ( 
.A(n_1159),
.B(n_65),
.Y(n_1184)
);

NAND4xp75_ASAP7_75t_L g1185 ( 
.A(n_1164),
.B(n_998),
.C(n_994),
.D(n_936),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1169),
.B(n_936),
.Y(n_1186)
);

NAND4xp75_ASAP7_75t_L g1187 ( 
.A(n_1151),
.B(n_994),
.C(n_936),
.D(n_939),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1166),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1162),
.Y(n_1189)
);

XNOR2xp5_ASAP7_75t_L g1190 ( 
.A(n_1150),
.B(n_66),
.Y(n_1190)
);

NAND5xp2_ASAP7_75t_L g1191 ( 
.A(n_1168),
.B(n_984),
.C(n_1010),
.D(n_75),
.E(n_76),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1171),
.B(n_997),
.Y(n_1192)
);

XNOR2xp5_ASAP7_75t_L g1193 ( 
.A(n_1157),
.B(n_68),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1173),
.B(n_1152),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1174),
.B(n_1167),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1175),
.B(n_997),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1188),
.B(n_922),
.Y(n_1197)
);

NOR3xp33_ASAP7_75t_L g1198 ( 
.A(n_1172),
.B(n_1179),
.C(n_1189),
.Y(n_1198)
);

NAND4xp75_ASAP7_75t_L g1199 ( 
.A(n_1181),
.B(n_1176),
.C(n_1177),
.D(n_1180),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1178),
.B(n_923),
.Y(n_1200)
);

NAND3x1_ASAP7_75t_SL g1201 ( 
.A(n_1184),
.B(n_74),
.C(n_77),
.Y(n_1201)
);

NAND4xp25_ASAP7_75t_L g1202 ( 
.A(n_1178),
.B(n_939),
.C(n_923),
.D(n_924),
.Y(n_1202)
);

NOR4xp75_ASAP7_75t_L g1203 ( 
.A(n_1185),
.B(n_79),
.C(n_85),
.D(n_87),
.Y(n_1203)
);

NAND4xp75_ASAP7_75t_L g1204 ( 
.A(n_1182),
.B(n_939),
.C(n_89),
.D(n_90),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1193),
.A2(n_927),
.B1(n_932),
.B2(n_923),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1192),
.B(n_927),
.Y(n_1206)
);

AOI31xp33_ASAP7_75t_L g1207 ( 
.A1(n_1190),
.A2(n_88),
.A3(n_91),
.B(n_92),
.Y(n_1207)
);

OAI322xp33_ASAP7_75t_L g1208 ( 
.A1(n_1186),
.A2(n_927),
.A3(n_914),
.B1(n_924),
.B2(n_919),
.C1(n_913),
.C2(n_915),
.Y(n_1208)
);

XNOR2x1_ASAP7_75t_L g1209 ( 
.A(n_1199),
.B(n_1186),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1195),
.B(n_1191),
.Y(n_1210)
);

XNOR2xp5_ASAP7_75t_L g1211 ( 
.A(n_1201),
.B(n_1183),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_SL g1212 ( 
.A1(n_1207),
.A2(n_1191),
.B(n_1183),
.Y(n_1212)
);

AND3x1_ASAP7_75t_L g1213 ( 
.A(n_1198),
.B(n_1187),
.C(n_95),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1194),
.A2(n_927),
.B1(n_932),
.B2(n_924),
.Y(n_1214)
);

NAND4xp75_ASAP7_75t_L g1215 ( 
.A(n_1197),
.B(n_93),
.C(n_96),
.D(n_97),
.Y(n_1215)
);

INVx1_ASAP7_75t_SL g1216 ( 
.A(n_1199),
.Y(n_1216)
);

AOI211xp5_ASAP7_75t_L g1217 ( 
.A1(n_1196),
.A2(n_927),
.B(n_99),
.C(n_100),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1200),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_R g1219 ( 
.A(n_1204),
.B(n_98),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1203),
.Y(n_1220)
);

O2A1O1Ixp5_ASAP7_75t_L g1221 ( 
.A1(n_1206),
.A2(n_101),
.B(n_103),
.C(n_108),
.Y(n_1221)
);

NAND3xp33_ASAP7_75t_L g1222 ( 
.A(n_1202),
.B(n_927),
.C(n_932),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1205),
.Y(n_1223)
);

AO22x2_ASAP7_75t_L g1224 ( 
.A1(n_1209),
.A2(n_1208),
.B1(n_113),
.B2(n_115),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_SL g1225 ( 
.A1(n_1216),
.A2(n_927),
.B1(n_932),
.B2(n_924),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1220),
.A2(n_932),
.B1(n_913),
.B2(n_924),
.Y(n_1226)
);

OAI22x1_ASAP7_75t_L g1227 ( 
.A1(n_1211),
.A2(n_914),
.B1(n_116),
.B2(n_123),
.Y(n_1227)
);

OA22x2_ASAP7_75t_L g1228 ( 
.A1(n_1212),
.A2(n_932),
.B1(n_914),
.B2(n_918),
.Y(n_1228)
);

OAI22x1_ASAP7_75t_L g1229 ( 
.A1(n_1210),
.A2(n_110),
.B1(n_124),
.B2(n_129),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1214),
.A2(n_932),
.B1(n_915),
.B2(n_987),
.Y(n_1230)
);

INVx1_ASAP7_75t_SL g1231 ( 
.A(n_1219),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1218),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1213),
.A2(n_915),
.B1(n_987),
.B2(n_139),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1229),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1232),
.A2(n_1223),
.B1(n_1222),
.B2(n_1217),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1224),
.Y(n_1236)
);

AOI22x1_ASAP7_75t_L g1237 ( 
.A1(n_1227),
.A2(n_1231),
.B1(n_1224),
.B2(n_1221),
.Y(n_1237)
);

AO22x1_ASAP7_75t_L g1238 ( 
.A1(n_1233),
.A2(n_1221),
.B1(n_1215),
.B2(n_140),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1226),
.B(n_134),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1236),
.A2(n_1225),
.B1(n_1228),
.B2(n_1230),
.Y(n_1240)
);

OAI22x1_ASAP7_75t_SL g1241 ( 
.A1(n_1234),
.A2(n_136),
.B1(n_143),
.B2(n_144),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1235),
.A2(n_974),
.B1(n_915),
.B2(n_938),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1237),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1243),
.A2(n_1239),
.B(n_1238),
.Y(n_1244)
);

AOI221xp5_ASAP7_75t_L g1245 ( 
.A1(n_1244),
.A2(n_1240),
.B1(n_1241),
.B2(n_1242),
.C(n_157),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1245),
.B(n_150),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1246),
.Y(n_1247)
);

AOI221xp5_ASAP7_75t_L g1248 ( 
.A1(n_1247),
.A2(n_152),
.B1(n_155),
.B2(n_160),
.C(n_161),
.Y(n_1248)
);

AOI211xp5_ASAP7_75t_L g1249 ( 
.A1(n_1248),
.A2(n_162),
.B(n_164),
.C(n_167),
.Y(n_1249)
);


endmodule