module real_jpeg_14306_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_213;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_3),
.A2(n_33),
.B1(n_55),
.B2(n_57),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_4),
.A2(n_41),
.B1(n_42),
.B2(n_74),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_4),
.A2(n_55),
.B1(n_57),
.B2(n_74),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_74),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_50),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_6),
.A2(n_50),
.B1(n_55),
.B2(n_57),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_50),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_7),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_71),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_7),
.A2(n_55),
.B1(n_57),
.B2(n_71),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_71),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_10),
.A2(n_35),
.B1(n_55),
.B2(n_57),
.Y(n_95)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_12),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_12),
.A2(n_55),
.B1(n_57),
.B2(n_84),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_84),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_13),
.A2(n_37),
.B(n_38),
.C(n_43),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_13),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_13),
.B(n_115),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_13),
.A2(n_40),
.B1(n_55),
.B2(n_57),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_13),
.A2(n_100),
.B1(n_104),
.B2(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_13),
.B(n_61),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_14),
.A2(n_41),
.B1(n_42),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_14),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_63),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_14),
.A2(n_55),
.B1(n_57),
.B2(n_63),
.Y(n_122)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_131),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_116),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_19),
.B(n_116),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_75),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_47),
.C(n_64),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_21),
.A2(n_22),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_23),
.A2(n_24),
.B1(n_36),
.B2(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_25),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_25),
.A2(n_80),
.B(n_103),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_25),
.A2(n_30),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_26),
.A2(n_27),
.B1(n_90),
.B2(n_91),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_26),
.B(n_40),
.C(n_91),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_26),
.B(n_185),
.Y(n_184)
);

CKINVDCx6p67_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_30),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_32),
.A2(n_81),
.B(n_104),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_34),
.Y(n_101)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_36),
.Y(n_213)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_37),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B(n_41),
.Y(n_38)
);

HAxp5_ASAP7_75t_SL g142 ( 
.A(n_40),
.B(n_42),
.CON(n_142),
.SN(n_142)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_40),
.B(n_104),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_40),
.B(n_93),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_42),
.B1(n_54),
.B2(n_58),
.Y(n_59)
);

NOR3xp33_ASAP7_75t_L g143 ( 
.A(n_41),
.B(n_55),
.C(n_58),
.Y(n_143)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_47),
.B(n_64),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B(n_60),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_49),
.A2(n_52),
.B1(n_61),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_51),
.A2(n_53),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_52),
.A2(n_62),
.B(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_52),
.A2(n_61),
.B1(n_142),
.B2(n_153),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_53),
.B(n_112),
.Y(n_111)
);

OA22x2_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_54),
.A2(n_57),
.B(n_141),
.C(n_143),
.Y(n_140)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_55),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_57),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_57),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_68),
.B1(n_69),
.B2(n_72),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_66),
.A2(n_73),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_66),
.A2(n_70),
.B1(n_115),
.B2(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_97),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_85),
.B2(n_96),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_79),
.A2(n_100),
.B(n_181),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_104),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_85),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_88),
.B1(n_94),
.B2(n_95),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_93),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_88),
.A2(n_94),
.B1(n_148),
.B2(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_88),
.A2(n_94),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_88),
.A2(n_94),
.B1(n_164),
.B2(n_174),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_94),
.B(n_122),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_109),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_105),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_105),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B(n_102),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_100),
.A2(n_104),
.B1(n_179),
.B2(n_187),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.C(n_128),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_117),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_120),
.B(n_128),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.C(n_126),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_121),
.B(n_124),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_126),
.B(n_216),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_223),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_219),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_209),
.B(n_218),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_165),
.B(n_208),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_160),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_137),
.B(n_160),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_150),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_145),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_139),
.B(n_145),
.C(n_150),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_140),
.B(n_144),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B(n_149),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_155),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_151),
.B(n_156),
.C(n_159),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.C(n_163),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_163),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_203),
.B(n_207),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_193),
.B(n_202),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_182),
.B(n_192),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_177),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_177),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_172),
.B1(n_175),
.B2(n_176),
.Y(n_169)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_175),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_188),
.B(n_191),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_190),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_195),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_198),
.C(n_201),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_200),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_206),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_217),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_217),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_214),
.C(n_215),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_222),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);


endmodule