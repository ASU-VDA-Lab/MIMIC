module fake_jpeg_589_n_411 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_411);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_411;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_56),
.Y(n_126)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_58),
.Y(n_157)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_61),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_26),
.B(n_7),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_62),
.B(n_65),
.Y(n_139)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_63),
.Y(n_150)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_26),
.B(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_68),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_34),
.Y(n_113)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_71),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_30),
.B(n_7),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_72),
.B(n_89),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_74),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_76),
.Y(n_162)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_29),
.Y(n_77)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_30),
.B(n_10),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_91),
.Y(n_114)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_80),
.Y(n_143)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_81),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_29),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_84),
.A2(n_2),
.B(n_3),
.Y(n_160)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_86),
.Y(n_163)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_43),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_10),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_45),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_54),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_35),
.B(n_29),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_99),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_31),
.B(n_11),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

BUFx2_ASAP7_75t_SL g175 ( 
.A(n_97),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_100),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_41),
.B(n_1),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_102),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_37),
.B(n_15),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_111),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_105),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_18),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_27),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_106),
.B(n_107),
.Y(n_169)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_21),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_23),
.Y(n_138)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_109),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_34),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_110),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_37),
.B(n_15),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_76),
.A2(n_38),
.B1(n_47),
.B2(n_18),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_112),
.A2(n_116),
.B1(n_119),
.B2(n_121),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_113),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_38),
.B1(n_47),
.B2(n_34),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_67),
.A2(n_21),
.B1(n_23),
.B2(n_44),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_86),
.A2(n_33),
.B1(n_94),
.B2(n_96),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_62),
.A2(n_72),
.B1(n_89),
.B2(n_51),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_122),
.A2(n_140),
.B1(n_146),
.B2(n_167),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_53),
.B1(n_51),
.B2(n_50),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_124),
.A2(n_136),
.B1(n_116),
.B2(n_150),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_95),
.A2(n_53),
.B1(n_50),
.B2(n_42),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_114),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_103),
.A2(n_42),
.B1(n_22),
.B2(n_36),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_22),
.B(n_36),
.Y(n_141)
);

BUFx24_ASAP7_75t_SL g189 ( 
.A(n_141),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_106),
.A2(n_19),
.B1(n_25),
.B2(n_44),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_65),
.A2(n_19),
.B1(n_25),
.B2(n_44),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_160),
.B(n_171),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_92),
.B(n_1),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_153),
.B(n_164),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_93),
.B(n_44),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_155),
.B(n_157),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_77),
.B(n_2),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_174),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_110),
.B(n_3),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_68),
.A2(n_5),
.B1(n_32),
.B2(n_90),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_84),
.A2(n_5),
.B1(n_71),
.B2(n_73),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_80),
.B(n_5),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_118),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_177),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_5),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_134),
.A2(n_175),
.B1(n_169),
.B2(n_165),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_180),
.A2(n_203),
.B1(n_192),
.B2(n_210),
.Y(n_268)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_181),
.Y(n_267)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_182),
.B(n_195),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_127),
.B(n_155),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_183),
.B(n_227),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_140),
.A2(n_122),
.B1(n_123),
.B2(n_146),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_184),
.A2(n_207),
.B1(n_190),
.B2(n_226),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_119),
.A2(n_132),
.B1(n_156),
.B2(n_168),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_185),
.A2(n_193),
.B1(n_219),
.B2(n_209),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_187),
.B(n_188),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_123),
.B(n_115),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_128),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_191),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_192),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_132),
.A2(n_156),
.B1(n_168),
.B2(n_120),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_147),
.Y(n_194)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_144),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_134),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_196),
.Y(n_233)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_198),
.Y(n_249)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_199),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_115),
.B(n_135),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_201),
.Y(n_236)
);

AOI32xp33_ASAP7_75t_L g201 ( 
.A1(n_125),
.A2(n_165),
.A3(n_129),
.B1(n_154),
.B2(n_163),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_202),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_169),
.A2(n_149),
.B1(n_151),
.B2(n_133),
.Y(n_203)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_143),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g257 ( 
.A(n_205),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_208),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_131),
.B(n_151),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_207),
.Y(n_230)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_150),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_152),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_209),
.B(n_213),
.Y(n_263)
);

INVx13_ASAP7_75t_L g210 ( 
.A(n_143),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_210),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_131),
.B(n_149),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_212),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_214),
.B(n_215),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_145),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_133),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_216),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_226),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_161),
.B(n_166),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_229),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_161),
.A2(n_166),
.B1(n_130),
.B2(n_170),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_126),
.B(n_157),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_220),
.B(n_221),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_126),
.B(n_143),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_137),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_222),
.Y(n_245)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_223),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_172),
.B(n_129),
.Y(n_224)
);

HAxp5_ASAP7_75t_SL g231 ( 
.A(n_224),
.B(n_225),
.CON(n_231),
.SN(n_231)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_172),
.B(n_129),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_130),
.B(n_137),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_112),
.B(n_121),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_139),
.B(n_158),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_228),
.B(n_211),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_127),
.B(n_141),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_229),
.A2(n_178),
.B(n_189),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_234),
.A2(n_239),
.B(n_259),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_204),
.A2(n_176),
.B(n_213),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_241),
.B(n_258),
.Y(n_300)
);

A2O1A1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_187),
.A2(n_176),
.B(n_183),
.C(n_186),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_L g277 ( 
.A1(n_242),
.A2(n_244),
.B(n_252),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_187),
.A2(n_218),
.B1(n_196),
.B2(n_212),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_246),
.A2(n_253),
.B1(n_230),
.B2(n_233),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_251),
.B(n_259),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_212),
.A2(n_207),
.B1(n_202),
.B2(n_199),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_197),
.A2(n_222),
.B1(n_181),
.B2(n_194),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_256),
.A2(n_266),
.B1(n_248),
.B2(n_245),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_177),
.B(n_226),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_177),
.B(n_215),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_248),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_191),
.A2(n_223),
.B1(n_198),
.B2(n_206),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_268),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_270),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_272),
.B(n_283),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_235),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_273),
.B(n_274),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_252),
.B(n_235),
.Y(n_274)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_275),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_239),
.A2(n_263),
.B1(n_244),
.B2(n_258),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_276),
.A2(n_281),
.B1(n_282),
.B2(n_297),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_277),
.B(n_299),
.Y(n_314)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_278),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_242),
.B(n_246),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_279),
.B(n_284),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_263),
.A2(n_236),
.B1(n_255),
.B2(n_261),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_236),
.A2(n_255),
.B1(n_261),
.B2(n_230),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_270),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_255),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_285),
.B(n_286),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_264),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_254),
.Y(n_287)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_287),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_247),
.B(n_232),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_288),
.B(n_289),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_242),
.B(n_233),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_232),
.B(n_262),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_290),
.B(n_298),
.Y(n_324)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_254),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_291),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_292),
.A2(n_296),
.B(n_260),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_294),
.B(n_303),
.Y(n_327)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_243),
.Y(n_295)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_295),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_253),
.A2(n_241),
.B1(n_234),
.B2(n_231),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_249),
.A2(n_245),
.B1(n_250),
.B2(n_243),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_265),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_268),
.B(n_240),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_238),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_301),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_265),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_302),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_262),
.B(n_238),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_306),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_300),
.A2(n_249),
.B1(n_260),
.B2(n_266),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_310),
.A2(n_313),
.B1(n_275),
.B2(n_297),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_279),
.B(n_240),
.C(n_257),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_316),
.C(n_272),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_300),
.A2(n_271),
.B1(n_250),
.B2(n_267),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_282),
.B(n_237),
.C(n_267),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_290),
.Y(n_320)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_320),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_274),
.B(n_237),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_322),
.B(n_284),
.Y(n_335)
);

AOI322xp5_ASAP7_75t_L g323 ( 
.A1(n_289),
.A2(n_256),
.A3(n_267),
.B1(n_285),
.B2(n_273),
.C1(n_286),
.C2(n_300),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_323),
.B(n_278),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_325),
.B(n_280),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_328),
.B(n_332),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_329),
.A2(n_345),
.B1(n_347),
.B2(n_309),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_305),
.A2(n_296),
.B1(n_294),
.B2(n_276),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_330),
.A2(n_304),
.B1(n_307),
.B2(n_326),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_301),
.Y(n_331)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_331),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_326),
.B(n_288),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_281),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_338),
.C(n_341),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_335),
.B(n_336),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_312),
.A2(n_292),
.B1(n_280),
.B2(n_293),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_337),
.B(n_339),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_292),
.C(n_299),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_303),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_315),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_340),
.B(n_344),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_314),
.B(n_299),
.C(n_295),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_283),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_342),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_319),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_312),
.A2(n_304),
.B1(n_310),
.B2(n_320),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_322),
.B(n_287),
.C(n_291),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_346),
.B(n_316),
.C(n_308),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_343),
.A2(n_306),
.B(n_327),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_357),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_343),
.A2(n_327),
.B(n_331),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_350),
.B(n_362),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_352),
.A2(n_353),
.B1(n_354),
.B2(n_317),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_330),
.A2(n_307),
.B1(n_311),
.B2(n_324),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_339),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_358),
.B(n_359),
.C(n_346),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_336),
.B(n_308),
.C(n_315),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_338),
.A2(n_333),
.B(n_341),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_364),
.B(n_365),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_351),
.B(n_335),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_363),
.Y(n_366)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_366),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_351),
.B(n_332),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_369),
.B(n_371),
.Y(n_384)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_363),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_370),
.B(n_373),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_359),
.B(n_334),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_334),
.C(n_344),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_372),
.B(n_376),
.Y(n_381)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_355),
.Y(n_373)
);

OAI22x1_ASAP7_75t_L g374 ( 
.A1(n_360),
.A2(n_313),
.B1(n_340),
.B2(n_317),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_374),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_375),
.B(n_353),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_348),
.B(n_318),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_368),
.A2(n_352),
.B1(n_361),
.B2(n_360),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_378),
.Y(n_394)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_380),
.Y(n_389)
);

FAx1_ASAP7_75t_SL g382 ( 
.A(n_369),
.B(n_349),
.CI(n_357),
.CON(n_382),
.SN(n_382)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_382),
.B(n_386),
.Y(n_391)
);

FAx1_ASAP7_75t_SL g386 ( 
.A(n_372),
.B(n_362),
.CI(n_350),
.CON(n_386),
.SN(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_356),
.Y(n_387)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_387),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_377),
.B(n_356),
.Y(n_388)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_388),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_383),
.B(n_364),
.C(n_376),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_390),
.B(n_393),
.C(n_384),
.Y(n_399)
);

INVxp33_ASAP7_75t_L g392 ( 
.A(n_379),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_392),
.B(n_355),
.Y(n_395)
);

XNOR2x1_ASAP7_75t_L g393 ( 
.A(n_384),
.B(n_354),
.Y(n_393)
);

AO21x2_ASAP7_75t_L g401 ( 
.A1(n_395),
.A2(n_385),
.B(n_389),
.Y(n_401)
);

AOI31xp67_ASAP7_75t_SL g398 ( 
.A1(n_392),
.A2(n_382),
.A3(n_358),
.B(n_386),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_398),
.B(n_400),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_399),
.B(n_391),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_390),
.B(n_383),
.C(n_371),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_401),
.B(n_403),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_396),
.B(n_394),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_404),
.B(n_393),
.Y(n_407)
);

NAND3xp33_ASAP7_75t_L g406 ( 
.A(n_402),
.B(n_397),
.C(n_367),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_406),
.B(n_407),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_405),
.B(n_395),
.C(n_401),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_409),
.A2(n_386),
.B(n_382),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_410),
.B(n_408),
.Y(n_411)
);


endmodule