module real_jpeg_4731_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g84 ( 
.A(n_0),
.Y(n_84)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_1),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_1),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_1),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_2),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_2),
.A2(n_44),
.B1(n_136),
.B2(n_140),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_2),
.A2(n_44),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_2),
.A2(n_44),
.B1(n_203),
.B2(n_205),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_3),
.A2(n_33),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_3),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_3),
.A2(n_132),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_3),
.A2(n_132),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_3),
.A2(n_132),
.B1(n_165),
.B2(n_270),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_4),
.A2(n_26),
.B1(n_103),
.B2(n_107),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_4),
.A2(n_26),
.B1(n_171),
.B2(n_174),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_4),
.A2(n_26),
.B1(n_211),
.B2(n_213),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_4),
.B(n_31),
.Y(n_278)
);

O2A1O1Ixp33_ASAP7_75t_L g335 ( 
.A1(n_4),
.A2(n_336),
.B(n_338),
.C(n_344),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_4),
.B(n_86),
.C(n_165),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_4),
.B(n_142),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_4),
.B(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_4),
.B(n_90),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_5),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_5),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_5),
.A2(n_219),
.B1(n_254),
.B2(n_257),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_5),
.A2(n_219),
.B1(n_351),
.B2(n_352),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_5),
.A2(n_219),
.B1(n_372),
.B2(n_374),
.Y(n_371)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_6),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_7),
.Y(n_167)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_7),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_7),
.Y(n_389)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_8),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_9),
.A2(n_15),
.B1(n_18),
.B2(n_20),
.Y(n_14)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_11),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_11),
.Y(n_231)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_13),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_13),
.Y(n_92)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_13),
.Y(n_99)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_446),
.Y(n_20)
);

OAI221xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_59),
.B1(n_63),
.B2(n_441),
.C(n_444),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_22),
.B(n_445),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_22),
.B(n_59),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_23),
.B(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_24),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_25),
.B(n_48),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B(n_28),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_26),
.B(n_29),
.Y(n_28)
);

OAI21xp33_ASAP7_75t_L g338 ( 
.A1(n_26),
.A2(n_339),
.B(n_341),
.Y(n_338)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_27),
.Y(n_228)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_28),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_29),
.Y(n_220)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_31),
.B(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_31),
.B(n_217),
.Y(n_248)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_36),
.B2(n_38),
.Y(n_31)
);

NAND2xp33_ASAP7_75t_SL g267 ( 
.A(n_32),
.B(n_118),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_33),
.A2(n_113),
.B1(n_116),
.B2(n_117),
.Y(n_112)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_35),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_35),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g212 ( 
.A(n_35),
.Y(n_212)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_41),
.A2(n_61),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_41),
.B(n_248),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_48),
.Y(n_41)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_48),
.B(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_55),
.B2(n_57),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_59),
.A2(n_159),
.B(n_186),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_59),
.A2(n_161),
.B1(n_186),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_59),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B(n_62),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_60),
.A2(n_72),
.B(n_227),
.Y(n_437)
);

A2O1A1O1Ixp25_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_241),
.B(n_430),
.C(n_433),
.D(n_440),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_221),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_187),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_66),
.B(n_187),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_158),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_143),
.B2(n_144),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_69),
.B(n_143),
.C(n_158),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_70),
.A2(n_71),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_71),
.B(n_76),
.C(n_109),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_71),
.B(n_224),
.C(n_239),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_72),
.B(n_216),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_73),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_108),
.B2(n_109),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_76),
.A2(n_77),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_76),
.A2(n_77),
.B1(n_250),
.B2(n_258),
.Y(n_249)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_77),
.B(n_247),
.C(n_250),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_77),
.B(n_235),
.C(n_238),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_100),
.B(n_101),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_78),
.A2(n_179),
.B(n_185),
.Y(n_178)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_79),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_79),
.B(n_102),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_79),
.B(n_350),
.Y(n_349)
);

NOR2x1_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_90),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_83),
.Y(n_351)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_84),
.Y(n_343)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_88),
.Y(n_181)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_90),
.B(n_149),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_90),
.B(n_350),
.Y(n_366)
);

AO22x1_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_93),
.B1(n_96),
.B2(n_98),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_93),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_94),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_95),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_97),
.Y(n_375)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_100),
.B(n_101),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_100),
.A2(n_148),
.B(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g184 ( 
.A(n_107),
.Y(n_184)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_129),
.B(n_133),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_110),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_110),
.B(n_253),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_110),
.A2(n_142),
.B(n_210),
.Y(n_306)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_111),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_119),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_114),
.Y(n_337)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_115),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_119),
.B(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_122),
.B1(n_123),
.B2(n_126),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_125),
.Y(n_354)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_142),
.B(n_156),
.Y(n_155)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_134),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_134),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_142),
.Y(n_134)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_138),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_141),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_142),
.B(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_144),
.A2(n_145),
.B(n_155),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_155),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_146),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_148),
.B(n_366),
.Y(n_410)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_156),
.B(n_236),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_156),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_160),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_178),
.Y(n_160)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_161),
.A2(n_178),
.B1(n_186),
.B2(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_161),
.B(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_161),
.A2(n_186),
.B1(n_335),
.B2(n_413),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_168),
.B(n_170),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_162),
.B(n_170),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_162),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_162),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_174),
.Y(n_270)
);

INVx4_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_178),
.Y(n_318)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g290 ( 
.A(n_185),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_185),
.B(n_349),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_192),
.C(n_194),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_188),
.A2(n_192),
.B1(n_193),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_188),
.Y(n_322)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_194),
.B(n_321),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_208),
.C(n_215),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_195),
.A2(n_196),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_207),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_197),
.B(n_207),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_198),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_200),
.B(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_201),
.A2(n_269),
.B(n_271),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_202),
.B(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx8_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g395 ( 
.A(n_206),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_208),
.B(n_215),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_209),
.B(n_252),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g237 ( 
.A(n_210),
.Y(n_237)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_211),
.Y(n_257)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_221),
.A2(n_431),
.B(n_432),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_240),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_222),
.B(n_240),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_239),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_232),
.B1(n_233),
.B2(n_238),
.Y(n_225)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_226),
.Y(n_238)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

AOI32xp33_ASAP7_75t_L g261 ( 
.A1(n_231),
.A2(n_262),
.A3(n_263),
.B1(n_266),
.B2(n_267),
.Y(n_261)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_236),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_422),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_311),
.C(n_325),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_298),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_284),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_245),
.B(n_284),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_259),
.C(n_274),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_246),
.B(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_255),
.Y(n_262)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_259),
.A2(n_260),
.B1(n_274),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_268),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_261),
.B(n_268),
.Y(n_293)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_269),
.A2(n_281),
.B(n_289),
.Y(n_288)
);

INVx8_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_273),
.Y(n_283)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_273),
.Y(n_397)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_274),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.C(n_279),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_275),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_297),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_279),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_280),
.B(n_387),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_281),
.B(n_370),
.Y(n_400)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_292),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_287),
.C(n_292),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_290),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_291),
.B(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_295),
.C(n_296),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_298),
.A2(n_425),
.B(n_426),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_310),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_299),
.B(n_310),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_302),
.C(n_303),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_307),
.C(n_308),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_306),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_306),
.A2(n_308),
.B1(n_436),
.B2(n_437),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_306),
.B(n_437),
.C(n_438),
.Y(n_443)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_307),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_323),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_312),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_320),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_313),
.B(n_324),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_313),
.B(n_324),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_313),
.B(n_320),
.Y(n_429)
);

FAx1_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_317),
.CI(n_319),
.CON(n_313),
.SN(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_323),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_355),
.B(n_421),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_330),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_327),
.B(n_330),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_334),
.C(n_346),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_331),
.B(n_417),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_334),
.A2(n_346),
.B1(n_347),
.B2(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_334),
.Y(n_418)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_335),
.Y(n_413)
);

INVx8_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx6_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_343),
.Y(n_363)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx6_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_415),
.B(n_420),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_357),
.A2(n_405),
.B(n_414),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_381),
.B(n_404),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_367),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_359),
.B(n_367),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_365),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_360),
.A2(n_361),
.B1(n_365),
.B2(n_384),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_364),
.Y(n_361)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_365),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_376),
.Y(n_367)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_368),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_388),
.Y(n_387)
);

INVx6_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_377),
.A2(n_378),
.B1(n_379),
.B2(n_380),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_377),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_378),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_378),
.B(n_379),
.C(n_407),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_382),
.A2(n_390),
.B(n_403),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_385),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_383),
.B(n_385),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_391),
.A2(n_399),
.B(n_402),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_398),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_396),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_394),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_400),
.B(n_401),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_408),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_406),
.B(n_408),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_412),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_410),
.B(n_411),
.C(n_412),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_416),
.B(n_419),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_416),
.B(n_419),
.Y(n_420)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g422 ( 
.A1(n_423),
.A2(n_424),
.B(n_427),
.C(n_428),
.D(n_429),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_439),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_434),
.B(n_439),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_438),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_443),
.Y(n_445)
);


endmodule