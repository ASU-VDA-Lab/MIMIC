module real_jpeg_27007_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_341, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_341;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_0),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_0),
.A2(n_27),
.B1(n_31),
.B2(n_46),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_0),
.A2(n_46),
.B1(n_59),
.B2(n_62),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_25),
.B1(n_53),
.B2(n_54),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_1),
.A2(n_25),
.B1(n_27),
.B2(n_31),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_1),
.A2(n_25),
.B1(n_59),
.B2(n_62),
.Y(n_99)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_2),
.Y(n_95)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_2),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_3),
.A2(n_27),
.B1(n_31),
.B2(n_37),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_3),
.A2(n_37),
.B1(n_59),
.B2(n_62),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_3),
.A2(n_37),
.B1(n_53),
.B2(n_54),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_5),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_5),
.A2(n_48),
.B1(n_59),
.B2(n_62),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_5),
.A2(n_27),
.B1(n_31),
.B2(n_48),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_8),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_8),
.A2(n_27),
.B1(n_31),
.B2(n_136),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_8),
.A2(n_53),
.B1(n_54),
.B2(n_136),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_8),
.A2(n_59),
.B1(n_62),
.B2(n_136),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_9),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_9),
.A2(n_27),
.B1(n_31),
.B2(n_110),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_9),
.A2(n_53),
.B1(n_54),
.B2(n_110),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_9),
.A2(n_59),
.B1(n_62),
.B2(n_110),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_10),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_10),
.A2(n_27),
.B1(n_31),
.B2(n_171),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_10),
.A2(n_53),
.B1(n_54),
.B2(n_171),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_10),
.A2(n_59),
.B1(n_62),
.B2(n_171),
.Y(n_256)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_12),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_12),
.B(n_26),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_12),
.B(n_31),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g212 ( 
.A1(n_12),
.A2(n_31),
.B(n_208),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_12),
.A2(n_53),
.B1(n_54),
.B2(n_169),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_12),
.A2(n_56),
.B(n_59),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_12),
.B(n_78),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_12),
.A2(n_114),
.B1(n_115),
.B2(n_256),
.Y(n_258)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

INVx11_ASAP7_75t_SL g61 ( 
.A(n_15),
.Y(n_61)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_339),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_83),
.B(n_337),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_38),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_20),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_32),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_21),
.A2(n_44),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_22),
.A2(n_33),
.B(n_82),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_22),
.A2(n_26),
.B(n_33),
.Y(n_339)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_26),
.B(n_29),
.C(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_29),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g168 ( 
.A(n_23),
.B(n_169),
.CON(n_168),
.SN(n_168)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_26),
.A2(n_33),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_27),
.A2(n_31),
.B1(n_68),
.B2(n_69),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_27),
.A2(n_34),
.B1(n_168),
.B2(n_182),
.Y(n_181)
);

AOI32xp33_ASAP7_75t_L g206 ( 
.A1(n_27),
.A2(n_53),
.A3(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_206)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_29),
.B(n_31),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_32),
.A2(n_45),
.B(n_49),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_33),
.A2(n_81),
.B(n_82),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_36),
.B(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_39),
.B(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_75),
.C(n_80),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_40),
.A2(n_41),
.B1(n_333),
.B2(n_335),
.Y(n_332)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_50),
.C(n_65),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_42),
.A2(n_43),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_44),
.A2(n_49),
.B1(n_109),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_44),
.A2(n_49),
.B1(n_135),
.B2(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_47),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_50),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_50),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_50),
.A2(n_65),
.B1(n_305),
.B2(n_319),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_58),
.B(n_63),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_51),
.A2(n_58),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_51),
.A2(n_102),
.B(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_51),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_51),
.A2(n_63),
.B(n_118),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_51),
.A2(n_58),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_51),
.A2(n_142),
.B(n_216),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_51),
.A2(n_58),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_51),
.A2(n_58),
.B1(n_215),
.B2(n_233),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_58),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_54),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g209 ( 
.A(n_54),
.B(n_68),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_54),
.A2(n_57),
.B(n_169),
.C(n_235),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_62),
.Y(n_58)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_58),
.A2(n_101),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_58),
.B(n_169),
.Y(n_254)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

BUFx4f_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_62),
.B(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_64),
.B(n_120),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_65),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_71),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_66),
.A2(n_77),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_67),
.B(n_72),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_67),
.A2(n_73),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_67),
.A2(n_73),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_67),
.A2(n_73),
.B1(n_165),
.B2(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_67),
.A2(n_73),
.B1(n_193),
.B2(n_212),
.Y(n_211)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_68),
.Y(n_207)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_71),
.A2(n_78),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_75),
.A2(n_76),
.B1(n_80),
.B2(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B(n_79),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_77),
.A2(n_79),
.B(n_132),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_77),
.A2(n_132),
.B(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_80),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_330),
.B(n_336),
.Y(n_83)
);

OAI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_300),
.A3(n_322),
.B1(n_328),
.B2(n_329),
.C(n_341),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_154),
.B(n_299),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_137),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_87),
.B(n_137),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_111),
.C(n_122),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_88),
.A2(n_89),
.B1(n_111),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_103),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_90),
.B(n_105),
.C(n_107),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_100),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_91),
.B(n_100),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_98),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_92),
.A2(n_184),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_93),
.A2(n_99),
.B(n_127),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_93),
.A2(n_94),
.B1(n_247),
.B2(n_249),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_99),
.Y(n_98)
);

INVx11_ASAP7_75t_L g197 ( 
.A(n_94),
.Y(n_197)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_95),
.A2(n_114),
.B1(n_125),
.B2(n_184),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_115),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_98),
.A2(n_114),
.B(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_106),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_111),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_117),
.B2(n_121),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_112),
.A2(n_113),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_117),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_113),
.A2(n_148),
.B(n_151),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B(n_116),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_125),
.B(n_126),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_114),
.A2(n_197),
.B1(n_248),
.B2(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_115),
.B(n_169),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_117),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_119),
.B(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_122),
.B(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_131),
.C(n_133),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_123),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_128),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_131),
.A2(n_133),
.B1(n_134),
.B2(n_289),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_131),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_152),
.B2(n_153),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_147),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_140),
.B(n_147),
.C(n_153),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_143),
.B(n_146),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_143),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_145),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_146),
.B(n_302),
.C(n_312),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_146),
.A2(n_302),
.B1(n_303),
.B2(n_327),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_146),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_152),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_293),
.B(n_298),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_198),
.B(n_279),
.C(n_292),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_185),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_157),
.B(n_185),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_172),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_159),
.B(n_160),
.C(n_172),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.C(n_167),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_167),
.B(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_170),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_180),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_174),
.B(n_178),
.C(n_180),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_183),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.C(n_191),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_186),
.A2(n_187),
.B1(n_274),
.B2(n_276),
.Y(n_273)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_191),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.C(n_196),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_196),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_278),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_271),
.B(n_277),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_226),
.B(n_270),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_217),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_202),
.B(n_217),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_210),
.C(n_213),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_203),
.A2(n_204),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_206),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_223),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_218),
.B(n_224),
.C(n_225),
.Y(n_272)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_264),
.B(n_269),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_244),
.B(n_263),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_236),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_229),
.B(n_236),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_234),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_230),
.A2(n_231),
.B1(n_234),
.B2(n_251),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_234),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_242),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_241),
.C(n_242),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_243),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_252),
.B(n_262),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_250),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_246),
.B(n_250),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_257),
.B(n_261),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_254),
.B(n_255),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_272),
.B(n_273),
.Y(n_277)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_274),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_280),
.B(n_281),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_290),
.B2(n_291),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_287),
.C(n_291),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_290),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_294),
.B(n_295),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_314),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_314),
.Y(n_329)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_304),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_303)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_304),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_307),
.C(n_309),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_309),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_309),
.A2(n_311),
.B1(n_316),
.B2(n_320),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_320),
.C(n_321),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_312),
.A2(n_313),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_321),
.Y(n_314)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_323),
.B(n_324),
.Y(n_328)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_332),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_333),
.Y(n_335)
);


endmodule