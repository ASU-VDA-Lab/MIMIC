module fake_netlist_6_2049_n_1705 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1705);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1705;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_109),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_59),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_136),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_57),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_60),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_23),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_0),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_122),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_80),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_58),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_97),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_68),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_43),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_71),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_32),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_15),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_81),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_70),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_10),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_49),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_49),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_113),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_69),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_119),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_72),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_34),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_148),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_98),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_103),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_99),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_89),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g188 ( 
.A(n_60),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_111),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_39),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_131),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_141),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_16),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_92),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_54),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_45),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_145),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_138),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_108),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_105),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_61),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_1),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_6),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_0),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_56),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_110),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_46),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_27),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_66),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_102),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_25),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_17),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_26),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_64),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_67),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_2),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_8),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_100),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_95),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_10),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_139),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_22),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_29),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_9),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_146),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_47),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_65),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_112),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_50),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_27),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_90),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_118),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_142),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_34),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_58),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_64),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_29),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_123),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_149),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_30),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_152),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_61),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_115),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_28),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_18),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_45),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_74),
.Y(n_247)
);

CKINVDCx6p67_ASAP7_75t_R g248 ( 
.A(n_96),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_14),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_23),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_32),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_5),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_137),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_8),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_38),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_147),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_41),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_75),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_41),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_128),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_3),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_40),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_28),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_134),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_43),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_132),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_53),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_143),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_140),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_14),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_62),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_62),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_86),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_73),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_116),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_88),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_135),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_52),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_77),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_19),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_36),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_56),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_20),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_124),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_24),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_107),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_25),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_40),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_129),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_151),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_63),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_36),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_30),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_93),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_85),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_50),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_91),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_84),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_24),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_82),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_125),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_33),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_5),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_33),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_42),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_290),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_153),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_167),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_167),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_167),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_155),
.Y(n_311)
);

INVxp33_ASAP7_75t_SL g312 ( 
.A(n_154),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_161),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_1),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_167),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_167),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_167),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_165),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_168),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_171),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_173),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_170),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_158),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_170),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_157),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_170),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_179),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_170),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_170),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_180),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_159),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_188),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_170),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_223),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_216),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_216),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_183),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_216),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_216),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_166),
.B(n_172),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_185),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_157),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_216),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_186),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_216),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_240),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_240),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_166),
.B(n_2),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_187),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_160),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_172),
.B(n_3),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_156),
.B(n_4),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_189),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_240),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_240),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_240),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_199),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_240),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_200),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_201),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_201),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_254),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_209),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_210),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_215),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_254),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_219),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_295),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_288),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_223),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_188),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_288),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_223),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_280),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_280),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_176),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_221),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_227),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_280),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_232),
.Y(n_380)
);

NAND2xp33_ASAP7_75t_SL g381 ( 
.A(n_352),
.B(n_283),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_308),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_368),
.Y(n_383)
);

BUFx8_ASAP7_75t_L g384 ( 
.A(n_334),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_333),
.B(n_233),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_308),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_368),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_338),
.B(n_239),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_355),
.B(n_241),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_368),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_368),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_368),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_340),
.B(n_243),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_334),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_368),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_309),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_309),
.B(n_163),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_310),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_373),
.B(n_253),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_331),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_310),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_373),
.B(n_256),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_314),
.B(n_188),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_315),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_306),
.B(n_197),
.Y(n_405)
);

NOR2x1_ASAP7_75t_L g406 ( 
.A(n_337),
.B(n_156),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_315),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_316),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_260),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_316),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_317),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_317),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_322),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_322),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_374),
.B(n_283),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_324),
.B(n_163),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_324),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_312),
.B(n_225),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_348),
.B(n_238),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_332),
.B(n_188),
.Y(n_420)
);

AND2x6_ASAP7_75t_L g421 ( 
.A(n_326),
.B(n_156),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_326),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_370),
.B(n_287),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_375),
.B(n_264),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_375),
.B(n_266),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_328),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_379),
.B(n_273),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_328),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_329),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_379),
.B(n_287),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_329),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_335),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_335),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_336),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_336),
.B(n_276),
.Y(n_435)
);

OA21x2_ASAP7_75t_L g436 ( 
.A1(n_339),
.A2(n_205),
.B(n_176),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_339),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_343),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_343),
.B(n_277),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_345),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_345),
.B(n_279),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_346),
.B(n_286),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_346),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_347),
.B(n_289),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_347),
.B(n_297),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_354),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_351),
.A2(n_193),
.B1(n_255),
.B2(n_282),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_354),
.Y(n_448)
);

BUFx8_ASAP7_75t_L g449 ( 
.A(n_337),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_436),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_436),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_394),
.Y(n_452)
);

INVx5_ASAP7_75t_L g453 ( 
.A(n_421),
.Y(n_453)
);

AOI21x1_ASAP7_75t_L g454 ( 
.A1(n_382),
.A2(n_358),
.B(n_356),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_419),
.A2(n_287),
.B1(n_205),
.B2(n_208),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_408),
.Y(n_456)
);

AND2x6_ASAP7_75t_L g457 ( 
.A(n_406),
.B(n_162),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_385),
.B(n_311),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_408),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_443),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_385),
.B(n_313),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_408),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_391),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_408),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_391),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_436),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_436),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_436),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_436),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_382),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_391),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_423),
.B(n_360),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_419),
.A2(n_230),
.B1(n_208),
.B2(n_213),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_SL g474 ( 
.A1(n_384),
.A2(n_332),
.B1(n_371),
.B2(n_323),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_386),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_423),
.B(n_360),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_386),
.Y(n_477)
);

OR2x6_ASAP7_75t_L g478 ( 
.A(n_406),
.B(n_162),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_391),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_396),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_435),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_391),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_391),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_394),
.Y(n_484)
);

BUFx10_ASAP7_75t_L g485 ( 
.A(n_418),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_410),
.Y(n_486)
);

OAI22xp33_ASAP7_75t_L g487 ( 
.A1(n_403),
.A2(n_371),
.B1(n_207),
.B2(n_257),
.Y(n_487)
);

NAND2xp33_ASAP7_75t_L g488 ( 
.A(n_393),
.B(n_318),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_400),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_418),
.B(n_320),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_423),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_391),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_430),
.B(n_361),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_384),
.Y(n_494)
);

NAND2xp33_ASAP7_75t_L g495 ( 
.A(n_393),
.B(n_321),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_391),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_443),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_410),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_399),
.B(n_323),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_392),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_400),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_396),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_410),
.Y(n_503)
);

INVx6_ASAP7_75t_L g504 ( 
.A(n_397),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_384),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_384),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_392),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_398),
.Y(n_508)
);

AND2x6_ASAP7_75t_L g509 ( 
.A(n_397),
.B(n_162),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_398),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_405),
.B(n_327),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_412),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_403),
.A2(n_381),
.B1(n_405),
.B2(n_430),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_415),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_430),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_392),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_392),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_381),
.A2(n_226),
.B1(n_213),
.B2(n_214),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_392),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_415),
.Y(n_520)
);

INVx4_ASAP7_75t_SL g521 ( 
.A(n_421),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_404),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_399),
.B(n_361),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_421),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_404),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_407),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_402),
.B(n_362),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_397),
.B(n_178),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_412),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_402),
.B(n_174),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_397),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_388),
.B(n_341),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_407),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_409),
.B(n_362),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_412),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_447),
.A2(n_420),
.B1(n_226),
.B2(n_230),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_416),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_414),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_384),
.B(n_344),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_414),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_389),
.B(n_439),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_416),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_420),
.B(n_357),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_447),
.A2(n_220),
.B1(n_177),
.B2(n_175),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_412),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_422),
.Y(n_546)
);

INVx5_ASAP7_75t_L g547 ( 
.A(n_421),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_422),
.Y(n_548)
);

BUFx10_ASAP7_75t_L g549 ( 
.A(n_416),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_416),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_439),
.B(n_359),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_449),
.B(n_364),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_426),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_449),
.B(n_380),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_409),
.B(n_337),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_449),
.B(n_378),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_424),
.B(n_366),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_443),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_426),
.Y(n_559)
);

CKINVDCx11_ASAP7_75t_R g560 ( 
.A(n_416),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_449),
.B(n_307),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_424),
.B(n_366),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_440),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_428),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_L g565 ( 
.A(n_425),
.B(n_295),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_425),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_440),
.Y(n_567)
);

AO22x2_ASAP7_75t_L g568 ( 
.A1(n_415),
.A2(n_174),
.B1(n_184),
.B2(n_178),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_440),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_449),
.B(n_377),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_427),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_427),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_441),
.B(n_442),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_428),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_441),
.A2(n_214),
.B1(n_234),
.B2(n_235),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_442),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_429),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_392),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_444),
.B(n_198),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_444),
.B(n_319),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_445),
.Y(n_581)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_421),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_440),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_429),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_445),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_431),
.B(n_330),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_401),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_431),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_401),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_434),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_401),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_434),
.B(n_349),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_432),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_432),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_437),
.B(n_353),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_452),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_581),
.B(n_437),
.Y(n_597)
);

AO22x1_ASAP7_75t_L g598 ( 
.A1(n_536),
.A2(n_235),
.B1(n_234),
.B2(n_236),
.Y(n_598)
);

NAND2x1p5_ASAP7_75t_L g599 ( 
.A(n_491),
.B(n_198),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_581),
.B(n_446),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_499),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_493),
.B(n_325),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_451),
.A2(n_466),
.B1(n_467),
.B2(n_450),
.Y(n_603)
);

NAND3xp33_ASAP7_75t_L g604 ( 
.A(n_513),
.B(n_350),
.C(n_363),
.Y(n_604)
);

NAND3xp33_ASAP7_75t_SL g605 ( 
.A(n_544),
.B(n_367),
.C(n_365),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_484),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_585),
.B(n_446),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_585),
.B(n_448),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_485),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_571),
.B(n_295),
.Y(n_610)
);

NOR3xp33_ASAP7_75t_L g611 ( 
.A(n_536),
.B(n_376),
.C(n_342),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_481),
.B(n_448),
.Y(n_612)
);

NOR2xp67_ASAP7_75t_L g613 ( 
.A(n_501),
.B(n_298),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_456),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_456),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_571),
.B(n_258),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_572),
.B(n_541),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_L g618 ( 
.A(n_576),
.B(n_191),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_456),
.Y(n_619)
);

NAND3xp33_ASAP7_75t_L g620 ( 
.A(n_473),
.B(n_169),
.C(n_164),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_491),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_459),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_514),
.B(n_261),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_572),
.B(n_182),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_573),
.B(n_411),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_491),
.B(n_295),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_531),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_566),
.B(n_190),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_532),
.B(n_411),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_566),
.A2(n_184),
.B1(n_174),
.B2(n_192),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_499),
.B(n_195),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_514),
.B(n_196),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_531),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_537),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_451),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_555),
.B(n_411),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_504),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_580),
.A2(n_300),
.B1(n_206),
.B2(n_301),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_537),
.Y(n_639)
);

BUFx6f_ASAP7_75t_SL g640 ( 
.A(n_501),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_537),
.Y(n_641)
);

AND2x4_ASAP7_75t_SL g642 ( 
.A(n_484),
.B(n_248),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_542),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_459),
.Y(n_644)
);

INVx4_ASAP7_75t_SL g645 ( 
.A(n_509),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_459),
.Y(n_646)
);

INVxp67_ASAP7_75t_L g647 ( 
.A(n_489),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_523),
.B(n_527),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_579),
.B(n_295),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_489),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_452),
.B(n_202),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_579),
.B(n_295),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_527),
.B(n_413),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_520),
.B(n_203),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_520),
.B(n_204),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_515),
.B(n_261),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_462),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_534),
.B(n_413),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_451),
.A2(n_293),
.B1(n_271),
.B2(n_236),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_542),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_458),
.B(n_211),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_534),
.B(n_557),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_550),
.Y(n_663)
);

AOI221xp5_ASAP7_75t_L g664 ( 
.A1(n_487),
.A2(n_237),
.B1(n_245),
.B2(n_265),
.C(n_271),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_592),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_579),
.B(n_191),
.Y(n_666)
);

OAI22xp33_ASAP7_75t_L g667 ( 
.A1(n_515),
.A2(n_293),
.B1(n_265),
.B2(n_305),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_550),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_550),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_493),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_562),
.B(n_461),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_470),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_511),
.B(n_212),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_470),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_579),
.B(n_191),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_475),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_551),
.B(n_417),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_588),
.B(n_417),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_475),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_549),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_490),
.B(n_217),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_549),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_586),
.B(n_595),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_485),
.B(n_222),
.Y(n_684)
);

NAND3xp33_ASAP7_75t_L g685 ( 
.A(n_455),
.B(n_272),
.C(n_224),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_485),
.B(n_229),
.Y(n_686)
);

OR2x6_ASAP7_75t_L g687 ( 
.A(n_505),
.B(n_237),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_485),
.B(n_242),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_477),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_477),
.Y(n_690)
);

INVx1_ASAP7_75t_SL g691 ( 
.A(n_472),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_543),
.B(n_244),
.Y(n_692)
);

OR2x6_ASAP7_75t_L g693 ( 
.A(n_505),
.B(n_245),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_588),
.B(n_417),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_488),
.B(n_246),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_450),
.B(n_191),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_495),
.A2(n_274),
.B1(n_206),
.B2(n_218),
.Y(n_697)
);

INVx5_ASAP7_75t_L g698 ( 
.A(n_509),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_588),
.B(n_417),
.Y(n_699)
);

OAI21xp33_ASAP7_75t_L g700 ( 
.A1(n_476),
.A2(n_305),
.B(n_267),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_462),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_480),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_476),
.B(n_249),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_544),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_504),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_474),
.B(n_261),
.Y(n_706)
);

BUFx5_ASAP7_75t_L g707 ( 
.A(n_467),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_480),
.B(n_250),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_468),
.B(n_191),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_530),
.A2(n_284),
.B1(n_218),
.B2(n_228),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_469),
.A2(n_565),
.B(n_471),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_469),
.B(n_191),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_502),
.B(n_395),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_502),
.B(n_251),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_508),
.B(n_395),
.Y(n_715)
);

INVx1_ASAP7_75t_SL g716 ( 
.A(n_560),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_549),
.B(n_191),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_508),
.B(n_252),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_539),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_464),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_464),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_510),
.B(n_259),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_530),
.A2(n_294),
.B1(n_284),
.B2(n_275),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_464),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_510),
.B(n_228),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_575),
.B(n_262),
.Y(n_726)
);

INVxp67_ASAP7_75t_SL g727 ( 
.A(n_465),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_522),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_528),
.B(n_231),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_525),
.B(n_231),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_525),
.B(n_247),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_526),
.B(n_263),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_533),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_533),
.B(n_247),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_504),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_538),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_540),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_540),
.B(n_270),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_546),
.B(n_278),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_504),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_494),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_528),
.B(n_269),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_506),
.B(n_518),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_530),
.A2(n_269),
.B1(n_294),
.B2(n_275),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_549),
.B(n_191),
.Y(n_745)
);

INVxp67_ASAP7_75t_L g746 ( 
.A(n_528),
.Y(n_746)
);

BUFx2_ASAP7_75t_L g747 ( 
.A(n_596),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_671),
.B(n_548),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_741),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_648),
.A2(n_530),
.B1(n_504),
.B2(n_554),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_662),
.B(n_553),
.Y(n_751)
);

OAI21xp33_ASAP7_75t_L g752 ( 
.A1(n_683),
.A2(n_285),
.B(n_281),
.Y(n_752)
);

O2A1O1Ixp5_ASAP7_75t_L g753 ( 
.A1(n_636),
.A2(n_559),
.B(n_564),
.C(n_553),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_616),
.B(n_617),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_650),
.Y(n_755)
);

NOR2xp67_ASAP7_75t_L g756 ( 
.A(n_647),
.B(n_552),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_606),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_711),
.A2(n_482),
.B(n_463),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_707),
.B(n_528),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_616),
.B(n_559),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_621),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_L g762 ( 
.A1(n_696),
.A2(n_530),
.B(n_564),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_617),
.B(n_574),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_683),
.A2(n_556),
.B1(n_570),
.B2(n_561),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_602),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_625),
.A2(n_482),
.B(n_516),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_707),
.B(n_574),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_661),
.B(n_577),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_661),
.B(n_577),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_698),
.A2(n_482),
.B(n_463),
.Y(n_770)
);

BUFx12f_ASAP7_75t_L g771 ( 
.A(n_651),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_624),
.B(n_478),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_664),
.A2(n_659),
.B(n_704),
.C(n_631),
.Y(n_773)
);

A2O1A1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_673),
.A2(n_590),
.B(n_584),
.C(n_274),
.Y(n_774)
);

NOR3xp33_ASAP7_75t_L g775 ( 
.A(n_605),
.B(n_301),
.C(n_590),
.Y(n_775)
);

AND2x2_ASAP7_75t_SL g776 ( 
.A(n_659),
.B(n_184),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_635),
.Y(n_777)
);

OR2x6_ASAP7_75t_L g778 ( 
.A(n_687),
.B(n_478),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_698),
.A2(n_578),
.B(n_516),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_707),
.B(n_584),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_601),
.B(n_478),
.Y(n_781)
);

OAI21xp33_ASAP7_75t_L g782 ( 
.A1(n_631),
.A2(n_624),
.B(n_632),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_698),
.A2(n_482),
.B(n_516),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_672),
.Y(n_784)
);

O2A1O1Ixp5_ASAP7_75t_L g785 ( 
.A1(n_696),
.A2(n_454),
.B(n_593),
.C(n_591),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_707),
.B(n_463),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_674),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_629),
.A2(n_516),
.B(n_519),
.Y(n_788)
);

NAND3xp33_ASAP7_75t_L g789 ( 
.A(n_638),
.B(n_478),
.C(n_292),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_691),
.B(n_478),
.Y(n_790)
);

NOR2x1p5_ASAP7_75t_L g791 ( 
.A(n_604),
.B(n_609),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_623),
.B(n_568),
.Y(n_792)
);

INVx4_ASAP7_75t_L g793 ( 
.A(n_680),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_655),
.B(n_291),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_670),
.B(n_521),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_653),
.A2(n_519),
.B(n_463),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_707),
.B(n_457),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_707),
.B(n_457),
.Y(n_798)
);

A2O1A1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_673),
.A2(n_268),
.B(n_192),
.C(n_194),
.Y(n_799)
);

INVx6_ASAP7_75t_L g800 ( 
.A(n_602),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_658),
.A2(n_519),
.B(n_578),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_665),
.B(n_465),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_681),
.A2(n_268),
.B(n_194),
.C(n_181),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_709),
.A2(n_492),
.B(n_465),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_603),
.B(n_519),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_676),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_687),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_677),
.A2(n_519),
.B(n_578),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_679),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_612),
.A2(n_578),
.B(n_497),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_689),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_690),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_632),
.B(n_465),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_680),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_637),
.A2(n_578),
.B(n_558),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_637),
.A2(n_558),
.B(n_497),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_702),
.B(n_457),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_728),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_705),
.Y(n_819)
);

A2O1A1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_681),
.A2(n_181),
.B(n_471),
.C(n_479),
.Y(n_820)
);

O2A1O1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_610),
.A2(n_594),
.B(n_591),
.C(n_589),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_712),
.A2(n_492),
.B(n_471),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_735),
.A2(n_558),
.B(n_460),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_611),
.A2(n_568),
.B1(n_457),
.B2(n_509),
.Y(n_824)
);

INVx4_ASAP7_75t_L g825 ( 
.A(n_680),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_735),
.A2(n_727),
.B(n_694),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_680),
.B(n_471),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_678),
.A2(n_497),
.B(n_558),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_699),
.A2(n_460),
.B(n_497),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_733),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_736),
.B(n_457),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_682),
.A2(n_460),
.B(n_492),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_682),
.A2(n_460),
.B(n_492),
.Y(n_833)
);

OAI21xp5_ASAP7_75t_L g834 ( 
.A1(n_626),
.A2(n_483),
.B(n_479),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_626),
.A2(n_483),
.B(n_479),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_610),
.A2(n_483),
.B(n_479),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_737),
.B(n_496),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_716),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_654),
.B(n_496),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_597),
.B(n_600),
.Y(n_840)
);

NOR2x1_ASAP7_75t_R g841 ( 
.A(n_706),
.B(n_296),
.Y(n_841)
);

A2O1A1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_695),
.A2(n_496),
.B(n_500),
.C(n_507),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_630),
.A2(n_589),
.B(n_587),
.C(n_583),
.Y(n_843)
);

INVx5_ASAP7_75t_L g844 ( 
.A(n_660),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_607),
.B(n_500),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_746),
.A2(n_568),
.B1(n_500),
.B2(n_507),
.Y(n_846)
);

INVx1_ASAP7_75t_SL g847 ( 
.A(n_642),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_641),
.B(n_521),
.Y(n_848)
);

OR2x2_ASAP7_75t_L g849 ( 
.A(n_654),
.B(n_299),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_641),
.B(n_521),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_717),
.A2(n_500),
.B(n_517),
.Y(n_851)
);

AND2x6_ASAP7_75t_L g852 ( 
.A(n_705),
.B(n_507),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_717),
.A2(n_745),
.B(n_660),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_628),
.B(n_568),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_745),
.A2(n_517),
.B(n_507),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_608),
.B(n_509),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_703),
.B(n_509),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_628),
.B(n_302),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_703),
.B(n_509),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_645),
.B(n_453),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_713),
.A2(n_715),
.B(n_740),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_684),
.B(n_303),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_740),
.A2(n_392),
.B(n_582),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_627),
.A2(n_392),
.B(n_582),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_656),
.B(n_568),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_633),
.A2(n_453),
.B(n_582),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_708),
.B(n_509),
.Y(n_867)
);

O2A1O1Ixp5_ASAP7_75t_L g868 ( 
.A1(n_666),
.A2(n_589),
.B(n_587),
.C(n_583),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_634),
.A2(n_453),
.B(n_582),
.Y(n_869)
);

O2A1O1Ixp33_ASAP7_75t_SL g870 ( 
.A1(n_649),
.A2(n_486),
.B(n_583),
.C(n_569),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_708),
.B(n_509),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_642),
.Y(n_872)
);

O2A1O1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_618),
.A2(n_587),
.B(n_569),
.C(n_567),
.Y(n_873)
);

NOR3xp33_ASAP7_75t_L g874 ( 
.A(n_684),
.B(n_304),
.C(n_372),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_639),
.A2(n_582),
.B(n_453),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_643),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_599),
.A2(n_248),
.B1(n_569),
.B2(n_567),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_663),
.A2(n_582),
.B(n_453),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_666),
.A2(n_567),
.B(n_563),
.C(n_486),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_714),
.B(n_486),
.Y(n_880)
);

A2O1A1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_695),
.A2(n_498),
.B(n_563),
.C(n_503),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_714),
.B(n_498),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_686),
.B(n_498),
.Y(n_883)
);

INVx6_ASAP7_75t_L g884 ( 
.A(n_729),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_718),
.B(n_503),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_729),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_645),
.B(n_453),
.Y(n_887)
);

O2A1O1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_675),
.A2(n_545),
.B(n_535),
.C(n_529),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_692),
.A2(n_529),
.B(n_512),
.C(n_545),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_718),
.B(n_503),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_722),
.B(n_512),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_692),
.A2(n_535),
.B(n_529),
.C(n_512),
.Y(n_892)
);

A2O1A1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_722),
.A2(n_369),
.B(n_372),
.C(n_358),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_668),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_599),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_732),
.B(n_432),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_686),
.B(n_4),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_726),
.B(n_688),
.Y(n_898)
);

NAND3xp33_ASAP7_75t_L g899 ( 
.A(n_688),
.B(n_738),
.C(n_732),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_719),
.B(n_6),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_614),
.A2(n_390),
.B(n_387),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_743),
.B(n_369),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_738),
.B(n_438),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_739),
.B(n_742),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_669),
.A2(n_582),
.B(n_547),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_742),
.A2(n_421),
.B1(n_521),
.B2(n_433),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_739),
.A2(n_356),
.B(n_433),
.C(n_438),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_649),
.A2(n_547),
.B(n_524),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_SL g909 ( 
.A1(n_652),
.A2(n_390),
.B(n_387),
.C(n_383),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_652),
.A2(n_547),
.B(n_524),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_697),
.A2(n_723),
.B(n_710),
.C(n_744),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_615),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_619),
.A2(n_547),
.B(n_524),
.Y(n_913)
);

NOR2x1p5_ASAP7_75t_SL g914 ( 
.A(n_622),
.B(n_644),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_646),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_754),
.B(n_613),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_886),
.B(n_645),
.Y(n_917)
);

AO21x1_ASAP7_75t_L g918 ( 
.A1(n_897),
.A2(n_734),
.B(n_731),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_782),
.B(n_898),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_899),
.A2(n_640),
.B1(n_687),
.B2(n_693),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_747),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_773),
.A2(n_640),
.B1(n_693),
.B2(n_725),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_755),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_772),
.B(n_657),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_777),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_858),
.B(n_700),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_776),
.A2(n_667),
.B1(n_685),
.B2(n_620),
.Y(n_927)
);

O2A1O1Ixp33_ASAP7_75t_SL g928 ( 
.A1(n_773),
.A2(n_667),
.B(n_730),
.C(n_721),
.Y(n_928)
);

O2A1O1Ixp5_ASAP7_75t_L g929 ( 
.A1(n_862),
.A2(n_598),
.B(n_720),
.C(n_701),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_858),
.B(n_693),
.Y(n_930)
);

CKINVDCx16_ASAP7_75t_R g931 ( 
.A(n_838),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_840),
.B(n_724),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_765),
.B(n_521),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_760),
.B(n_438),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_755),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_748),
.B(n_433),
.Y(n_936)
);

OR2x6_ASAP7_75t_L g937 ( 
.A(n_778),
.B(n_443),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_768),
.B(n_421),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_749),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_800),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_759),
.A2(n_547),
.B(n_524),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_L g942 ( 
.A1(n_776),
.A2(n_897),
.B1(n_854),
.B2(n_862),
.Y(n_942)
);

INVxp67_ASAP7_75t_SL g943 ( 
.A(n_814),
.Y(n_943)
);

A2O1A1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_900),
.A2(n_390),
.B(n_387),
.C(n_383),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_769),
.B(n_421),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_771),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_761),
.B(n_120),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_904),
.A2(n_547),
.B1(n_524),
.B2(n_453),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_784),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_800),
.Y(n_950)
);

AOI33xp33_ASAP7_75t_L g951 ( 
.A1(n_787),
.A2(n_261),
.A3(n_9),
.B1(n_11),
.B2(n_12),
.B3(n_13),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_814),
.Y(n_952)
);

OR2x4_ASAP7_75t_L g953 ( 
.A(n_900),
.B(n_7),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_800),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_874),
.A2(n_421),
.B1(n_443),
.B2(n_383),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_874),
.A2(n_421),
.B1(n_443),
.B2(n_383),
.Y(n_956)
);

NOR3xp33_ASAP7_75t_SL g957 ( 
.A(n_752),
.B(n_7),
.C(n_11),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_814),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_857),
.B(n_443),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_849),
.A2(n_12),
.B(n_13),
.C(n_15),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_859),
.B(n_867),
.Y(n_961)
);

O2A1O1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_775),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_806),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_781),
.B(n_19),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_775),
.A2(n_443),
.B1(n_150),
.B2(n_133),
.Y(n_965)
);

NOR2xp67_ASAP7_75t_SL g966 ( 
.A(n_844),
.B(n_20),
.Y(n_966)
);

INVx4_ASAP7_75t_L g967 ( 
.A(n_848),
.Y(n_967)
);

AND2x4_ASAP7_75t_SL g968 ( 
.A(n_793),
.B(n_130),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_751),
.B(n_21),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_757),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_813),
.A2(n_127),
.B1(n_126),
.B2(n_117),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_848),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_902),
.B(n_21),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_790),
.B(n_22),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_850),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_809),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_850),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_805),
.A2(n_104),
.B(n_101),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_763),
.B(n_26),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_807),
.Y(n_980)
);

OAI21xp33_ASAP7_75t_L g981 ( 
.A1(n_794),
.A2(n_31),
.B(n_35),
.Y(n_981)
);

INVxp67_ASAP7_75t_SL g982 ( 
.A(n_819),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_811),
.Y(n_983)
);

INVxp67_ASAP7_75t_L g984 ( 
.A(n_841),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_813),
.A2(n_94),
.B1(n_87),
.B2(n_83),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_912),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_839),
.B(n_31),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_911),
.A2(n_35),
.B(n_37),
.C(n_38),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_884),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_812),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_871),
.B(n_79),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_839),
.B(n_37),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_818),
.B(n_39),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_815),
.A2(n_78),
.B(n_76),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_894),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_778),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_830),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_883),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_802),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_792),
.A2(n_762),
.B(n_753),
.C(n_865),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_802),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_895),
.B(n_48),
.Y(n_1002)
);

NOR2xp67_ASAP7_75t_SL g1003 ( 
.A(n_844),
.B(n_51),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_780),
.A2(n_797),
.B(n_798),
.Y(n_1004)
);

NAND2xp33_ASAP7_75t_R g1005 ( 
.A(n_778),
.B(n_51),
.Y(n_1005)
);

INVx4_ASAP7_75t_L g1006 ( 
.A(n_793),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_895),
.B(n_880),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_756),
.B(n_52),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_882),
.B(n_53),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_753),
.A2(n_54),
.B(n_55),
.C(n_57),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_872),
.B(n_55),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_805),
.A2(n_844),
.B1(n_884),
.B2(n_750),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_844),
.B(n_59),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_SL g1014 ( 
.A(n_847),
.B(n_63),
.Y(n_1014)
);

BUFx4f_ASAP7_75t_SL g1015 ( 
.A(n_825),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_876),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_789),
.A2(n_853),
.B(n_774),
.C(n_891),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_791),
.B(n_884),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_885),
.A2(n_890),
.B1(n_856),
.B2(n_819),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_894),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_837),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_896),
.B(n_903),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_799),
.A2(n_803),
.B(n_868),
.C(n_817),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_825),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_795),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_810),
.A2(n_826),
.B(n_786),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_915),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_845),
.B(n_795),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_785),
.Y(n_1029)
);

NAND3xp33_ASAP7_75t_SL g1030 ( 
.A(n_824),
.B(n_831),
.C(n_861),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_767),
.B(n_852),
.Y(n_1031)
);

NAND2x1p5_ASAP7_75t_L g1032 ( 
.A(n_827),
.B(n_860),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_915),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_915),
.B(n_786),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_816),
.A2(n_823),
.B(n_788),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_852),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_758),
.A2(n_808),
.B(n_766),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_868),
.A2(n_785),
.B(n_824),
.C(n_879),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_843),
.Y(n_1039)
);

OAI22x1_ASAP7_75t_L g1040 ( 
.A1(n_906),
.A2(n_846),
.B1(n_860),
.B2(n_887),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_852),
.B(n_801),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_821),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_804),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_822),
.B(n_835),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_SL g1045 ( 
.A1(n_877),
.A2(n_836),
.B1(n_834),
.B2(n_901),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_851),
.B(n_855),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_796),
.B(n_889),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_949),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_1022),
.A2(n_833),
.B(n_832),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_1035),
.A2(n_828),
.B(n_829),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_921),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_926),
.A2(n_930),
.B1(n_919),
.B2(n_942),
.Y(n_1052)
);

INVx4_ASAP7_75t_L g1053 ( 
.A(n_1015),
.Y(n_1053)
);

OAI221xp5_ASAP7_75t_L g1054 ( 
.A1(n_926),
.A2(n_893),
.B1(n_820),
.B2(n_907),
.C(n_842),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_961),
.A2(n_1026),
.B(n_1037),
.Y(n_1055)
);

INVx2_ASAP7_75t_SL g1056 ( 
.A(n_921),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_919),
.B(n_892),
.Y(n_1057)
);

NOR4xp25_ASAP7_75t_L g1058 ( 
.A(n_960),
.B(n_881),
.C(n_870),
.D(n_873),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_988),
.A2(n_909),
.B(n_870),
.C(n_888),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_970),
.Y(n_1060)
);

AOI21x1_ASAP7_75t_L g1061 ( 
.A1(n_959),
.A2(n_770),
.B(n_779),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_SL g1062 ( 
.A(n_939),
.B(n_910),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_942),
.A2(n_783),
.B1(n_864),
.B2(n_863),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_980),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_961),
.A2(n_866),
.B(n_869),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_969),
.A2(n_914),
.B(n_878),
.C(n_905),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_927),
.A2(n_875),
.B1(n_908),
.B2(n_913),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_969),
.A2(n_909),
.B(n_916),
.C(n_987),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_1047),
.A2(n_1019),
.B(n_1017),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_923),
.B(n_935),
.Y(n_1070)
);

OR2x6_ASAP7_75t_L g1071 ( 
.A(n_937),
.B(n_939),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_1017),
.A2(n_1041),
.B(n_1004),
.Y(n_1072)
);

CKINVDCx11_ASAP7_75t_R g1073 ( 
.A(n_931),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_1046),
.A2(n_1045),
.B(n_959),
.Y(n_1074)
);

OAI22x1_ASAP7_75t_L g1075 ( 
.A1(n_974),
.A2(n_964),
.B1(n_996),
.B2(n_1013),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_970),
.B(n_1027),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_963),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_976),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_974),
.B(n_964),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1044),
.A2(n_1030),
.B(n_932),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_983),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_973),
.B(n_1016),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1007),
.B(n_999),
.Y(n_1083)
);

AO21x2_ASAP7_75t_L g1084 ( 
.A1(n_918),
.A2(n_944),
.B(n_1038),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_992),
.A2(n_927),
.B(n_978),
.C(n_981),
.Y(n_1085)
);

AOI21x1_ASAP7_75t_L g1086 ( 
.A1(n_991),
.A2(n_1044),
.B(n_924),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_1032),
.A2(n_991),
.B(n_924),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_1001),
.B(n_920),
.Y(n_1088)
);

INVx3_ASAP7_75t_SL g1089 ( 
.A(n_1011),
.Y(n_1089)
);

BUFx4_ASAP7_75t_SL g1090 ( 
.A(n_946),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1038),
.A2(n_936),
.B(n_1029),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_SL g1092 ( 
.A1(n_962),
.A2(n_994),
.B(n_1031),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1029),
.A2(n_934),
.B(n_1028),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_922),
.A2(n_988),
.B(n_1009),
.C(n_929),
.Y(n_1094)
);

BUFx4_ASAP7_75t_SL g1095 ( 
.A(n_940),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_979),
.A2(n_1000),
.B(n_965),
.C(n_1034),
.Y(n_1096)
);

AO22x2_ASAP7_75t_L g1097 ( 
.A1(n_998),
.A2(n_1013),
.B1(n_1008),
.B2(n_1002),
.Y(n_1097)
);

AO31x2_ASAP7_75t_L g1098 ( 
.A1(n_944),
.A2(n_1023),
.A3(n_1000),
.B(n_1010),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_1034),
.A2(n_957),
.B(n_993),
.C(n_1021),
.Y(n_1099)
);

AO31x2_ASAP7_75t_L g1100 ( 
.A1(n_1023),
.A2(n_1010),
.A3(n_1040),
.B(n_1042),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_SL g1101 ( 
.A1(n_971),
.A2(n_985),
.B(n_1039),
.C(n_945),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_928),
.A2(n_938),
.B(n_1043),
.Y(n_1102)
);

INVxp67_ASAP7_75t_L g1103 ( 
.A(n_1014),
.Y(n_1103)
);

OA21x2_ASAP7_75t_L g1104 ( 
.A1(n_956),
.A2(n_955),
.B(n_1020),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_990),
.B(n_997),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1036),
.A2(n_982),
.B(n_943),
.Y(n_1106)
);

OR2x6_ASAP7_75t_L g1107 ( 
.A(n_937),
.B(n_1024),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_940),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_941),
.A2(n_948),
.B(n_937),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_1015),
.B(n_1024),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_956),
.A2(n_925),
.B(n_986),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_947),
.A2(n_1025),
.B(n_995),
.C(n_951),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_958),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_950),
.B(n_954),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_953),
.A2(n_947),
.B1(n_968),
.B2(n_975),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_968),
.A2(n_1024),
.B(n_1033),
.Y(n_1116)
);

NAND3xp33_ASAP7_75t_L g1117 ( 
.A(n_1005),
.B(n_951),
.C(n_1003),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_972),
.B(n_977),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_1011),
.A2(n_984),
.B(n_1018),
.C(n_989),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_972),
.B(n_977),
.Y(n_1120)
);

BUFx12f_ASAP7_75t_L g1121 ( 
.A(n_958),
.Y(n_1121)
);

AO21x2_ASAP7_75t_L g1122 ( 
.A1(n_917),
.A2(n_966),
.B(n_933),
.Y(n_1122)
);

AO21x2_ASAP7_75t_L g1123 ( 
.A1(n_917),
.A2(n_933),
.B(n_953),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_967),
.B(n_975),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_967),
.B(n_975),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1006),
.A2(n_952),
.B(n_975),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_989),
.A2(n_950),
.B(n_954),
.C(n_1005),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_972),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_977),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1006),
.A2(n_1022),
.B(n_961),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_SL g1131 ( 
.A(n_926),
.B(n_782),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1035),
.A2(n_1037),
.B(n_1026),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1035),
.A2(n_1037),
.B(n_1026),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_989),
.B(n_940),
.Y(n_1134)
);

INVx4_ASAP7_75t_L g1135 ( 
.A(n_1015),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_919),
.B(n_671),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_930),
.B(n_601),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_919),
.B(n_683),
.Y(n_1138)
);

INVxp67_ASAP7_75t_SL g1139 ( 
.A(n_921),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_921),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_926),
.A2(n_683),
.B(n_782),
.C(n_862),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1022),
.A2(n_961),
.B(n_1026),
.Y(n_1142)
);

AOI221x1_ASAP7_75t_L g1143 ( 
.A1(n_988),
.A2(n_782),
.B1(n_897),
.B2(n_899),
.C(n_683),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1022),
.A2(n_961),
.B(n_1026),
.Y(n_1144)
);

AO32x2_ASAP7_75t_L g1145 ( 
.A1(n_1012),
.A2(n_922),
.A3(n_998),
.B1(n_1045),
.B2(n_536),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1022),
.A2(n_961),
.B(n_1026),
.Y(n_1146)
);

BUFx10_ASAP7_75t_L g1147 ( 
.A(n_953),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_919),
.B(n_683),
.Y(n_1148)
);

NAND3xp33_ASAP7_75t_L g1149 ( 
.A(n_926),
.B(n_683),
.C(n_782),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_919),
.B(n_671),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1035),
.A2(n_1037),
.B(n_1026),
.Y(n_1151)
);

OAI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_926),
.A2(n_683),
.B1(n_899),
.B2(n_764),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_926),
.A2(n_683),
.B1(n_782),
.B2(n_899),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_926),
.A2(n_782),
.B(n_683),
.C(n_899),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1017),
.A2(n_899),
.B(n_926),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_926),
.A2(n_782),
.B(n_683),
.C(n_899),
.Y(n_1156)
);

INVxp67_ASAP7_75t_SL g1157 ( 
.A(n_921),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_919),
.B(n_671),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_926),
.A2(n_683),
.B1(n_782),
.B2(n_858),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1035),
.A2(n_1037),
.B(n_1026),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1017),
.A2(n_899),
.B(n_926),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_921),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_926),
.A2(n_683),
.B(n_782),
.C(n_862),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1022),
.A2(n_961),
.B(n_1026),
.Y(n_1164)
);

AO21x1_ASAP7_75t_L g1165 ( 
.A1(n_926),
.A2(n_897),
.B(n_987),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_926),
.A2(n_782),
.B(n_683),
.C(n_899),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_918),
.A2(n_944),
.A3(n_1038),
.B(n_1023),
.Y(n_1167)
);

AOI21xp33_ASAP7_75t_L g1168 ( 
.A1(n_926),
.A2(n_782),
.B(n_899),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1022),
.A2(n_961),
.B(n_1026),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1022),
.A2(n_961),
.B(n_1026),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_R g1171 ( 
.A(n_931),
.B(n_749),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1035),
.A2(n_1037),
.B(n_1026),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_921),
.Y(n_1173)
);

AO21x1_ASAP7_75t_L g1174 ( 
.A1(n_926),
.A2(n_897),
.B(n_987),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_918),
.A2(n_944),
.A3(n_1038),
.B(n_1023),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_926),
.A2(n_683),
.B(n_782),
.C(n_862),
.Y(n_1176)
);

OAI22x1_ASAP7_75t_L g1177 ( 
.A1(n_926),
.A2(n_764),
.B1(n_683),
.B2(n_897),
.Y(n_1177)
);

AO32x2_ASAP7_75t_L g1178 ( 
.A1(n_1012),
.A2(n_922),
.A3(n_998),
.B1(n_1045),
.B2(n_536),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_942),
.A2(n_776),
.B1(n_773),
.B2(n_659),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_1100),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1177),
.A2(n_1149),
.B1(n_1131),
.B2(n_1159),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1149),
.A2(n_1152),
.B1(n_1079),
.B2(n_1153),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1148),
.A2(n_1176),
.B1(n_1141),
.B2(n_1163),
.Y(n_1183)
);

INVx6_ASAP7_75t_L g1184 ( 
.A(n_1053),
.Y(n_1184)
);

NAND2xp33_ASAP7_75t_SL g1185 ( 
.A(n_1171),
.B(n_1053),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_1121),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1105),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1048),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1052),
.A2(n_1156),
.B1(n_1154),
.B2(n_1166),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1077),
.Y(n_1190)
);

NAND2x1p5_ASAP7_75t_L g1191 ( 
.A(n_1110),
.B(n_1135),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1179),
.A2(n_1088),
.B1(n_1085),
.B2(n_1138),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1131),
.A2(n_1179),
.B1(n_1168),
.B2(n_1155),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1137),
.B(n_1082),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1136),
.A2(n_1150),
.B1(n_1158),
.B2(n_1099),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_SL g1196 ( 
.A1(n_1117),
.A2(n_1161),
.B1(n_1155),
.B2(n_1115),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1078),
.Y(n_1197)
);

CKINVDCx11_ASAP7_75t_R g1198 ( 
.A(n_1073),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_SL g1199 ( 
.A1(n_1117),
.A2(n_1161),
.B1(n_1115),
.B2(n_1158),
.Y(n_1199)
);

CKINVDCx11_ASAP7_75t_R g1200 ( 
.A(n_1108),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_1140),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1168),
.A2(n_1165),
.B1(n_1174),
.B2(n_1075),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1081),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_1064),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1136),
.A2(n_1150),
.B1(n_1071),
.B2(n_1083),
.Y(n_1205)
);

BUFx8_ASAP7_75t_L g1206 ( 
.A(n_1051),
.Y(n_1206)
);

INVx6_ASAP7_75t_L g1207 ( 
.A(n_1135),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_SL g1208 ( 
.A1(n_1097),
.A2(n_1147),
.B1(n_1123),
.B2(n_1103),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_SL g1209 ( 
.A1(n_1097),
.A2(n_1147),
.B1(n_1123),
.B2(n_1083),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1071),
.A2(n_1139),
.B1(n_1157),
.B2(n_1107),
.Y(n_1210)
);

CKINVDCx11_ASAP7_75t_R g1211 ( 
.A(n_1089),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_1134),
.Y(n_1212)
);

OAI21xp33_ASAP7_75t_SL g1213 ( 
.A1(n_1107),
.A2(n_1057),
.B(n_1087),
.Y(n_1213)
);

CKINVDCx11_ASAP7_75t_R g1214 ( 
.A(n_1090),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1162),
.B(n_1076),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1056),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1071),
.A2(n_1112),
.B1(n_1096),
.B2(n_1070),
.Y(n_1217)
);

INVx4_ASAP7_75t_L g1218 ( 
.A(n_1113),
.Y(n_1218)
);

CKINVDCx14_ASAP7_75t_R g1219 ( 
.A(n_1114),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_1173),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1057),
.A2(n_1069),
.B1(n_1092),
.B2(n_1074),
.Y(n_1221)
);

BUFx8_ASAP7_75t_L g1222 ( 
.A(n_1060),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1094),
.A2(n_1119),
.B1(n_1127),
.B2(n_1116),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1084),
.A2(n_1080),
.B1(n_1054),
.B2(n_1072),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1084),
.A2(n_1130),
.B1(n_1143),
.B2(n_1062),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_1113),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1111),
.Y(n_1227)
);

INVx5_ASAP7_75t_L g1228 ( 
.A(n_1113),
.Y(n_1228)
);

OAI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1145),
.A2(n_1178),
.B1(n_1120),
.B2(n_1118),
.Y(n_1229)
);

CKINVDCx6p67_ASAP7_75t_R g1230 ( 
.A(n_1129),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1091),
.A2(n_1093),
.B1(n_1122),
.B2(n_1169),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1128),
.Y(n_1232)
);

CKINVDCx6p67_ASAP7_75t_R g1233 ( 
.A(n_1118),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_1120),
.Y(n_1234)
);

INVx6_ASAP7_75t_L g1235 ( 
.A(n_1095),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_SL g1236 ( 
.A1(n_1145),
.A2(n_1178),
.B1(n_1063),
.B2(n_1104),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1100),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1068),
.A2(n_1125),
.B1(n_1124),
.B2(n_1106),
.Y(n_1238)
);

INVx6_ASAP7_75t_L g1239 ( 
.A(n_1126),
.Y(n_1239)
);

BUFx8_ASAP7_75t_L g1240 ( 
.A(n_1145),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1086),
.B(n_1101),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_SL g1242 ( 
.A1(n_1178),
.A2(n_1063),
.B1(n_1104),
.B2(n_1067),
.Y(n_1242)
);

OAI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1102),
.A2(n_1142),
.B1(n_1170),
.B2(n_1144),
.Y(n_1243)
);

AOI21xp33_ASAP7_75t_L g1244 ( 
.A1(n_1059),
.A2(n_1067),
.B(n_1164),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_SL g1245 ( 
.A1(n_1146),
.A2(n_1098),
.B1(n_1055),
.B2(n_1109),
.Y(n_1245)
);

BUFx10_ASAP7_75t_L g1246 ( 
.A(n_1058),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_SL g1247 ( 
.A1(n_1098),
.A2(n_1175),
.B1(n_1167),
.B2(n_1160),
.Y(n_1247)
);

OAI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1049),
.A2(n_1065),
.B1(n_1061),
.B2(n_1167),
.Y(n_1248)
);

BUFx4f_ASAP7_75t_SL g1249 ( 
.A(n_1058),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_1066),
.Y(n_1250)
);

CKINVDCx11_ASAP7_75t_R g1251 ( 
.A(n_1167),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1132),
.Y(n_1252)
);

BUFx8_ASAP7_75t_L g1253 ( 
.A(n_1133),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1151),
.B(n_1172),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1050),
.A2(n_782),
.B1(n_926),
.B2(n_1149),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1107),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1121),
.Y(n_1257)
);

CKINVDCx6p67_ASAP7_75t_R g1258 ( 
.A(n_1073),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_1140),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1105),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1108),
.Y(n_1261)
);

OAI22xp33_ASAP7_75t_R g1262 ( 
.A1(n_1088),
.A2(n_323),
.B1(n_314),
.B2(n_683),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1149),
.A2(n_782),
.B1(n_926),
.B2(n_683),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1177),
.A2(n_683),
.B1(n_782),
.B2(n_926),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1105),
.Y(n_1265)
);

BUFx2_ASAP7_75t_SL g1266 ( 
.A(n_1108),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1177),
.A2(n_683),
.B1(n_782),
.B2(n_926),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1159),
.B(n_782),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1149),
.A2(n_782),
.B1(n_926),
.B2(n_683),
.Y(n_1269)
);

OAI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1159),
.A2(n_1131),
.B1(n_1179),
.B2(n_1148),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1159),
.A2(n_683),
.B1(n_942),
.B2(n_1153),
.Y(n_1271)
);

AO22x1_ASAP7_75t_L g1272 ( 
.A1(n_1079),
.A2(n_683),
.B1(n_506),
.B2(n_494),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1149),
.A2(n_782),
.B1(n_926),
.B2(n_683),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_SL g1274 ( 
.A1(n_1159),
.A2(n_683),
.B(n_474),
.Y(n_1274)
);

INVx8_ASAP7_75t_L g1275 ( 
.A(n_1121),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1105),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1148),
.B(n_683),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1105),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_1073),
.Y(n_1279)
);

INVx2_ASAP7_75t_SL g1280 ( 
.A(n_1095),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1149),
.A2(n_782),
.B1(n_926),
.B2(n_683),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1148),
.B(n_683),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1148),
.B(n_683),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1107),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1148),
.B(n_683),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_1171),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1121),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1095),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1140),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1159),
.A2(n_1131),
.B1(n_1179),
.B2(n_1148),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_SL g1291 ( 
.A1(n_1159),
.A2(n_683),
.B1(n_474),
.B2(n_953),
.Y(n_1291)
);

INVx1_ASAP7_75t_SL g1292 ( 
.A(n_1140),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_1121),
.Y(n_1293)
);

OR2x2_ASAP7_75t_L g1294 ( 
.A(n_1180),
.B(n_1237),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1195),
.B(n_1205),
.Y(n_1295)
);

AO21x2_ASAP7_75t_L g1296 ( 
.A1(n_1243),
.A2(n_1248),
.B(n_1244),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1236),
.B(n_1242),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1256),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1253),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1213),
.Y(n_1300)
);

BUFx2_ASAP7_75t_SL g1301 ( 
.A(n_1234),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1229),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1277),
.B(n_1282),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1229),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1246),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1236),
.B(n_1242),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_1240),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1246),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1253),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1247),
.B(n_1193),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1231),
.A2(n_1224),
.B(n_1252),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1193),
.B(n_1192),
.Y(n_1312)
);

INVxp67_ASAP7_75t_SL g1313 ( 
.A(n_1240),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1254),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1247),
.B(n_1196),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1256),
.B(n_1284),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1199),
.B(n_1270),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1227),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1188),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1249),
.A2(n_1273),
.B1(n_1269),
.B2(n_1263),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1190),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1249),
.A2(n_1273),
.B1(n_1269),
.B2(n_1263),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1197),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1250),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1284),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1231),
.A2(n_1224),
.B(n_1225),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1203),
.Y(n_1327)
);

AO21x2_ASAP7_75t_L g1328 ( 
.A1(n_1243),
.A2(n_1248),
.B(n_1241),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1196),
.B(n_1221),
.Y(n_1329)
);

AO21x2_ASAP7_75t_L g1330 ( 
.A1(n_1270),
.A2(n_1290),
.B(n_1183),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1210),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1271),
.A2(n_1281),
.B(n_1268),
.Y(n_1332)
);

OR2x6_ASAP7_75t_L g1333 ( 
.A(n_1223),
.B(n_1189),
.Y(n_1333)
);

OAI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1274),
.A2(n_1283),
.B1(n_1285),
.B2(n_1217),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1225),
.A2(n_1221),
.B(n_1255),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1262),
.A2(n_1291),
.B1(n_1281),
.B2(n_1182),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1238),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_1187),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1251),
.Y(n_1339)
);

INVxp67_ASAP7_75t_L g1340 ( 
.A(n_1260),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1255),
.A2(n_1202),
.B(n_1181),
.Y(n_1341)
);

INVx2_ASAP7_75t_SL g1342 ( 
.A(n_1239),
.Y(n_1342)
);

BUFx2_ASAP7_75t_SL g1343 ( 
.A(n_1228),
.Y(n_1343)
);

AO21x1_ASAP7_75t_SL g1344 ( 
.A1(n_1202),
.A2(n_1182),
.B(n_1267),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1199),
.B(n_1209),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1264),
.A2(n_1245),
.B(n_1191),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1265),
.Y(n_1347)
);

BUFx8_ASAP7_75t_L g1348 ( 
.A(n_1280),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1276),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1278),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1228),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1228),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1289),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1233),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1215),
.Y(n_1355)
);

O2A1O1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1290),
.A2(n_1204),
.B(n_1292),
.C(n_1259),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1209),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1201),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1208),
.B(n_1194),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1232),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1208),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1232),
.Y(n_1362)
);

INVxp67_ASAP7_75t_SL g1363 ( 
.A(n_1232),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1185),
.A2(n_1184),
.B(n_1207),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1218),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1212),
.B(n_1219),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1266),
.B(n_1216),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1272),
.B(n_1212),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1226),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1212),
.B(n_1261),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1184),
.B(n_1207),
.Y(n_1371)
);

AO31x2_ASAP7_75t_L g1372 ( 
.A1(n_1207),
.A2(n_1230),
.A3(n_1275),
.B(n_1206),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1222),
.Y(n_1373)
);

OR2x6_ASAP7_75t_L g1374 ( 
.A(n_1333),
.B(n_1275),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1336),
.A2(n_1235),
.B1(n_1220),
.B2(n_1258),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1355),
.B(n_1288),
.Y(n_1376)
);

OR2x6_ASAP7_75t_L g1377 ( 
.A(n_1333),
.B(n_1275),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1363),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1355),
.B(n_1286),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_SL g1380 ( 
.A1(n_1333),
.A2(n_1235),
.B1(n_1279),
.B2(n_1293),
.Y(n_1380)
);

A2O1A1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1332),
.A2(n_1186),
.B(n_1287),
.C(n_1257),
.Y(n_1381)
);

NAND4xp25_ASAP7_75t_L g1382 ( 
.A(n_1303),
.B(n_1198),
.C(n_1222),
.D(n_1206),
.Y(n_1382)
);

AND2x2_ASAP7_75t_SL g1383 ( 
.A(n_1329),
.B(n_1186),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1359),
.B(n_1200),
.Y(n_1384)
);

NOR2x1_ASAP7_75t_L g1385 ( 
.A(n_1368),
.B(n_1257),
.Y(n_1385)
);

A2O1A1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_1332),
.A2(n_1356),
.B(n_1317),
.C(n_1329),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1359),
.B(n_1293),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1333),
.A2(n_1211),
.B(n_1235),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1319),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1333),
.A2(n_1287),
.B(n_1293),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1319),
.Y(n_1391)
);

OA21x2_ASAP7_75t_L g1392 ( 
.A1(n_1341),
.A2(n_1214),
.B(n_1326),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1333),
.A2(n_1337),
.B(n_1320),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1302),
.B(n_1304),
.Y(n_1394)
);

AOI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1320),
.A2(n_1322),
.B1(n_1334),
.B2(n_1312),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1339),
.B(n_1307),
.Y(n_1396)
);

A2O1A1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1356),
.A2(n_1317),
.B(n_1329),
.C(n_1337),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1321),
.Y(n_1398)
);

A2O1A1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1295),
.A2(n_1312),
.B(n_1324),
.C(n_1322),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1339),
.B(n_1307),
.Y(n_1400)
);

A2O1A1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1295),
.A2(n_1324),
.B(n_1345),
.C(n_1341),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1302),
.B(n_1304),
.Y(n_1402)
);

CKINVDCx16_ASAP7_75t_R g1403 ( 
.A(n_1301),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1316),
.B(n_1298),
.Y(n_1404)
);

AO32x2_ASAP7_75t_L g1405 ( 
.A1(n_1342),
.A2(n_1351),
.A3(n_1352),
.B1(n_1306),
.B2(n_1297),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1370),
.B(n_1301),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1323),
.B(n_1327),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1313),
.A2(n_1315),
.B1(n_1345),
.B2(n_1310),
.Y(n_1408)
);

O2A1O1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1330),
.A2(n_1368),
.B(n_1308),
.C(n_1305),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1366),
.B(n_1325),
.Y(n_1410)
);

AO32x2_ASAP7_75t_L g1411 ( 
.A1(n_1342),
.A2(n_1352),
.A3(n_1351),
.B1(n_1306),
.B2(n_1297),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1325),
.B(n_1360),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1360),
.B(n_1363),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1341),
.A2(n_1326),
.B(n_1311),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1358),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_SL g1416 ( 
.A(n_1299),
.B(n_1309),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1353),
.B(n_1318),
.Y(n_1417)
);

AOI221xp5_ASAP7_75t_L g1418 ( 
.A1(n_1315),
.A2(n_1357),
.B1(n_1361),
.B2(n_1310),
.C(n_1297),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1358),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1370),
.B(n_1367),
.Y(n_1420)
);

AOI221xp5_ASAP7_75t_L g1421 ( 
.A1(n_1357),
.A2(n_1361),
.B1(n_1306),
.B2(n_1330),
.C(n_1340),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_SL g1422 ( 
.A1(n_1373),
.A2(n_1338),
.B(n_1371),
.C(n_1299),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1360),
.B(n_1316),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1347),
.B(n_1349),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1331),
.B(n_1362),
.Y(n_1425)
);

AO21x1_ASAP7_75t_L g1426 ( 
.A1(n_1349),
.A2(n_1350),
.B(n_1369),
.Y(n_1426)
);

CKINVDCx20_ASAP7_75t_R g1427 ( 
.A(n_1348),
.Y(n_1427)
);

A2O1A1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1346),
.A2(n_1335),
.B(n_1326),
.C(n_1300),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1414),
.B(n_1405),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1405),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1395),
.A2(n_1330),
.B1(n_1331),
.B2(n_1296),
.Y(n_1431)
);

AND2x4_ASAP7_75t_SL g1432 ( 
.A(n_1374),
.B(n_1299),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1405),
.B(n_1328),
.Y(n_1433)
);

NOR2x1_ASAP7_75t_SL g1434 ( 
.A(n_1374),
.B(n_1328),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_SL g1435 ( 
.A1(n_1393),
.A2(n_1330),
.B1(n_1300),
.B2(n_1328),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1389),
.Y(n_1436)
);

INVxp67_ASAP7_75t_SL g1437 ( 
.A(n_1426),
.Y(n_1437)
);

INVxp67_ASAP7_75t_L g1438 ( 
.A(n_1378),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1391),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1395),
.A2(n_1344),
.B1(n_1296),
.B2(n_1335),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1398),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1411),
.B(n_1296),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1428),
.B(n_1296),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1411),
.B(n_1314),
.Y(n_1444)
);

INVx3_ASAP7_75t_L g1445 ( 
.A(n_1404),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1411),
.B(n_1314),
.Y(n_1446)
);

CKINVDCx16_ASAP7_75t_R g1447 ( 
.A(n_1403),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1392),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1407),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1417),
.B(n_1294),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1393),
.A2(n_1344),
.B1(n_1335),
.B2(n_1346),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1424),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1394),
.B(n_1294),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1402),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1430),
.B(n_1396),
.Y(n_1455)
);

OAI31xp33_ASAP7_75t_SL g1456 ( 
.A1(n_1435),
.A2(n_1421),
.A3(n_1408),
.B(n_1418),
.Y(n_1456)
);

NAND2x1_ASAP7_75t_L g1457 ( 
.A(n_1430),
.B(n_1377),
.Y(n_1457)
);

OAI31xp33_ASAP7_75t_L g1458 ( 
.A1(n_1440),
.A2(n_1386),
.A3(n_1399),
.B(n_1401),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1444),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1444),
.Y(n_1460)
);

INVx1_ASAP7_75t_SL g1461 ( 
.A(n_1450),
.Y(n_1461)
);

OAI221xp5_ASAP7_75t_L g1462 ( 
.A1(n_1435),
.A2(n_1375),
.B1(n_1397),
.B2(n_1388),
.C(n_1380),
.Y(n_1462)
);

OR2x6_ASAP7_75t_SL g1463 ( 
.A(n_1443),
.B(n_1408),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1436),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1444),
.Y(n_1465)
);

INVx4_ASAP7_75t_L g1466 ( 
.A(n_1432),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1447),
.B(n_1382),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1446),
.Y(n_1468)
);

OAI221xp5_ASAP7_75t_L g1469 ( 
.A1(n_1440),
.A2(n_1375),
.B1(n_1388),
.B2(n_1409),
.C(n_1381),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1452),
.B(n_1412),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1451),
.A2(n_1431),
.B1(n_1383),
.B2(n_1377),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1436),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1429),
.B(n_1423),
.Y(n_1473)
);

OAI221xp5_ASAP7_75t_L g1474 ( 
.A1(n_1431),
.A2(n_1390),
.B1(n_1382),
.B2(n_1416),
.C(n_1384),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1432),
.Y(n_1475)
);

OAI21xp33_ASAP7_75t_SL g1476 ( 
.A1(n_1437),
.A2(n_1390),
.B(n_1364),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_SL g1477 ( 
.A(n_1447),
.B(n_1416),
.Y(n_1477)
);

AOI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1451),
.A2(n_1387),
.B1(n_1420),
.B2(n_1346),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1439),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1439),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1430),
.B(n_1415),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1441),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1452),
.B(n_1425),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1446),
.B(n_1400),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1454),
.B(n_1413),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1454),
.B(n_1419),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1450),
.B(n_1410),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1429),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1429),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1432),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1464),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1483),
.B(n_1470),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1464),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1472),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1459),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1461),
.B(n_1454),
.Y(n_1496)
);

NOR3xp33_ASAP7_75t_SL g1497 ( 
.A(n_1474),
.B(n_1406),
.C(n_1373),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1481),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1472),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1461),
.B(n_1454),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1481),
.B(n_1450),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1455),
.Y(n_1502)
);

INVxp67_ASAP7_75t_SL g1503 ( 
.A(n_1486),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1459),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1463),
.Y(n_1505)
);

INVx6_ASAP7_75t_L g1506 ( 
.A(n_1466),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1483),
.B(n_1438),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1489),
.B(n_1437),
.Y(n_1508)
);

BUFx2_ASAP7_75t_L g1509 ( 
.A(n_1463),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1470),
.B(n_1438),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1479),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1486),
.B(n_1449),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1479),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1473),
.B(n_1445),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1473),
.B(n_1445),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1467),
.B(n_1379),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1475),
.B(n_1434),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1459),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1474),
.B(n_1376),
.Y(n_1519)
);

INVx1_ASAP7_75t_SL g1520 ( 
.A(n_1463),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1480),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1455),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1480),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1460),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1482),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1489),
.B(n_1453),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_R g1527 ( 
.A(n_1477),
.B(n_1427),
.Y(n_1527)
);

INVxp67_ASAP7_75t_SL g1528 ( 
.A(n_1485),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1519),
.B(n_1456),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1503),
.B(n_1456),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1495),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1509),
.B(n_1488),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1509),
.B(n_1488),
.Y(n_1533)
);

NAND2x1p5_ASAP7_75t_L g1534 ( 
.A(n_1505),
.B(n_1466),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1498),
.B(n_1489),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1527),
.Y(n_1536)
);

CKINVDCx16_ASAP7_75t_R g1537 ( 
.A(n_1505),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1501),
.B(n_1487),
.Y(n_1538)
);

INVx2_ASAP7_75t_SL g1539 ( 
.A(n_1506),
.Y(n_1539)
);

AOI211xp5_ASAP7_75t_L g1540 ( 
.A1(n_1520),
.A2(n_1462),
.B(n_1469),
.C(n_1458),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1495),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1501),
.B(n_1487),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1502),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1492),
.B(n_1458),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1491),
.Y(n_1545)
);

INVxp67_ASAP7_75t_L g1546 ( 
.A(n_1516),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1491),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1493),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1493),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1494),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1494),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1499),
.Y(n_1552)
);

AND2x4_ASAP7_75t_SL g1553 ( 
.A(n_1497),
.B(n_1466),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1499),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1520),
.B(n_1460),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1508),
.B(n_1460),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1495),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1511),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1508),
.B(n_1465),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1511),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1513),
.Y(n_1561)
);

O2A1O1Ixp33_ASAP7_75t_L g1562 ( 
.A1(n_1507),
.A2(n_1462),
.B(n_1469),
.C(n_1443),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1528),
.B(n_1484),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1504),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1526),
.B(n_1465),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1526),
.B(n_1465),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1513),
.Y(n_1567)
);

AO22x1_ASAP7_75t_L g1568 ( 
.A1(n_1517),
.A2(n_1385),
.B1(n_1490),
.B2(n_1475),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1522),
.B(n_1468),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1517),
.B(n_1475),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_1537),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1538),
.B(n_1512),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1532),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1540),
.B(n_1536),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1545),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1532),
.B(n_1517),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1533),
.B(n_1517),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1538),
.B(n_1510),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1542),
.B(n_1504),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1533),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1547),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1534),
.B(n_1570),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1529),
.B(n_1484),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1542),
.B(n_1504),
.Y(n_1584)
);

INVxp67_ASAP7_75t_L g1585 ( 
.A(n_1543),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1535),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1548),
.Y(n_1587)
);

INVx3_ASAP7_75t_L g1588 ( 
.A(n_1534),
.Y(n_1588)
);

NAND2x1_ASAP7_75t_L g1589 ( 
.A(n_1570),
.B(n_1506),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1535),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1570),
.B(n_1506),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1549),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1550),
.Y(n_1593)
);

AND3x2_ASAP7_75t_L g1594 ( 
.A(n_1546),
.B(n_1477),
.C(n_1448),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1530),
.A2(n_1476),
.B(n_1457),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1551),
.Y(n_1596)
);

OAI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1562),
.A2(n_1478),
.B(n_1476),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1539),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1563),
.B(n_1518),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1552),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1555),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1554),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1558),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1555),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1560),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1571),
.A2(n_1553),
.B1(n_1544),
.B2(n_1478),
.Y(n_1606)
);

A2O1A1Ixp33_ASAP7_75t_L g1607 ( 
.A1(n_1597),
.A2(n_1553),
.B(n_1443),
.C(n_1457),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1573),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1571),
.B(n_1539),
.Y(n_1609)
);

NAND2x1p5_ASAP7_75t_L g1610 ( 
.A(n_1588),
.B(n_1309),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1597),
.A2(n_1471),
.B1(n_1506),
.B2(n_1448),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1575),
.Y(n_1612)
);

OAI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1574),
.A2(n_1506),
.B1(n_1448),
.B2(n_1569),
.C(n_1561),
.Y(n_1613)
);

AOI211xp5_ASAP7_75t_L g1614 ( 
.A1(n_1595),
.A2(n_1585),
.B(n_1582),
.C(n_1588),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1582),
.B(n_1514),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1591),
.Y(n_1616)
);

INVxp67_ASAP7_75t_L g1617 ( 
.A(n_1598),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1598),
.B(n_1567),
.Y(n_1618)
);

AOI221x1_ASAP7_75t_L g1619 ( 
.A1(n_1588),
.A2(n_1557),
.B1(n_1531),
.B2(n_1564),
.C(n_1541),
.Y(n_1619)
);

OAI31xp33_ASAP7_75t_L g1620 ( 
.A1(n_1588),
.A2(n_1569),
.A3(n_1559),
.B(n_1556),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1583),
.B(n_1568),
.Y(n_1621)
);

A2O1A1Ixp33_ASAP7_75t_L g1622 ( 
.A1(n_1589),
.A2(n_1433),
.B(n_1442),
.C(n_1309),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1576),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1578),
.B(n_1565),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1580),
.B(n_1578),
.Y(n_1625)
);

INVxp67_ASAP7_75t_SL g1626 ( 
.A(n_1580),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1580),
.B(n_1490),
.Y(n_1627)
);

AO22x1_ASAP7_75t_L g1628 ( 
.A1(n_1591),
.A2(n_1348),
.B1(n_1490),
.B2(n_1466),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1575),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1601),
.B(n_1514),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1626),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1606),
.A2(n_1589),
.B1(n_1601),
.B2(n_1604),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1626),
.B(n_1601),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1608),
.Y(n_1634)
);

O2A1O1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1611),
.A2(n_1605),
.B(n_1592),
.C(n_1596),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1618),
.Y(n_1636)
);

XOR2xp5_ASAP7_75t_L g1637 ( 
.A(n_1609),
.B(n_1367),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1618),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1616),
.B(n_1604),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1617),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1610),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1615),
.B(n_1576),
.Y(n_1642)
);

NAND2x1p5_ASAP7_75t_L g1643 ( 
.A(n_1627),
.B(n_1612),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1624),
.B(n_1604),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1629),
.Y(n_1645)
);

OAI21xp33_ASAP7_75t_SL g1646 ( 
.A1(n_1620),
.A2(n_1577),
.B(n_1586),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1617),
.B(n_1586),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1610),
.Y(n_1648)
);

NAND3xp33_ASAP7_75t_L g1649 ( 
.A(n_1614),
.B(n_1594),
.C(n_1587),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1640),
.B(n_1636),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1636),
.B(n_1623),
.Y(n_1651)
);

XNOR2x2_ASAP7_75t_L g1652 ( 
.A(n_1649),
.B(n_1613),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1637),
.A2(n_1607),
.B1(n_1621),
.B2(n_1625),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1633),
.Y(n_1654)
);

O2A1O1Ixp33_ASAP7_75t_L g1655 ( 
.A1(n_1632),
.A2(n_1622),
.B(n_1625),
.C(n_1602),
.Y(n_1655)
);

AOI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1635),
.A2(n_1622),
.B1(n_1630),
.B2(n_1586),
.C(n_1590),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1637),
.B(n_1627),
.Y(n_1657)
);

INVxp67_ASAP7_75t_L g1658 ( 
.A(n_1638),
.Y(n_1658)
);

OAI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1638),
.A2(n_1577),
.B1(n_1572),
.B2(n_1590),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1638),
.B(n_1590),
.Y(n_1660)
);

NOR4xp25_ASAP7_75t_L g1661 ( 
.A(n_1658),
.B(n_1634),
.C(n_1631),
.D(n_1645),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1657),
.B(n_1650),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1654),
.B(n_1634),
.Y(n_1663)
);

INVxp67_ASAP7_75t_SL g1664 ( 
.A(n_1660),
.Y(n_1664)
);

OAI21xp5_ASAP7_75t_SL g1665 ( 
.A1(n_1655),
.A2(n_1643),
.B(n_1639),
.Y(n_1665)
);

AOI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1653),
.A2(n_1646),
.B1(n_1647),
.B2(n_1643),
.C(n_1633),
.Y(n_1666)
);

NAND3xp33_ASAP7_75t_L g1667 ( 
.A(n_1656),
.B(n_1633),
.C(n_1644),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1651),
.Y(n_1668)
);

NAND3xp33_ASAP7_75t_L g1669 ( 
.A(n_1659),
.B(n_1644),
.C(n_1641),
.Y(n_1669)
);

AOI211xp5_ASAP7_75t_L g1670 ( 
.A1(n_1652),
.A2(n_1628),
.B(n_1642),
.C(n_1641),
.Y(n_1670)
);

AOI211xp5_ASAP7_75t_L g1671 ( 
.A1(n_1665),
.A2(n_1642),
.B(n_1648),
.C(n_1602),
.Y(n_1671)
);

OAI211xp5_ASAP7_75t_L g1672 ( 
.A1(n_1666),
.A2(n_1619),
.B(n_1648),
.C(n_1643),
.Y(n_1672)
);

NAND4xp25_ASAP7_75t_L g1673 ( 
.A(n_1670),
.B(n_1605),
.C(n_1603),
.D(n_1600),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1667),
.A2(n_1572),
.B1(n_1599),
.B2(n_1600),
.Y(n_1674)
);

NAND3xp33_ASAP7_75t_L g1675 ( 
.A(n_1669),
.B(n_1662),
.C(n_1661),
.Y(n_1675)
);

NAND4xp25_ASAP7_75t_L g1676 ( 
.A(n_1668),
.B(n_1603),
.C(n_1581),
.D(n_1596),
.Y(n_1676)
);

AOI211xp5_ASAP7_75t_L g1677 ( 
.A1(n_1664),
.A2(n_1593),
.B(n_1581),
.C(n_1587),
.Y(n_1677)
);

O2A1O1Ixp33_ASAP7_75t_L g1678 ( 
.A1(n_1675),
.A2(n_1663),
.B(n_1592),
.C(n_1593),
.Y(n_1678)
);

OAI31xp33_ASAP7_75t_L g1679 ( 
.A1(n_1672),
.A2(n_1599),
.A3(n_1584),
.B(n_1579),
.Y(n_1679)
);

NOR3xp33_ASAP7_75t_SL g1680 ( 
.A(n_1673),
.B(n_1371),
.C(n_1348),
.Y(n_1680)
);

AOI211xp5_ASAP7_75t_L g1681 ( 
.A1(n_1674),
.A2(n_1584),
.B(n_1579),
.C(n_1353),
.Y(n_1681)
);

AOI221x1_ASAP7_75t_L g1682 ( 
.A1(n_1676),
.A2(n_1531),
.B1(n_1564),
.B2(n_1541),
.C(n_1557),
.Y(n_1682)
);

OAI31xp33_ASAP7_75t_L g1683 ( 
.A1(n_1671),
.A2(n_1559),
.A3(n_1556),
.B(n_1566),
.Y(n_1683)
);

OAI211xp5_ASAP7_75t_SL g1684 ( 
.A1(n_1677),
.A2(n_1566),
.B(n_1565),
.C(n_1354),
.Y(n_1684)
);

XNOR2x1_ASAP7_75t_L g1685 ( 
.A(n_1679),
.B(n_1348),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1680),
.B(n_1515),
.Y(n_1686)
);

NOR2x1_ASAP7_75t_L g1687 ( 
.A(n_1678),
.B(n_1521),
.Y(n_1687)
);

NOR2x1_ASAP7_75t_L g1688 ( 
.A(n_1684),
.B(n_1521),
.Y(n_1688)
);

NOR2x1_ASAP7_75t_L g1689 ( 
.A(n_1681),
.B(n_1523),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1685),
.B(n_1683),
.Y(n_1690)
);

AOI22x1_ASAP7_75t_L g1691 ( 
.A1(n_1686),
.A2(n_1682),
.B1(n_1343),
.B2(n_1524),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1689),
.B(n_1496),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1690),
.B(n_1687),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1693),
.Y(n_1694)
);

XNOR2xp5_ASAP7_75t_L g1695 ( 
.A(n_1694),
.B(n_1691),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1694),
.A2(n_1692),
.B1(n_1688),
.B2(n_1518),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1695),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1696),
.A2(n_1524),
.B1(n_1518),
.B2(n_1525),
.Y(n_1698)
);

NAND3xp33_ASAP7_75t_L g1699 ( 
.A(n_1697),
.B(n_1525),
.C(n_1523),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1698),
.Y(n_1700)
);

OAI21x1_ASAP7_75t_L g1701 ( 
.A1(n_1700),
.A2(n_1524),
.B(n_1500),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1701),
.A2(n_1699),
.B(n_1422),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1702),
.Y(n_1703)
);

OAI221xp5_ASAP7_75t_R g1704 ( 
.A1(n_1703),
.A2(n_1372),
.B1(n_1434),
.B2(n_1496),
.C(n_1500),
.Y(n_1704)
);

AOI211xp5_ASAP7_75t_L g1705 ( 
.A1(n_1704),
.A2(n_1354),
.B(n_1365),
.C(n_1369),
.Y(n_1705)
);


endmodule