module real_aes_6501_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_0), .B(n_105), .C(n_106), .Y(n_104) );
INVx1_ASAP7_75t_L g123 ( .A(n_0), .Y(n_123) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_1), .A2(n_155), .B(n_158), .C(n_238), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_2), .A2(n_184), .B(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g484 ( .A(n_3), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_4), .B(n_214), .Y(n_213) );
AOI21xp33_ASAP7_75t_L g467 ( .A1(n_5), .A2(n_184), .B(n_468), .Y(n_467) );
AND2x6_ASAP7_75t_L g155 ( .A(n_6), .B(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g251 ( .A(n_7), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_8), .B(n_41), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_9), .A2(n_183), .B(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_10), .B(n_167), .Y(n_240) );
INVx1_ASAP7_75t_L g472 ( .A(n_11), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_12), .B(n_208), .Y(n_507) );
INVx1_ASAP7_75t_L g147 ( .A(n_13), .Y(n_147) );
INVx1_ASAP7_75t_L g519 ( .A(n_14), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_15), .A2(n_78), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_15), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_16), .A2(n_192), .B(n_273), .C(n_275), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_17), .B(n_214), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_18), .B(n_450), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_19), .B(n_184), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_20), .B(n_198), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_21), .A2(n_208), .B(n_259), .C(n_261), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_22), .B(n_214), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_23), .B(n_167), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_24), .A2(n_194), .B(n_275), .C(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_25), .B(n_167), .Y(n_222) );
CKINVDCx16_ASAP7_75t_R g149 ( .A(n_26), .Y(n_149) );
INVx1_ASAP7_75t_L g221 ( .A(n_27), .Y(n_221) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_28), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_29), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_30), .B(n_167), .Y(n_485) );
INVx1_ASAP7_75t_L g190 ( .A(n_31), .Y(n_190) );
INVx1_ASAP7_75t_L g462 ( .A(n_32), .Y(n_462) );
INVx2_ASAP7_75t_L g153 ( .A(n_33), .Y(n_153) );
AOI222xp33_ASAP7_75t_SL g125 ( .A1(n_34), .A2(n_126), .B1(n_129), .B2(n_722), .C1(n_723), .C2(n_725), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_35), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_36), .A2(n_208), .B(n_209), .C(n_211), .Y(n_207) );
INVxp67_ASAP7_75t_L g193 ( .A(n_37), .Y(n_193) );
CKINVDCx14_ASAP7_75t_R g206 ( .A(n_38), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_39), .A2(n_158), .B(n_220), .C(n_224), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_40), .A2(n_155), .B(n_158), .C(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g461 ( .A(n_42), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_43), .A2(n_169), .B(n_249), .C(n_250), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_44), .B(n_167), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_45), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_46), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_47), .A2(n_102), .B1(n_111), .B2(n_738), .Y(n_101) );
INVx1_ASAP7_75t_L g257 ( .A(n_48), .Y(n_257) );
CKINVDCx16_ASAP7_75t_R g463 ( .A(n_49), .Y(n_463) );
OAI22xp5_ASAP7_75t_SL g733 ( .A1(n_50), .A2(n_60), .B1(n_734), .B2(n_735), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_50), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_51), .B(n_184), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_52), .A2(n_158), .B1(n_261), .B2(n_460), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_53), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g481 ( .A(n_54), .Y(n_481) );
CKINVDCx14_ASAP7_75t_R g247 ( .A(n_55), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_56), .A2(n_211), .B(n_249), .C(n_471), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_57), .Y(n_124) );
INVx1_ASAP7_75t_L g469 ( .A(n_58), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_59), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_60), .Y(n_735) );
INVx1_ASAP7_75t_L g156 ( .A(n_61), .Y(n_156) );
INVx1_ASAP7_75t_L g146 ( .A(n_62), .Y(n_146) );
INVx1_ASAP7_75t_SL g210 ( .A(n_63), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_64), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_65), .B(n_214), .Y(n_263) );
INVx1_ASAP7_75t_L g162 ( .A(n_66), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_SL g449 ( .A1(n_67), .A2(n_211), .B(n_450), .C(n_451), .Y(n_449) );
INVxp67_ASAP7_75t_L g452 ( .A(n_68), .Y(n_452) );
INVx1_ASAP7_75t_L g108 ( .A(n_69), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_70), .A2(n_184), .B(n_246), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_71), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_72), .A2(n_184), .B(n_270), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_73), .Y(n_465) );
INVx1_ASAP7_75t_L g525 ( .A(n_74), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_75), .A2(n_183), .B(n_185), .Y(n_182) );
CKINVDCx16_ASAP7_75t_R g218 ( .A(n_76), .Y(n_218) );
INVx1_ASAP7_75t_L g271 ( .A(n_77), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_78), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_79), .A2(n_155), .B(n_158), .C(n_527), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_80), .A2(n_184), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g274 ( .A(n_81), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_82), .B(n_191), .Y(n_496) );
INVx2_ASAP7_75t_L g144 ( .A(n_83), .Y(n_144) );
INVx1_ASAP7_75t_L g239 ( .A(n_84), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_85), .B(n_450), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_86), .A2(n_155), .B(n_158), .C(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g105 ( .A(n_87), .Y(n_105) );
OR2x2_ASAP7_75t_L g120 ( .A(n_87), .B(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g437 ( .A(n_87), .B(n_122), .Y(n_437) );
A2O1A1Ixp33_ASAP7_75t_L g157 ( .A1(n_88), .A2(n_158), .B(n_161), .C(n_171), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_89), .B(n_176), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_90), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_91), .A2(n_155), .B(n_158), .C(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_92), .Y(n_511) );
INVx1_ASAP7_75t_L g448 ( .A(n_93), .Y(n_448) );
CKINVDCx16_ASAP7_75t_R g516 ( .A(n_94), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_95), .B(n_191), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_96), .B(n_142), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_97), .B(n_142), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_98), .B(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g260 ( .A(n_99), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_100), .A2(n_184), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_103), .Y(n_739) );
OR2x2_ASAP7_75t_SL g103 ( .A(n_104), .B(n_109), .Y(n_103) );
OR2x2_ASAP7_75t_L g721 ( .A(n_105), .B(n_122), .Y(n_721) );
NOR2x2_ASAP7_75t_L g727 ( .A(n_105), .B(n_121), .Y(n_727) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g122 ( .A(n_110), .B(n_123), .Y(n_122) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AOI22xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_125), .B1(n_728), .B2(n_730), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_117), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g729 ( .A(n_115), .Y(n_729) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_117), .A2(n_731), .B(n_736), .Y(n_730) );
NOR2xp33_ASAP7_75t_SL g117 ( .A(n_118), .B(n_124), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g737 ( .A(n_120), .Y(n_737) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g722 ( .A(n_126), .Y(n_722) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_437), .B1(n_438), .B2(n_719), .Y(n_129) );
OAI22xp5_ASAP7_75t_SL g731 ( .A1(n_130), .A2(n_131), .B1(n_732), .B2(n_733), .Y(n_731) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g723 ( .A1(n_131), .A2(n_437), .B1(n_719), .B2(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_371), .Y(n_131) );
NAND5xp2_ASAP7_75t_L g132 ( .A(n_133), .B(n_300), .C(n_330), .D(n_351), .E(n_357), .Y(n_132) );
AOI221xp5_ASAP7_75t_SL g133 ( .A1(n_134), .A2(n_230), .B1(n_264), .B2(n_266), .C(n_277), .Y(n_133) );
INVxp67_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_227), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_199), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_SL g351 ( .A1(n_138), .A2(n_215), .B(n_352), .C(n_355), .Y(n_351) );
AND2x2_ASAP7_75t_L g421 ( .A(n_138), .B(n_216), .Y(n_421) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_177), .Y(n_138) );
AND2x2_ASAP7_75t_L g279 ( .A(n_139), .B(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g283 ( .A(n_139), .B(n_280), .Y(n_283) );
OR2x2_ASAP7_75t_L g309 ( .A(n_139), .B(n_216), .Y(n_309) );
AND2x2_ASAP7_75t_L g311 ( .A(n_139), .B(n_202), .Y(n_311) );
AND2x2_ASAP7_75t_L g329 ( .A(n_139), .B(n_201), .Y(n_329) );
INVx1_ASAP7_75t_L g362 ( .A(n_139), .Y(n_362) );
INVx2_ASAP7_75t_SL g139 ( .A(n_140), .Y(n_139) );
BUFx2_ASAP7_75t_L g229 ( .A(n_140), .Y(n_229) );
AND2x2_ASAP7_75t_L g265 ( .A(n_140), .B(n_202), .Y(n_265) );
AND2x2_ASAP7_75t_L g418 ( .A(n_140), .B(n_216), .Y(n_418) );
AO21x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_148), .B(n_173), .Y(n_140) );
INVx3_ASAP7_75t_L g214 ( .A(n_141), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_141), .B(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_141), .B(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_SL g498 ( .A(n_141), .B(n_499), .Y(n_498) );
INVx4_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_142), .Y(n_203) );
OA21x2_ASAP7_75t_L g445 ( .A1(n_142), .A2(n_446), .B(n_453), .Y(n_445) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g180 ( .A(n_143), .Y(n_180) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AND2x2_ASAP7_75t_SL g176 ( .A(n_144), .B(n_145), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
OAI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_157), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_150), .A2(n_176), .B(n_218), .C(n_219), .Y(n_217) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_150), .A2(n_236), .B(n_237), .Y(n_235) );
OAI22xp33_ASAP7_75t_L g458 ( .A1(n_150), .A2(n_172), .B1(n_459), .B2(n_463), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_150), .A2(n_481), .B(n_482), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_150), .A2(n_525), .B(n_526), .Y(n_524) );
NAND2x1p5_ASAP7_75t_L g150 ( .A(n_151), .B(n_155), .Y(n_150) );
AND2x4_ASAP7_75t_L g184 ( .A(n_151), .B(n_155), .Y(n_184) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_154), .Y(n_151) );
INVx1_ASAP7_75t_L g195 ( .A(n_152), .Y(n_195) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g159 ( .A(n_153), .Y(n_159) );
INVx1_ASAP7_75t_L g262 ( .A(n_153), .Y(n_262) );
INVx1_ASAP7_75t_L g160 ( .A(n_154), .Y(n_160) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_154), .Y(n_165) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_154), .Y(n_167) );
INVx3_ASAP7_75t_L g192 ( .A(n_154), .Y(n_192) );
INVx1_ASAP7_75t_L g450 ( .A(n_154), .Y(n_450) );
INVx4_ASAP7_75t_SL g172 ( .A(n_155), .Y(n_172) );
BUFx3_ASAP7_75t_L g224 ( .A(n_155), .Y(n_224) );
INVx5_ASAP7_75t_L g187 ( .A(n_158), .Y(n_187) );
AND2x6_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
BUFx3_ASAP7_75t_L g170 ( .A(n_159), .Y(n_170) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_159), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_166), .C(n_168), .Y(n_161) );
O2A1O1Ixp5_ASAP7_75t_L g238 ( .A1(n_163), .A2(n_168), .B(n_239), .C(n_240), .Y(n_238) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
OAI22xp5_ASAP7_75t_SL g460 ( .A1(n_164), .A2(n_165), .B1(n_461), .B2(n_462), .Y(n_460) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx4_ASAP7_75t_L g194 ( .A(n_165), .Y(n_194) );
INVx4_ASAP7_75t_L g208 ( .A(n_167), .Y(n_208) );
INVx2_ASAP7_75t_L g249 ( .A(n_167), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_168), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_168), .A2(n_528), .B(n_529), .Y(n_527) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g275 ( .A(n_170), .Y(n_275) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_SL g185 ( .A1(n_172), .A2(n_186), .B(n_187), .C(n_188), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g205 ( .A1(n_172), .A2(n_187), .B(n_206), .C(n_207), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_SL g246 ( .A1(n_172), .A2(n_187), .B(n_247), .C(n_248), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_SL g256 ( .A1(n_172), .A2(n_187), .B(n_257), .C(n_258), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_SL g270 ( .A1(n_172), .A2(n_187), .B(n_271), .C(n_272), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g447 ( .A1(n_172), .A2(n_187), .B(n_448), .C(n_449), .Y(n_447) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_172), .A2(n_187), .B(n_469), .C(n_470), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_172), .A2(n_187), .B(n_516), .C(n_517), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
INVx1_ASAP7_75t_L g198 ( .A(n_175), .Y(n_198) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_175), .A2(n_503), .B(n_510), .Y(n_502) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g234 ( .A(n_176), .Y(n_234) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_176), .A2(n_245), .B(n_252), .Y(n_244) );
OA21x2_ASAP7_75t_L g513 ( .A1(n_176), .A2(n_514), .B(n_520), .Y(n_513) );
AND2x2_ASAP7_75t_L g299 ( .A(n_177), .B(n_200), .Y(n_299) );
OR2x2_ASAP7_75t_L g303 ( .A(n_177), .B(n_216), .Y(n_303) );
AND2x2_ASAP7_75t_L g328 ( .A(n_177), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g375 ( .A(n_177), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_177), .B(n_337), .Y(n_423) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_181), .B(n_196), .Y(n_177) );
INVx1_ASAP7_75t_L g281 ( .A(n_178), .Y(n_281) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_178), .A2(n_524), .B(n_530), .Y(n_523) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AOI21xp5_ASAP7_75t_SL g492 ( .A1(n_179), .A2(n_493), .B(n_494), .Y(n_492) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_180), .A2(n_458), .B(n_464), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_180), .B(n_465), .Y(n_464) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_180), .A2(n_480), .B(n_487), .Y(n_479) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
OA21x2_ASAP7_75t_L g280 ( .A1(n_182), .A2(n_197), .B(n_281), .Y(n_280) );
BUFx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_189), .B(n_195), .Y(n_188) );
OAI22xp33_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B1(n_193), .B2(n_194), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_191), .A2(n_221), .B(n_222), .C(n_223), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_191), .A2(n_484), .B(n_485), .C(n_486), .Y(n_483) );
INVx5_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_192), .B(n_251), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_192), .B(n_452), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_192), .B(n_472), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_194), .B(n_260), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_194), .B(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_194), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g223 ( .A(n_195), .Y(n_223) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OAI322xp33_ASAP7_75t_L g424 ( .A1(n_199), .A2(n_360), .A3(n_383), .B1(n_404), .B2(n_425), .C1(n_427), .C2(n_428), .Y(n_424) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_200), .B(n_280), .Y(n_427) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_215), .Y(n_200) );
AND2x2_ASAP7_75t_L g228 ( .A(n_201), .B(n_229), .Y(n_228) );
AND2x4_ASAP7_75t_L g296 ( .A(n_201), .B(n_216), .Y(n_296) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g337 ( .A(n_202), .B(n_216), .Y(n_337) );
AND2x2_ASAP7_75t_L g381 ( .A(n_202), .B(n_215), .Y(n_381) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_213), .Y(n_202) );
OA21x2_ASAP7_75t_L g254 ( .A1(n_203), .A2(n_255), .B(n_263), .Y(n_254) );
OA21x2_ASAP7_75t_L g268 ( .A1(n_203), .A2(n_269), .B(n_276), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_208), .B(n_210), .Y(n_209) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_212), .Y(n_508) );
OA21x2_ASAP7_75t_L g466 ( .A1(n_214), .A2(n_467), .B(n_473), .Y(n_466) );
AND2x2_ASAP7_75t_L g264 ( .A(n_215), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g282 ( .A(n_215), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_215), .B(n_311), .Y(n_435) );
INVx3_ASAP7_75t_SL g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g227 ( .A(n_216), .B(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_216), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g349 ( .A(n_216), .B(n_280), .Y(n_349) );
AND2x2_ASAP7_75t_L g376 ( .A(n_216), .B(n_311), .Y(n_376) );
OR2x2_ASAP7_75t_L g432 ( .A(n_216), .B(n_283), .Y(n_432) );
OR2x6_ASAP7_75t_L g216 ( .A(n_217), .B(n_225), .Y(n_216) );
INVx1_ASAP7_75t_SL g318 ( .A(n_227), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_228), .B(n_349), .Y(n_350) );
AND2x2_ASAP7_75t_L g384 ( .A(n_228), .B(n_374), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_228), .B(n_307), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_228), .B(n_429), .Y(n_428) );
OAI31xp33_ASAP7_75t_L g402 ( .A1(n_230), .A2(n_264), .A3(n_403), .B(n_405), .Y(n_402) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_243), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_231), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g385 ( .A(n_231), .B(n_320), .Y(n_385) );
OR2x2_ASAP7_75t_L g392 ( .A(n_231), .B(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g404 ( .A(n_231), .B(n_293), .Y(n_404) );
CKINVDCx16_ASAP7_75t_R g231 ( .A(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g338 ( .A(n_232), .B(n_339), .Y(n_338) );
BUFx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g266 ( .A(n_233), .B(n_267), .Y(n_266) );
INVx4_ASAP7_75t_L g287 ( .A(n_233), .Y(n_287) );
AND2x2_ASAP7_75t_L g324 ( .A(n_233), .B(n_268), .Y(n_324) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_241), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_234), .B(n_488), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_234), .B(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_234), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g323 ( .A(n_243), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_SL g393 ( .A(n_243), .Y(n_393) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_253), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_244), .B(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g293 ( .A(n_244), .B(n_254), .Y(n_293) );
INVx2_ASAP7_75t_L g313 ( .A(n_244), .Y(n_313) );
AND2x2_ASAP7_75t_L g327 ( .A(n_244), .B(n_254), .Y(n_327) );
AND2x2_ASAP7_75t_L g334 ( .A(n_244), .B(n_290), .Y(n_334) );
BUFx3_ASAP7_75t_L g344 ( .A(n_244), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_244), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g289 ( .A(n_253), .Y(n_289) );
AND2x2_ASAP7_75t_L g297 ( .A(n_253), .B(n_287), .Y(n_297) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g267 ( .A(n_254), .B(n_268), .Y(n_267) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_254), .Y(n_321) );
INVx2_ASAP7_75t_L g486 ( .A(n_261), .Y(n_486) );
INVx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx2_ASAP7_75t_SL g304 ( .A(n_265), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_265), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_265), .B(n_374), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_266), .B(n_344), .Y(n_397) );
INVx1_ASAP7_75t_SL g431 ( .A(n_266), .Y(n_431) );
INVx1_ASAP7_75t_SL g339 ( .A(n_267), .Y(n_339) );
INVx1_ASAP7_75t_SL g290 ( .A(n_268), .Y(n_290) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_268), .Y(n_301) );
OR2x2_ASAP7_75t_L g312 ( .A(n_268), .B(n_287), .Y(n_312) );
AND2x2_ASAP7_75t_L g326 ( .A(n_268), .B(n_287), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_268), .B(n_316), .Y(n_378) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_282), .B(n_284), .C(n_295), .Y(n_277) );
AOI31xp33_ASAP7_75t_L g394 ( .A1(n_278), .A2(n_395), .A3(n_396), .B(n_397), .Y(n_394) );
AND2x2_ASAP7_75t_L g367 ( .A(n_279), .B(n_296), .Y(n_367) );
BUFx3_ASAP7_75t_L g307 ( .A(n_280), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_280), .B(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g343 ( .A(n_280), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_280), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g298 ( .A(n_283), .Y(n_298) );
OAI222xp33_ASAP7_75t_L g407 ( .A1(n_283), .A2(n_408), .B1(n_411), .B2(n_412), .C1(n_413), .C2(n_414), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_285), .B(n_291), .Y(n_284) );
INVx1_ASAP7_75t_L g413 ( .A(n_285), .Y(n_413) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_287), .B(n_290), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_287), .B(n_313), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_287), .B(n_288), .Y(n_383) );
INVx1_ASAP7_75t_L g434 ( .A(n_287), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_288), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g436 ( .A(n_288), .Y(n_436) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx2_ASAP7_75t_L g316 ( .A(n_289), .Y(n_316) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_290), .Y(n_359) );
AOI32xp33_ASAP7_75t_L g295 ( .A1(n_291), .A2(n_296), .A3(n_297), .B1(n_298), .B2(n_299), .Y(n_295) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_293), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g370 ( .A(n_293), .Y(n_370) );
OR2x2_ASAP7_75t_L g411 ( .A(n_293), .B(n_312), .Y(n_411) );
INVx1_ASAP7_75t_L g347 ( .A(n_294), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_296), .B(n_307), .Y(n_332) );
INVx3_ASAP7_75t_L g341 ( .A(n_296), .Y(n_341) );
AOI322xp5_ASAP7_75t_L g357 ( .A1(n_296), .A2(n_341), .A3(n_358), .B1(n_360), .B2(n_363), .C1(n_367), .C2(n_368), .Y(n_357) );
AND2x2_ASAP7_75t_L g333 ( .A(n_297), .B(n_334), .Y(n_333) );
INVxp67_ASAP7_75t_L g410 ( .A(n_297), .Y(n_410) );
A2O1A1O1Ixp25_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_302), .B(n_305), .C(n_313), .D(n_314), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_301), .B(n_344), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
OAI221xp5_ASAP7_75t_L g314 ( .A1(n_303), .A2(n_315), .B1(n_318), .B2(n_319), .C(n_322), .Y(n_314) );
INVx1_ASAP7_75t_SL g429 ( .A(n_303), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_310), .B(n_312), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_307), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OAI221xp5_ASAP7_75t_SL g399 ( .A1(n_309), .A2(n_393), .B1(n_400), .B2(n_401), .C(n_402), .Y(n_399) );
OAI222xp33_ASAP7_75t_L g430 ( .A1(n_310), .A2(n_431), .B1(n_432), .B2(n_433), .C1(n_435), .C2(n_436), .Y(n_430) );
AND2x2_ASAP7_75t_L g388 ( .A(n_311), .B(n_374), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_311), .A2(n_326), .B(n_373), .Y(n_400) );
INVx1_ASAP7_75t_L g414 ( .A(n_311), .Y(n_414) );
INVx2_ASAP7_75t_SL g317 ( .A(n_312), .Y(n_317) );
AND2x2_ASAP7_75t_L g320 ( .A(n_313), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_SL g354 ( .A(n_316), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_316), .B(n_326), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_317), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_317), .B(n_327), .Y(n_356) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OAI21xp5_ASAP7_75t_SL g322 ( .A1(n_323), .A2(n_325), .B(n_328), .Y(n_322) );
INVx1_ASAP7_75t_SL g340 ( .A(n_324), .Y(n_340) );
AND2x2_ASAP7_75t_L g387 ( .A(n_324), .B(n_370), .Y(n_387) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
AND2x2_ASAP7_75t_L g426 ( .A(n_326), .B(n_344), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_327), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_SL g412 ( .A(n_328), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .B1(n_335), .B2(n_342), .C(n_345), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_338), .B1(n_340), .B2(n_341), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OAI22xp33_ASAP7_75t_L g345 ( .A1(n_339), .A2(n_346), .B1(n_348), .B2(n_350), .Y(n_345) );
OR2x2_ASAP7_75t_L g416 ( .A(n_340), .B(n_344), .Y(n_416) );
OR2x2_ASAP7_75t_L g419 ( .A(n_340), .B(n_354), .Y(n_419) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OAI221xp5_ASAP7_75t_L g415 ( .A1(n_361), .A2(n_416), .B1(n_417), .B2(n_419), .C(n_420), .Y(n_415) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVxp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND3xp33_ASAP7_75t_SL g371 ( .A(n_372), .B(n_386), .C(n_398), .Y(n_371) );
AOI222xp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_377), .B1(n_379), .B2(n_382), .C1(n_384), .C2(n_385), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_374), .B(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g396 ( .A(n_376), .Y(n_396) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B1(n_389), .B2(n_391), .C(n_394), .Y(n_386) );
INVx1_ASAP7_75t_L g401 ( .A(n_387), .Y(n_401) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OAI21xp33_ASAP7_75t_L g420 ( .A1(n_391), .A2(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
NOR5xp2_ASAP7_75t_L g398 ( .A(n_399), .B(n_407), .C(n_415), .D(n_424), .E(n_430), .Y(n_398) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVxp67_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g724 ( .A(n_438), .Y(n_724) );
AND2x2_ASAP7_75t_SL g438 ( .A(n_439), .B(n_656), .Y(n_438) );
NOR4xp25_ASAP7_75t_L g439 ( .A(n_440), .B(n_586), .C(n_617), .D(n_636), .Y(n_439) );
NAND4xp25_ASAP7_75t_L g440 ( .A(n_441), .B(n_544), .C(n_559), .D(n_577), .Y(n_440) );
AOI222xp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_489), .B1(n_521), .B2(n_532), .C1(n_537), .C2(n_539), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_474), .Y(n_442) );
INVx1_ASAP7_75t_L g600 ( .A(n_443), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_454), .Y(n_443) );
AND2x2_ASAP7_75t_L g475 ( .A(n_444), .B(n_466), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_444), .B(n_478), .Y(n_629) );
INVx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g536 ( .A(n_445), .B(n_456), .Y(n_536) );
AND2x2_ASAP7_75t_L g545 ( .A(n_445), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g571 ( .A(n_445), .Y(n_571) );
AND2x2_ASAP7_75t_L g592 ( .A(n_445), .B(n_456), .Y(n_592) );
BUFx2_ASAP7_75t_L g615 ( .A(n_445), .Y(n_615) );
AND2x2_ASAP7_75t_L g639 ( .A(n_445), .B(n_457), .Y(n_639) );
AND2x2_ASAP7_75t_L g703 ( .A(n_445), .B(n_466), .Y(n_703) );
AND2x2_ASAP7_75t_L g604 ( .A(n_454), .B(n_535), .Y(n_604) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_455), .B(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_466), .Y(n_455) );
OR2x2_ASAP7_75t_L g564 ( .A(n_456), .B(n_479), .Y(n_564) );
AND2x2_ASAP7_75t_L g576 ( .A(n_456), .B(n_535), .Y(n_576) );
BUFx2_ASAP7_75t_L g708 ( .A(n_456), .Y(n_708) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g477 ( .A(n_457), .B(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g558 ( .A(n_457), .B(n_479), .Y(n_558) );
AND2x2_ASAP7_75t_L g611 ( .A(n_457), .B(n_466), .Y(n_611) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_457), .Y(n_647) );
AND2x2_ASAP7_75t_L g534 ( .A(n_466), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_SL g546 ( .A(n_466), .Y(n_546) );
INVx2_ASAP7_75t_L g557 ( .A(n_466), .Y(n_557) );
BUFx2_ASAP7_75t_L g581 ( .A(n_466), .Y(n_581) );
AND2x2_ASAP7_75t_SL g638 ( .A(n_466), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
AOI332xp33_ASAP7_75t_L g559 ( .A1(n_475), .A2(n_560), .A3(n_564), .B1(n_565), .B2(n_569), .B3(n_572), .C1(n_573), .C2(n_575), .Y(n_559) );
NAND2x1_ASAP7_75t_L g644 ( .A(n_475), .B(n_535), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_475), .B(n_549), .Y(n_695) );
A2O1A1Ixp33_ASAP7_75t_SL g577 ( .A1(n_476), .A2(n_578), .B(n_581), .C(n_582), .Y(n_577) );
AND2x2_ASAP7_75t_L g716 ( .A(n_476), .B(n_557), .Y(n_716) );
INVx3_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
OR2x2_ASAP7_75t_L g613 ( .A(n_477), .B(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g618 ( .A(n_477), .B(n_615), .Y(n_618) );
INVx1_ASAP7_75t_L g549 ( .A(n_478), .Y(n_549) );
AND2x2_ASAP7_75t_L g652 ( .A(n_478), .B(n_611), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_478), .B(n_592), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_478), .B(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_478), .B(n_570), .Y(n_678) );
INVx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx3_ASAP7_75t_L g535 ( .A(n_479), .Y(n_535) );
OAI31xp33_ASAP7_75t_L g717 ( .A1(n_489), .A2(n_638), .A3(n_645), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_500), .Y(n_489) );
AND2x2_ASAP7_75t_L g521 ( .A(n_490), .B(n_522), .Y(n_521) );
NAND2x1_ASAP7_75t_SL g540 ( .A(n_490), .B(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_490), .Y(n_627) );
AND2x2_ASAP7_75t_L g632 ( .A(n_490), .B(n_543), .Y(n_632) );
INVx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_491), .A2(n_545), .B(n_547), .C(n_550), .Y(n_544) );
OR2x2_ASAP7_75t_L g561 ( .A(n_491), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g574 ( .A(n_491), .Y(n_574) );
AND2x2_ASAP7_75t_L g580 ( .A(n_491), .B(n_523), .Y(n_580) );
INVx2_ASAP7_75t_L g598 ( .A(n_491), .Y(n_598) );
AND2x2_ASAP7_75t_L g609 ( .A(n_491), .B(n_563), .Y(n_609) );
AND2x2_ASAP7_75t_L g641 ( .A(n_491), .B(n_599), .Y(n_641) );
AND2x2_ASAP7_75t_L g645 ( .A(n_491), .B(n_568), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_491), .B(n_500), .Y(n_650) );
AND2x2_ASAP7_75t_L g684 ( .A(n_491), .B(n_685), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_491), .B(n_587), .Y(n_718) );
OR2x6_ASAP7_75t_L g491 ( .A(n_492), .B(n_498), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_500), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g626 ( .A(n_500), .Y(n_626) );
AND2x2_ASAP7_75t_L g688 ( .A(n_500), .B(n_609), .Y(n_688) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_512), .Y(n_500) );
OR2x2_ASAP7_75t_L g542 ( .A(n_501), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g552 ( .A(n_501), .B(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_501), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g660 ( .A(n_501), .Y(n_660) );
AND2x2_ASAP7_75t_L g677 ( .A(n_501), .B(n_523), .Y(n_677) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g568 ( .A(n_502), .B(n_512), .Y(n_568) );
AND2x2_ASAP7_75t_L g597 ( .A(n_502), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g608 ( .A(n_502), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_502), .B(n_563), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_509), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B(n_508), .Y(n_505) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g522 ( .A(n_513), .B(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g543 ( .A(n_513), .Y(n_543) );
AND2x2_ASAP7_75t_L g599 ( .A(n_513), .B(n_563), .Y(n_599) );
INVx1_ASAP7_75t_L g701 ( .A(n_521), .Y(n_701) );
INVx1_ASAP7_75t_L g705 ( .A(n_522), .Y(n_705) );
INVx2_ASAP7_75t_L g563 ( .A(n_523), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_533), .B(n_536), .Y(n_532) );
INVx1_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_534), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_534), .B(n_639), .Y(n_697) );
OR2x2_ASAP7_75t_L g538 ( .A(n_535), .B(n_536), .Y(n_538) );
INVx1_ASAP7_75t_SL g590 ( .A(n_535), .Y(n_590) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AOI221xp5_ASAP7_75t_L g593 ( .A1(n_541), .A2(n_594), .B1(n_596), .B2(n_600), .C(n_601), .Y(n_593) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
OR2x2_ASAP7_75t_L g621 ( .A(n_542), .B(n_585), .Y(n_621) );
INVx2_ASAP7_75t_L g553 ( .A(n_543), .Y(n_553) );
INVx1_ASAP7_75t_L g579 ( .A(n_543), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_543), .B(n_563), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_543), .B(n_566), .Y(n_673) );
INVx1_ASAP7_75t_L g681 ( .A(n_543), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_545), .B(n_549), .Y(n_595) );
AND2x4_ASAP7_75t_L g570 ( .A(n_546), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g683 ( .A(n_549), .B(n_639), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_551), .B(n_554), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_552), .B(n_584), .Y(n_583) );
INVxp67_ASAP7_75t_L g691 ( .A(n_553), .Y(n_691) );
INVxp67_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g591 ( .A(n_557), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g663 ( .A(n_557), .B(n_639), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_557), .B(n_576), .Y(n_669) );
AOI322xp5_ASAP7_75t_L g623 ( .A1(n_558), .A2(n_592), .A3(n_599), .B1(n_624), .B2(n_627), .C1(n_628), .C2(n_630), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_558), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g689 ( .A(n_561), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g635 ( .A(n_562), .Y(n_635) );
INVx2_ASAP7_75t_L g566 ( .A(n_563), .Y(n_566) );
INVx1_ASAP7_75t_L g625 ( .A(n_563), .Y(n_625) );
CKINVDCx16_ASAP7_75t_R g572 ( .A(n_564), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
AND2x2_ASAP7_75t_L g661 ( .A(n_566), .B(n_574), .Y(n_661) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g573 ( .A(n_568), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g616 ( .A(n_568), .B(n_609), .Y(n_616) );
AND2x2_ASAP7_75t_L g620 ( .A(n_568), .B(n_580), .Y(n_620) );
OAI21xp33_ASAP7_75t_SL g630 ( .A1(n_569), .A2(n_631), .B(n_633), .Y(n_630) );
OAI22xp33_ASAP7_75t_L g700 ( .A1(n_569), .A2(n_701), .B1(n_702), .B2(n_704), .Y(n_700) );
INVx3_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g575 ( .A(n_570), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_570), .B(n_590), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_572), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx1_ASAP7_75t_L g712 ( .A(n_579), .Y(n_712) );
INVx4_ASAP7_75t_L g585 ( .A(n_580), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_580), .B(n_607), .Y(n_655) );
INVx1_ASAP7_75t_SL g667 ( .A(n_581), .Y(n_667) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NOR2xp67_ASAP7_75t_L g680 ( .A(n_585), .B(n_681), .Y(n_680) );
OAI211xp5_ASAP7_75t_SL g586 ( .A1(n_587), .A2(n_588), .B(n_593), .C(n_610), .Y(n_586) );
OAI221xp5_ASAP7_75t_SL g706 ( .A1(n_588), .A2(n_626), .B1(n_705), .B2(n_707), .C(n_709), .Y(n_706) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_590), .B(n_703), .Y(n_702) );
OAI31xp33_ASAP7_75t_L g682 ( .A1(n_591), .A2(n_668), .A3(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g622 ( .A(n_592), .Y(n_622) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
INVx1_ASAP7_75t_L g672 ( .A(n_597), .Y(n_672) );
AND2x2_ASAP7_75t_L g685 ( .A(n_599), .B(n_608), .Y(n_685) );
AOI21xp33_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_603), .B(n_605), .Y(n_601) );
INVx1_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
INVxp67_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_609), .B(n_712), .Y(n_711) );
OAI21xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B(n_616), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI221xp5_ASAP7_75t_SL g617 ( .A1(n_618), .A2(n_619), .B1(n_621), .B2(n_622), .C(n_623), .Y(n_617) );
A2O1A1Ixp33_ASAP7_75t_L g686 ( .A1(n_618), .A2(n_687), .B(n_689), .C(n_692), .Y(n_686) );
CKINVDCx16_ASAP7_75t_R g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_621), .B(n_671), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
INVx1_ASAP7_75t_L g648 ( .A(n_629), .Y(n_648) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g634 ( .A(n_632), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g676 ( .A(n_632), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OAI211xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_640), .B(n_642), .C(n_651), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI221xp5_ASAP7_75t_L g713 ( .A1(n_640), .A2(n_650), .B1(n_714), .B2(n_715), .C(n_717), .Y(n_713) );
INVx1_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B1(n_646), .B2(n_649), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI21xp5_ASAP7_75t_SL g651 ( .A1(n_652), .A2(n_653), .B(n_654), .Y(n_651) );
INVx1_ASAP7_75t_SL g714 ( .A(n_653), .Y(n_714) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NOR4xp25_ASAP7_75t_L g656 ( .A(n_657), .B(n_686), .C(n_706), .D(n_713), .Y(n_656) );
OAI211xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_662), .B(n_664), .C(n_682), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .Y(n_658) );
INVxp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
O2A1O1Ixp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_668), .B(n_670), .C(n_674), .Y(n_664) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_SL g693 ( .A(n_671), .Y(n_693) );
OR2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
OR2x2_ASAP7_75t_L g704 ( .A(n_672), .B(n_705), .Y(n_704) );
OAI21xp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_678), .B(n_679), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_694), .B1(n_696), .B2(n_698), .C(n_700), .Y(n_692) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_703), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
endmodule