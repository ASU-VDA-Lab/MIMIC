module real_aes_3640_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g249 ( .A(n_0), .Y(n_249) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_0), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g159 ( .A1(n_1), .A2(n_18), .B1(n_84), .B2(n_151), .Y(n_159) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_2), .A2(n_51), .B1(n_572), .B2(n_576), .Y(n_571) );
INVx2_ASAP7_75t_L g130 ( .A(n_3), .Y(n_130) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_4), .A2(n_72), .B1(n_546), .B2(n_549), .Y(n_545) );
INVx1_ASAP7_75t_SL g206 ( .A(n_5), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_6), .A2(n_65), .B1(n_534), .B2(n_536), .Y(n_533) );
AO22x1_ASAP7_75t_L g588 ( .A1(n_7), .A2(n_50), .B1(n_589), .B2(n_590), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_8), .B(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_9), .B(n_225), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_10), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_11), .A2(n_557), .B(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g530 ( .A(n_12), .Y(n_530) );
INVxp67_ASAP7_75t_L g543 ( .A(n_12), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_12), .B(n_57), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_13), .A2(n_44), .B1(n_220), .B2(n_221), .Y(n_219) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_14), .Y(n_600) );
AO22x1_ASAP7_75t_L g577 ( .A1(n_15), .A2(n_48), .B1(n_578), .B2(n_581), .Y(n_577) );
OA21x2_ASAP7_75t_L g111 ( .A1(n_16), .A2(n_55), .B(n_112), .Y(n_111) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_16), .A2(n_55), .B(n_112), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_17), .B(n_515), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_19), .B(n_126), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g114 ( .A1(n_20), .A2(n_61), .B1(n_115), .B2(n_118), .Y(n_114) );
INVx2_ASAP7_75t_L g155 ( .A(n_21), .Y(n_155) );
AOI22xp5_ASAP7_75t_L g160 ( .A1(n_22), .A2(n_25), .B1(n_161), .B2(n_163), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_23), .B(n_511), .Y(n_510) );
BUFx3_ASAP7_75t_L g612 ( .A(n_24), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_26), .A2(n_52), .B1(n_123), .B2(n_125), .Y(n_122) );
O2A1O1Ixp5_ASAP7_75t_L g148 ( .A1(n_27), .A2(n_88), .B(n_149), .C(n_150), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_28), .Y(n_192) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_29), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_30), .A2(n_63), .B1(n_228), .B2(n_230), .Y(n_227) );
INVx1_ASAP7_75t_L g142 ( .A(n_31), .Y(n_142) );
INVx1_ASAP7_75t_L g516 ( .A(n_32), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_32), .B(n_56), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_33), .A2(n_507), .B1(n_592), .B2(n_625), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_33), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_34), .B(n_138), .Y(n_244) );
INVx2_ASAP7_75t_L g152 ( .A(n_35), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_36), .Y(n_194) );
INVx1_ASAP7_75t_L g559 ( .A(n_37), .Y(n_559) );
INVx2_ASAP7_75t_L g272 ( .A(n_38), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_39), .B(n_242), .Y(n_241) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_39), .Y(n_637) );
INVx1_ASAP7_75t_SL g210 ( .A(n_40), .Y(n_210) );
INVx1_ASAP7_75t_L g188 ( .A(n_41), .Y(n_188) );
AO22x1_ASAP7_75t_L g582 ( .A1(n_42), .A2(n_75), .B1(n_583), .B2(n_586), .Y(n_582) );
INVx1_ASAP7_75t_L g112 ( .A(n_43), .Y(n_112) );
AND2x4_ASAP7_75t_L g91 ( .A(n_45), .B(n_92), .Y(n_91) );
AND2x4_ASAP7_75t_L g146 ( .A(n_45), .B(n_92), .Y(n_146) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_45), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_46), .A2(n_596), .B1(n_599), .B2(n_600), .Y(n_595) );
INVx2_ASAP7_75t_L g598 ( .A(n_46), .Y(n_598) );
INVx1_ASAP7_75t_L g215 ( .A(n_47), .Y(n_215) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_49), .Y(n_89) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_53), .B(n_208), .Y(n_276) );
OA22x2_ASAP7_75t_L g520 ( .A1(n_54), .A2(n_57), .B1(n_515), .B2(n_519), .Y(n_520) );
INVx1_ASAP7_75t_L g554 ( .A(n_54), .Y(n_554) );
INVx1_ASAP7_75t_L g532 ( .A(n_56), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_56), .B(n_552), .Y(n_568) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_56), .Y(n_615) );
OAI21xp33_ASAP7_75t_L g555 ( .A1(n_57), .A2(n_62), .B(n_544), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_58), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_59), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_60), .B(n_119), .Y(n_212) );
INVx1_ASAP7_75t_L g518 ( .A(n_62), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_62), .B(n_74), .Y(n_566) );
BUFx6f_ASAP7_75t_L g85 ( .A(n_64), .Y(n_85) );
INVx1_ASAP7_75t_L g117 ( .A(n_64), .Y(n_117) );
BUFx5_ASAP7_75t_L g162 ( .A(n_64), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_66), .B(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g275 ( .A(n_67), .Y(n_275) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_68), .Y(n_602) );
INVx1_ASAP7_75t_L g279 ( .A(n_69), .Y(n_279) );
INVx2_ASAP7_75t_L g198 ( .A(n_70), .Y(n_198) );
INVx2_ASAP7_75t_SL g92 ( .A(n_71), .Y(n_92) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_73), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_74), .B(n_525), .Y(n_524) );
AO32x2_ASAP7_75t_L g157 ( .A1(n_76), .A2(n_90), .A3(n_153), .B1(n_158), .B2(n_165), .Y(n_157) );
AO22x2_ASAP7_75t_L g298 ( .A1(n_76), .A2(n_158), .B1(n_299), .B2(n_301), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_93), .B(n_502), .Y(n_77) );
BUFx2_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
AND2x2_ASAP7_75t_L g79 ( .A(n_80), .B(n_90), .Y(n_79) );
OA21x2_ASAP7_75t_L g632 ( .A1(n_80), .A2(n_633), .B(n_634), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g80 ( .A(n_81), .B(n_86), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx2_ASAP7_75t_L g144 ( .A(n_84), .Y(n_144) );
INVxp67_ASAP7_75t_SL g230 ( .A(n_84), .Y(n_230) );
INVx2_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx3_ASAP7_75t_L g119 ( .A(n_85), .Y(n_119) );
INVx6_ASAP7_75t_L g126 ( .A(n_85), .Y(n_126) );
INVx2_ASAP7_75t_L g186 ( .A(n_85), .Y(n_186) );
HB1xp67_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_87), .B(n_145), .Y(n_190) );
INVx4_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
OAI22xp5_ASAP7_75t_L g158 ( .A1(n_88), .A2(n_159), .B1(n_160), .B2(n_164), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_88), .A2(n_239), .B(n_241), .Y(n_238) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_89), .Y(n_121) );
INVx3_ASAP7_75t_L g128 ( .A(n_89), .Y(n_128) );
INVx4_ASAP7_75t_L g139 ( .A(n_89), .Y(n_139) );
INVx1_ASAP7_75t_L g232 ( .A(n_89), .Y(n_232) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
AND2x2_ASAP7_75t_L g107 ( .A(n_91), .B(n_108), .Y(n_107) );
INVx3_ASAP7_75t_L g203 ( .A(n_91), .Y(n_203) );
AND2x2_ASAP7_75t_L g299 ( .A(n_91), .B(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_92), .Y(n_620) );
INVxp33_ASAP7_75t_SL g93 ( .A(n_94), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
OR2x2_ASAP7_75t_L g97 ( .A(n_98), .B(n_396), .Y(n_97) );
NAND3xp33_ASAP7_75t_L g98 ( .A(n_99), .B(n_293), .C(n_348), .Y(n_98) );
AOI211xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_172), .B(n_261), .C(n_291), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g100 ( .A(n_101), .B(n_168), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_156), .Y(n_102) );
AND2x4_ASAP7_75t_L g354 ( .A(n_103), .B(n_318), .Y(n_354) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g296 ( .A(n_104), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_105), .B(n_132), .Y(n_104) );
OR2x2_ASAP7_75t_L g170 ( .A(n_105), .B(n_132), .Y(n_170) );
AND2x2_ASAP7_75t_L g347 ( .A(n_105), .B(n_298), .Y(n_347) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g266 ( .A(n_106), .Y(n_266) );
INVx1_ASAP7_75t_L g323 ( .A(n_106), .Y(n_323) );
AOI21x1_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_113), .B(n_129), .Y(n_106) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_109), .B(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx4_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g131 ( .A(n_111), .Y(n_131) );
BUFx3_ASAP7_75t_L g196 ( .A(n_111), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_120), .B1(n_122), .B2(n_127), .Y(n_113) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g182 ( .A(n_116), .Y(n_182) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g124 ( .A(n_117), .Y(n_124) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g163 ( .A(n_119), .Y(n_163) );
INVx1_ASAP7_75t_L g221 ( .A(n_119), .Y(n_221) );
INVx1_ASAP7_75t_L g240 ( .A(n_119), .Y(n_240) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g164 ( .A(n_121), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_121), .A2(n_205), .B(n_206), .C(n_207), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_121), .B(n_223), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_121), .A2(n_182), .B(n_275), .C(n_276), .Y(n_274) );
INVx3_ASAP7_75t_L g149 ( .A(n_123), .Y(n_149) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g208 ( .A(n_124), .Y(n_208) );
INVx1_ASAP7_75t_L g271 ( .A(n_125), .Y(n_271) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g136 ( .A(n_126), .Y(n_136) );
INVx2_ASAP7_75t_SL g151 ( .A(n_126), .Y(n_151) );
INVx2_ASAP7_75t_L g193 ( .A(n_126), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_127), .B(n_145), .Y(n_183) );
NOR3xp33_ASAP7_75t_L g187 ( .A(n_127), .B(n_145), .C(n_188), .Y(n_187) );
INVx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_128), .A2(n_210), .B(n_211), .C(n_212), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_128), .A2(n_271), .B(n_272), .C(n_273), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
BUFx3_ASAP7_75t_L g153 ( .A(n_131), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_131), .B(n_155), .Y(n_154) );
INVx3_ASAP7_75t_L g236 ( .A(n_131), .Y(n_236) );
INVx1_ASAP7_75t_L g280 ( .A(n_132), .Y(n_280) );
INVx2_ASAP7_75t_L g286 ( .A(n_132), .Y(n_286) );
AND2x2_ASAP7_75t_L g308 ( .A(n_132), .B(n_302), .Y(n_308) );
AND2x2_ASAP7_75t_L g317 ( .A(n_132), .B(n_268), .Y(n_317) );
AO31x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_147), .A3(n_153), .B(n_154), .Y(n_132) );
AOI221x1_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_137), .B1(n_141), .B2(n_143), .C(n_145), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
AND2x2_ASAP7_75t_L g141 ( .A(n_138), .B(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_139), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx4_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
INVx2_ASAP7_75t_L g301 ( .A(n_153), .Y(n_301) );
INVx2_ASAP7_75t_L g171 ( .A(n_156), .Y(n_171) );
AND2x2_ASAP7_75t_L g307 ( .A(n_156), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g341 ( .A(n_156), .B(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g419 ( .A(n_156), .B(n_322), .Y(n_419) );
AND2x2_ASAP7_75t_L g472 ( .A(n_156), .B(n_317), .Y(n_472) );
AND2x2_ASAP7_75t_SL g488 ( .A(n_156), .B(n_267), .Y(n_488) );
BUFx3_ASAP7_75t_L g498 ( .A(n_156), .Y(n_498) );
BUFx8_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g284 ( .A(n_157), .Y(n_284) );
AND2x2_ASAP7_75t_L g388 ( .A(n_157), .B(n_389), .Y(n_388) );
OAI22xp33_ASAP7_75t_L g191 ( .A1(n_161), .A2(n_192), .B1(n_193), .B2(n_194), .Y(n_191) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g211 ( .A(n_162), .Y(n_211) );
INVx2_ASAP7_75t_L g220 ( .A(n_162), .Y(n_220) );
INVx2_ASAP7_75t_L g242 ( .A(n_162), .Y(n_242) );
INVx1_ASAP7_75t_L g246 ( .A(n_162), .Y(n_246) );
INVx1_ASAP7_75t_L g205 ( .A(n_163), .Y(n_205) );
INVxp67_ASAP7_75t_L g260 ( .A(n_165), .Y(n_260) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_166), .B(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g214 ( .A(n_167), .Y(n_214) );
NOR2xp67_ASAP7_75t_L g223 ( .A(n_167), .B(n_203), .Y(n_223) );
BUFx3_ASAP7_75t_L g225 ( .A(n_167), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_167), .B(n_203), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_167), .B(n_203), .Y(n_277) );
INVx1_ASAP7_75t_L g300 ( .A(n_167), .Y(n_300) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NAND3xp33_ASAP7_75t_SL g483 ( .A(n_169), .B(n_484), .C(n_487), .Y(n_483) );
OR2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
INVx2_ASAP7_75t_L g362 ( .A(n_170), .Y(n_362) );
NAND2x1_ASAP7_75t_L g172 ( .A(n_173), .B(n_251), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_173), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_216), .Y(n_174) );
INVx1_ASAP7_75t_L g309 ( .A(n_175), .Y(n_309) );
AND2x2_ASAP7_75t_L g439 ( .A(n_175), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g477 ( .A(n_175), .B(n_330), .Y(n_477) );
AND2x4_ASAP7_75t_L g175 ( .A(n_176), .B(n_199), .Y(n_175) );
OR2x2_ASAP7_75t_L g344 ( .A(n_176), .B(n_258), .Y(n_344) );
AND2x2_ASAP7_75t_L g431 ( .A(n_176), .B(n_305), .Y(n_431) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g332 ( .A(n_177), .B(n_290), .Y(n_332) );
BUFx2_ASAP7_75t_L g336 ( .A(n_177), .Y(n_336) );
OR2x2_ASAP7_75t_L g353 ( .A(n_177), .B(n_201), .Y(n_353) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_195), .B(n_197), .Y(n_177) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_178), .A2(n_197), .B(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_189), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_183), .B1(n_184), .B2(n_187), .Y(n_179) );
NOR2xp67_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g229 ( .A(n_186), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_193), .B(n_248), .Y(n_247) );
INVx3_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g383 ( .A(n_200), .B(n_234), .Y(n_383) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g256 ( .A(n_201), .Y(n_256) );
INVx2_ASAP7_75t_L g290 ( .A(n_201), .Y(n_290) );
AND2x2_ASAP7_75t_L g364 ( .A(n_201), .B(n_259), .Y(n_364) );
INVx1_ASAP7_75t_L g416 ( .A(n_201), .Y(n_416) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_201), .Y(n_450) );
AO31x2_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_204), .A3(n_209), .B(n_213), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_210), .A2(n_602), .B1(n_603), .B2(n_604), .Y(n_601) );
INVx1_ASAP7_75t_L g604 ( .A(n_210), .Y(n_604) );
NOR2xp33_ASAP7_75t_SL g213 ( .A(n_214), .B(n_215), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_214), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_216), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g368 ( .A(n_216), .B(n_364), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_216), .B(n_336), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_216), .B(n_335), .Y(n_499) );
NAND2xp67_ASAP7_75t_L g500 ( .A(n_216), .B(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_233), .Y(n_216) );
INVx1_ASAP7_75t_L g254 ( .A(n_217), .Y(n_254) );
INVx2_ASAP7_75t_L g305 ( .A(n_217), .Y(n_305) );
INVx1_ASAP7_75t_L g313 ( .A(n_217), .Y(n_313) );
AND2x2_ASAP7_75t_L g375 ( .A(n_217), .B(n_234), .Y(n_375) );
NAND2x1p5_ASAP7_75t_L g217 ( .A(n_218), .B(n_226), .Y(n_217) );
AND2x2_ASAP7_75t_SL g412 ( .A(n_218), .B(n_226), .Y(n_412) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_222), .B(n_224), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_223), .B(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_231), .Y(n_226) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
OR2x2_ASAP7_75t_L g315 ( .A(n_233), .B(n_259), .Y(n_315) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g258 ( .A(n_234), .Y(n_258) );
INVx1_ASAP7_75t_L g339 ( .A(n_234), .Y(n_339) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_234), .Y(n_407) );
AND2x4_ASAP7_75t_L g234 ( .A(n_235), .B(n_237), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_243), .B(n_250), .Y(n_237) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_247), .Y(n_243) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_252), .A2(n_445), .B1(n_447), .B2(n_449), .Y(n_444) );
AND2x4_ASAP7_75t_L g252 ( .A(n_253), .B(n_257), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
BUFx3_ASAP7_75t_L g359 ( .A(n_254), .Y(n_359) );
AND2x2_ASAP7_75t_L g406 ( .A(n_255), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
AND2x2_ASAP7_75t_L g415 ( .A(n_258), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g304 ( .A(n_259), .B(n_305), .Y(n_304) );
AOI21xp33_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_281), .B(n_287), .Y(n_261) );
OAI21xp5_ASAP7_75t_L g384 ( .A1(n_262), .A2(n_385), .B(n_386), .Y(n_384) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
AND2x4_ASAP7_75t_L g282 ( .A(n_264), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_264), .B(n_297), .Y(n_417) );
INVx4_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g373 ( .A(n_265), .B(n_267), .Y(n_373) );
INVx2_ASAP7_75t_L g424 ( .A(n_265), .Y(n_424) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_265), .B(n_308), .Y(n_478) );
BUFx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g389 ( .A(n_266), .Y(n_389) );
INVx2_ASAP7_75t_L g292 ( .A(n_267), .Y(n_292) );
INVx2_ASAP7_75t_L g342 ( .A(n_267), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_267), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_267), .B(n_332), .Y(n_435) );
AND2x4_ASAP7_75t_L g267 ( .A(n_268), .B(n_280), .Y(n_267) );
INVx2_ASAP7_75t_L g302 ( .A(n_268), .Y(n_302) );
INVx1_ASAP7_75t_L g325 ( .A(n_268), .Y(n_325) );
BUFx3_ASAP7_75t_L g356 ( .A(n_268), .Y(n_356) );
AND2x4_ASAP7_75t_L g426 ( .A(n_268), .B(n_284), .Y(n_426) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AO31x2_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_274), .A3(n_277), .B(n_278), .Y(n_269) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g372 ( .A(n_283), .Y(n_372) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_284), .B(n_389), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_285), .B(n_381), .Y(n_380) );
INVx2_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g322 ( .A(n_286), .B(n_323), .Y(n_322) );
BUFx3_ASAP7_75t_L g366 ( .A(n_286), .Y(n_366) );
INVx1_ASAP7_75t_L g448 ( .A(n_286), .Y(n_448) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NOR2xp67_ASAP7_75t_L g378 ( .A(n_289), .B(n_344), .Y(n_378) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g394 ( .A(n_290), .B(n_381), .Y(n_394) );
INVxp67_ASAP7_75t_SL g494 ( .A(n_290), .Y(n_494) );
NOR3xp33_ASAP7_75t_L g293 ( .A(n_294), .B(n_310), .C(n_319), .Y(n_293) );
OAI22xp33_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_303), .B1(n_306), .B2(n_309), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx2_ASAP7_75t_L g469 ( .A(n_296), .Y(n_469) );
AND2x4_ASAP7_75t_L g361 ( .A(n_297), .B(n_362), .Y(n_361) );
INVx4_ASAP7_75t_L g377 ( .A(n_297), .Y(n_377) );
AND2x4_ASAP7_75t_L g297 ( .A(n_298), .B(n_302), .Y(n_297) );
INVx1_ASAP7_75t_L g318 ( .A(n_298), .Y(n_318) );
INVx1_ASAP7_75t_L g326 ( .A(n_298), .Y(n_326) );
AND2x4_ASAP7_75t_L g355 ( .A(n_298), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g367 ( .A(n_302), .B(n_323), .Y(n_367) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_304), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g467 ( .A(n_304), .B(n_383), .Y(n_467) );
BUFx2_ASAP7_75t_L g330 ( .A(n_305), .Y(n_330) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_305), .Y(n_456) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NOR2x1_ASAP7_75t_L g320 ( .A(n_307), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g387 ( .A(n_308), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g427 ( .A(n_308), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g462 ( .A(n_308), .B(n_381), .Y(n_462) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_316), .Y(n_310) );
INVx3_ASAP7_75t_L g385 ( .A(n_311), .Y(n_385) );
AND2x4_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
AND2x2_ASAP7_75t_L g409 ( .A(n_312), .B(n_364), .Y(n_409) );
INVx1_ASAP7_75t_L g491 ( .A(n_312), .Y(n_491) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g382 ( .A(n_313), .B(n_383), .Y(n_382) );
INVxp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g392 ( .A(n_315), .Y(n_392) );
INVxp67_ASAP7_75t_SL g457 ( .A(n_315), .Y(n_457) );
OR2x6_ASAP7_75t_L g493 ( .A(n_315), .B(n_494), .Y(n_493) );
OAI31xp33_ASAP7_75t_L g408 ( .A1(n_316), .A2(n_328), .A3(n_409), .B(n_410), .Y(n_408) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx2_ASAP7_75t_L g403 ( .A(n_317), .Y(n_403) );
INVx2_ASAP7_75t_L g486 ( .A(n_317), .Y(n_486) );
OAI21xp5_ASAP7_75t_SL g319 ( .A1(n_320), .A2(n_327), .B(n_333), .Y(n_319) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
INVxp67_ASAP7_75t_SL g496 ( .A(n_322), .Y(n_496) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_323), .Y(n_358) );
INVx2_ASAP7_75t_L g381 ( .A(n_323), .Y(n_381) );
AOI33xp33_ASAP7_75t_L g376 ( .A1(n_324), .A2(n_377), .A3(n_378), .B1(n_379), .B2(n_380), .B3(n_382), .Y(n_376) );
AND2x2_ASAP7_75t_L g443 ( .A(n_324), .B(n_381), .Y(n_443) );
AND2x2_ASAP7_75t_L g445 ( .A(n_324), .B(n_446), .Y(n_445) );
AND2x4_ASAP7_75t_SL g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVxp67_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
NOR2x1p5_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g363 ( .A(n_330), .B(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g357 ( .A(n_332), .B(n_358), .Y(n_357) );
NAND2x1p5_ASAP7_75t_L g420 ( .A(n_332), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g481 ( .A(n_332), .B(n_375), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_340), .B1(n_343), .B2(n_345), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g401 ( .A(n_336), .B(n_375), .Y(n_401) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_338), .B(n_359), .Y(n_433) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g440 ( .A(n_339), .B(n_412), .Y(n_440) );
AND2x2_ASAP7_75t_L g474 ( .A(n_339), .B(n_412), .Y(n_474) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NOR2xp67_ASAP7_75t_SL g410 ( .A(n_344), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVxp67_ASAP7_75t_L g434 ( .A(n_347), .Y(n_434) );
NOR3xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_369), .C(n_384), .Y(n_348) );
OAI21xp5_ASAP7_75t_SL g349 ( .A1(n_350), .A2(n_359), .B(n_360), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_354), .B1(n_355), .B2(n_357), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g501 ( .A(n_353), .Y(n_501) );
INVx2_ASAP7_75t_L g452 ( .A(n_355), .Y(n_452) );
INVx1_ASAP7_75t_L g485 ( .A(n_358), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_363), .B1(n_365), .B2(n_368), .Y(n_360) );
AND2x2_ASAP7_75t_L g374 ( .A(n_364), .B(n_375), .Y(n_374) );
OAI21xp5_ASAP7_75t_L g479 ( .A1(n_365), .A2(n_480), .B(n_481), .Y(n_479) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_376), .Y(n_369) );
OAI21xp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_373), .B(n_374), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g395 ( .A(n_375), .Y(n_395) );
AND2x2_ASAP7_75t_L g449 ( .A(n_375), .B(n_450), .Y(n_449) );
NOR3xp33_ASAP7_75t_L g393 ( .A(n_377), .B(n_394), .C(n_395), .Y(n_393) );
OAI221xp5_ASAP7_75t_L g437 ( .A1(n_377), .A2(n_438), .B1(n_441), .B2(n_442), .C(n_444), .Y(n_437) );
INVx2_ASAP7_75t_L g399 ( .A(n_379), .Y(n_399) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g446 ( .A(n_381), .Y(n_446) );
BUFx3_ASAP7_75t_L g471 ( .A(n_381), .Y(n_471) );
AND2x2_ASAP7_75t_L g480 ( .A(n_383), .B(n_431), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_390), .B(n_393), .Y(n_386) );
AND2x4_ASAP7_75t_SL g447 ( .A(n_388), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g454 ( .A(n_394), .Y(n_454) );
NAND4xp25_ASAP7_75t_L g396 ( .A(n_397), .B(n_436), .C(n_464), .D(n_482), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_398), .B(n_413), .Y(n_397) );
OAI221xp5_ASAP7_75t_SL g398 ( .A1(n_399), .A2(n_400), .B1(n_402), .B2(n_405), .C(n_408), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g428 ( .A(n_404), .Y(n_428) );
INVx1_ASAP7_75t_L g459 ( .A(n_404), .Y(n_459) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g430 ( .A(n_407), .Y(n_430) );
INVx1_ASAP7_75t_SL g441 ( .A(n_409), .Y(n_441) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g421 ( .A(n_412), .Y(n_421) );
OAI221xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_417), .B1(n_418), .B2(n_420), .C(n_422), .Y(n_413) );
AND2x2_ASAP7_75t_L g473 ( .A(n_416), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g463 ( .A(n_420), .Y(n_463) );
O2A1O1Ixp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_427), .B(n_429), .C(n_432), .Y(n_422) );
NOR2x1_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B(n_435), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_451), .Y(n_436) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVxp67_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
OAI21xp33_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B(n_458), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
AND2x4_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B1(n_462), .B2(n_463), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AOI221xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_468), .B1(n_470), .B2(n_473), .C(n_475), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
OAI21xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_478), .B(n_479), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_489), .B1(n_495), .B2(n_497), .Y(n_482) );
OR2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_492), .Y(n_489) );
INVxp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVxp67_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OAI21xp33_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .B(n_500), .Y(n_497) );
OAI221xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_606), .B1(n_623), .B2(n_626), .C(n_628), .Y(n_502) );
XOR2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_593), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_507), .B1(n_591), .B2(n_592), .Y(n_504) );
INVx1_ASAP7_75t_L g591 ( .A(n_505), .Y(n_591) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g592 ( .A(n_507), .Y(n_592) );
AO22x1_ASAP7_75t_L g636 ( .A1(n_507), .A2(n_592), .B1(n_637), .B2(n_638), .Y(n_636) );
INVxp33_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_569), .Y(n_508) );
AND4x1_ASAP7_75t_L g509 ( .A(n_510), .B(n_533), .C(n_545), .D(n_556), .Y(n_509) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_521), .Y(n_511) );
AND2x4_ASAP7_75t_L g534 ( .A(n_512), .B(n_535), .Y(n_534) );
AND2x4_ASAP7_75t_L g572 ( .A(n_512), .B(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g578 ( .A(n_512), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_520), .Y(n_512) );
INVx1_ASAP7_75t_L g548 ( .A(n_513), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_517), .Y(n_513) );
NAND2xp33_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
INVx2_ASAP7_75t_L g519 ( .A(n_515), .Y(n_519) );
INVx3_ASAP7_75t_L g525 ( .A(n_515), .Y(n_525) );
NAND2xp33_ASAP7_75t_L g531 ( .A(n_515), .B(n_532), .Y(n_531) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_515), .Y(n_539) );
INVx1_ASAP7_75t_L g544 ( .A(n_515), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_516), .B(n_554), .Y(n_553) );
INVxp67_ASAP7_75t_L g616 ( .A(n_516), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g542 ( .A1(n_518), .A2(n_543), .B(n_544), .Y(n_542) );
AND2x2_ASAP7_75t_L g541 ( .A(n_520), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g547 ( .A(n_520), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g585 ( .A(n_520), .Y(n_585) );
AND2x4_ASAP7_75t_L g549 ( .A(n_521), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g557 ( .A(n_521), .B(n_547), .Y(n_557) );
AND2x4_ASAP7_75t_L g590 ( .A(n_521), .B(n_584), .Y(n_590) );
AND2x4_ASAP7_75t_L g521 ( .A(n_522), .B(n_527), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x4_ASAP7_75t_L g535 ( .A(n_523), .B(n_527), .Y(n_535) );
AND2x2_ASAP7_75t_L g537 ( .A(n_523), .B(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g574 ( .A(n_523), .B(n_575), .Y(n_574) );
AND2x4_ASAP7_75t_L g579 ( .A(n_523), .B(n_580), .Y(n_579) );
AND2x4_ASAP7_75t_L g523 ( .A(n_524), .B(n_526), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_525), .B(n_530), .Y(n_529) );
INVxp67_ASAP7_75t_L g552 ( .A(n_525), .Y(n_552) );
NAND3xp33_ASAP7_75t_L g567 ( .A(n_526), .B(n_551), .C(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g575 ( .A(n_528), .Y(n_575) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
AND2x4_ASAP7_75t_L g546 ( .A(n_535), .B(n_547), .Y(n_546) );
AND2x4_ASAP7_75t_L g589 ( .A(n_535), .B(n_584), .Y(n_589) );
AND2x4_ASAP7_75t_L g536 ( .A(n_537), .B(n_541), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g563 ( .A(n_539), .Y(n_563) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_540), .Y(n_613) );
AND2x4_ASAP7_75t_L g584 ( .A(n_548), .B(n_585), .Y(n_584) );
AND2x4_ASAP7_75t_L g576 ( .A(n_550), .B(n_573), .Y(n_576) );
AND2x4_ASAP7_75t_L g581 ( .A(n_550), .B(n_579), .Y(n_581) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_555), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_554), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx4_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AO21x2_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_564), .B(n_567), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NOR4xp25_ASAP7_75t_L g569 ( .A(n_570), .B(n_577), .C(n_582), .D(n_588), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g587 ( .A(n_574), .Y(n_587) );
INVx1_ASAP7_75t_L g580 ( .A(n_575), .Y(n_580) );
AND2x4_ASAP7_75t_L g583 ( .A(n_579), .B(n_584), .Y(n_583) );
AND2x4_ASAP7_75t_L g586 ( .A(n_584), .B(n_587), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_595), .B1(n_601), .B2(n_605), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_601), .Y(n_605) );
CKINVDCx14_ASAP7_75t_R g603 ( .A(n_602), .Y(n_603) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
BUFx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_618), .Y(n_609) );
INVxp67_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g635 ( .A(n_611), .B(n_618), .Y(n_635) );
AOI211xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B(n_614), .C(n_617), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
OR2x2_ASAP7_75t_L g627 ( .A(n_619), .B(n_622), .Y(n_627) );
INVx1_ASAP7_75t_L g633 ( .A(n_619), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_619), .B(n_621), .Y(n_634) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B1(n_635), .B2(n_636), .Y(n_628) );
CKINVDCx20_ASAP7_75t_R g630 ( .A(n_631), .Y(n_630) );
BUFx3_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
CKINVDCx5p33_ASAP7_75t_R g638 ( .A(n_637), .Y(n_638) );
endmodule