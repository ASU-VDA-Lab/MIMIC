module fake_jpeg_771_n_691 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_691);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_691;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_7),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_12),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_23),
.B(n_11),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_60),
.B(n_66),
.Y(n_145)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_65),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_23),
.B(n_53),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_71),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_72),
.Y(n_168)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_73),
.Y(n_171)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_74),
.Y(n_142)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_77),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_23),
.B(n_11),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_78),
.B(n_86),
.Y(n_148)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_79),
.Y(n_225)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_81),
.Y(n_172)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_83),
.Y(n_220)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_85),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_11),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_87),
.Y(n_174)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_88),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_89),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_90),
.Y(n_185)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_91),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_92),
.Y(n_197)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_94),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_95),
.Y(n_187)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_96),
.Y(n_173)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_22),
.B(n_10),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_32),
.Y(n_137)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_46),
.Y(n_100)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_100),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_102),
.Y(n_178)
);

BUFx12f_ASAP7_75t_SL g103 ( 
.A(n_24),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_103),
.B(n_128),
.Y(n_150)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_105),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_106),
.Y(n_189)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_107),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_108),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_27),
.Y(n_109)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_109),
.Y(n_226)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_110),
.Y(n_183)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_20),
.Y(n_111)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_24),
.Y(n_112)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_112),
.Y(n_193)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_113),
.Y(n_207)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_114),
.Y(n_216)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_35),
.Y(n_115)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_58),
.Y(n_117)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_27),
.Y(n_119)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_119),
.Y(n_201)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_35),
.Y(n_120)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_121),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_22),
.B(n_12),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_26),
.Y(n_152)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_20),
.Y(n_123)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_35),
.Y(n_124)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_124),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_27),
.Y(n_125)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_125),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_20),
.Y(n_126)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_38),
.Y(n_127)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_127),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_28),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_28),
.Y(n_129)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_129),
.Y(n_208)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_28),
.Y(n_130)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_130),
.Y(n_213)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_29),
.Y(n_131)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_131),
.Y(n_217)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_38),
.Y(n_132)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_132),
.Y(n_218)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_38),
.Y(n_133)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_133),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_137),
.B(n_144),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_60),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_117),
.A2(n_59),
.B1(n_50),
.B2(n_26),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g305 ( 
.A1(n_149),
.A2(n_158),
.B1(n_165),
.B2(n_188),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_152),
.B(n_154),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_78),
.B(n_47),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_86),
.B(n_21),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_155),
.B(n_157),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_66),
.B(n_21),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_68),
.A2(n_59),
.B1(n_50),
.B2(n_26),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_89),
.B(n_32),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_162),
.B(n_179),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_124),
.A2(n_50),
.B1(n_30),
.B2(n_49),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_L g167 ( 
.A1(n_73),
.A2(n_56),
.B1(n_54),
.B2(n_44),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_167),
.A2(n_108),
.B1(n_114),
.B2(n_79),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_71),
.B(n_55),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_71),
.B(n_55),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_181),
.B(n_186),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_109),
.B(n_51),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_132),
.A2(n_29),
.B1(n_49),
.B2(n_42),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_109),
.B(n_51),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_195),
.B(n_196),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_126),
.B(n_44),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_64),
.A2(n_70),
.B1(n_118),
.B2(n_81),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_202),
.A2(n_223),
.B1(n_43),
.B2(n_1),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_100),
.B(n_41),
.C(n_47),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_209),
.B(n_43),
.C(n_94),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_133),
.A2(n_42),
.B1(n_30),
.B2(n_31),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_211),
.A2(n_212),
.B1(n_221),
.B2(n_225),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_77),
.A2(n_42),
.B1(n_29),
.B2(n_49),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_119),
.B(n_41),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_219),
.B(n_230),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_91),
.A2(n_37),
.B1(n_31),
.B2(n_30),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_72),
.B(n_56),
.Y(n_222)
);

AND2x2_ASAP7_75t_SL g265 ( 
.A(n_222),
.B(n_0),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_87),
.A2(n_54),
.B1(n_37),
.B2(n_31),
.Y(n_223)
);

OA22x2_ASAP7_75t_L g224 ( 
.A1(n_90),
.A2(n_52),
.B1(n_37),
.B2(n_43),
.Y(n_224)
);

AO22x2_ASAP7_75t_L g255 ( 
.A1(n_224),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_255)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_95),
.Y(n_229)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_229),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_101),
.B(n_52),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_125),
.B(n_52),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_231),
.B(n_4),
.Y(n_289)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_106),
.Y(n_232)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_163),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_234),
.Y(n_367)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_235),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_236),
.A2(n_253),
.B1(n_263),
.B2(n_272),
.Y(n_353)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_239),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_240),
.Y(n_319)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_241),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_214),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_242),
.B(n_254),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_169),
.Y(n_243)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_243),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_150),
.B(n_121),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_244),
.Y(n_365)
);

BUFx4f_ASAP7_75t_SL g245 ( 
.A(n_214),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_245),
.Y(n_325)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_134),
.Y(n_246)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_246),
.Y(n_340)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_136),
.Y(n_247)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_247),
.Y(n_369)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_249),
.Y(n_366)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_250),
.Y(n_345)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_177),
.Y(n_252)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_252),
.Y(n_380)
);

AO21x2_ASAP7_75t_L g374 ( 
.A1(n_255),
.A2(n_275),
.B(n_283),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_224),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_256),
.A2(n_315),
.B1(n_317),
.B2(n_174),
.Y(n_356)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_226),
.Y(n_257)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_257),
.Y(n_321)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_197),
.Y(n_258)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_258),
.Y(n_324)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_180),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_259),
.Y(n_328)
);

BUFx8_ASAP7_75t_L g260 ( 
.A(n_214),
.Y(n_260)
);

INVx11_ASAP7_75t_L g348 ( 
.A(n_260),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_150),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_261),
.Y(n_381)
);

AOI222xp33_ASAP7_75t_L g262 ( 
.A1(n_145),
.A2(n_12),
.B1(n_18),
.B2(n_17),
.C1(n_16),
.C2(n_15),
.Y(n_262)
);

NOR3xp33_ASAP7_75t_L g349 ( 
.A(n_262),
.B(n_265),
.C(n_276),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_148),
.A2(n_12),
.B1(n_18),
.B2(n_17),
.Y(n_263)
);

OR2x2_ASAP7_75t_SL g266 ( 
.A(n_139),
.B(n_6),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_266),
.Y(n_344)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_216),
.Y(n_268)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_268),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_205),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_269),
.B(n_299),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_138),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_270),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_203),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_271),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_223),
.A2(n_6),
.B1(n_18),
.B2(n_17),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_167),
.A2(n_19),
.B1(n_16),
.B2(n_15),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_273),
.A2(n_298),
.B1(n_311),
.B2(n_204),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_210),
.A2(n_13),
.B1(n_1),
.B2(n_2),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_274),
.A2(n_287),
.B1(n_303),
.B2(n_304),
.Y(n_368)
);

OAI22xp33_ASAP7_75t_L g275 ( 
.A1(n_149),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_275)
);

NAND2x1_ASAP7_75t_SL g276 ( 
.A(n_200),
.B(n_3),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_138),
.Y(n_277)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_277),
.Y(n_331)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_197),
.Y(n_278)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_278),
.Y(n_358)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_203),
.Y(n_279)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_279),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_140),
.Y(n_281)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_281),
.Y(n_375)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_220),
.Y(n_282)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_282),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_165),
.A2(n_13),
.B1(n_4),
.B2(n_5),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_135),
.B(n_3),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_284),
.B(n_286),
.Y(n_339)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_217),
.Y(n_285)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_285),
.Y(n_379)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_183),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_224),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_289),
.B(n_290),
.Y(n_352)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_164),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_166),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_291),
.B(n_294),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_215),
.A2(n_4),
.B1(n_5),
.B2(n_193),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_292),
.A2(n_189),
.B(n_276),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_143),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_293),
.Y(n_326)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_190),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_176),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_295),
.B(n_296),
.Y(n_376)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_191),
.Y(n_296)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_140),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_297),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_142),
.A2(n_4),
.B1(n_160),
.B2(n_161),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_207),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_227),
.Y(n_300)
);

INVx11_ASAP7_75t_L g351 ( 
.A(n_300),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_147),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_301),
.Y(n_355)
);

NAND2x1_ASAP7_75t_L g302 ( 
.A(n_151),
.B(n_192),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_302),
.B(n_308),
.Y(n_342)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_227),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_226),
.Y(n_304)
);

INVx5_ASAP7_75t_L g306 ( 
.A(n_182),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_306),
.Y(n_360)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_168),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_310),
.Y(n_329)
);

NAND2x1_ASAP7_75t_L g308 ( 
.A(n_184),
.B(n_170),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_205),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_309),
.B(n_318),
.Y(n_332)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_198),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_171),
.A2(n_185),
.B1(n_204),
.B2(n_172),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_198),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_312),
.B(n_313),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_156),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_178),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_314),
.B(n_187),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_218),
.A2(n_228),
.B1(n_158),
.B2(n_173),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_206),
.B(n_194),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_316),
.B(n_185),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_159),
.A2(n_211),
.B1(n_188),
.B2(n_212),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_201),
.Y(n_318)
);

FAx1_ASAP7_75t_SL g320 ( 
.A(n_251),
.B(n_221),
.CI(n_146),
.CON(n_320),
.SN(n_320)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_320),
.B(n_341),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_SL g327 ( 
.A(n_233),
.B(n_182),
.C(n_146),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_327),
.B(n_361),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_330),
.A2(n_334),
.B1(n_306),
.B2(n_257),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_256),
.A2(n_171),
.B1(n_153),
.B2(n_168),
.Y(n_334)
);

O2A1O1Ixp33_ASAP7_75t_L g336 ( 
.A1(n_255),
.A2(n_141),
.B(n_175),
.C(n_201),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_336),
.A2(n_370),
.B(n_260),
.Y(n_410)
);

FAx1_ASAP7_75t_SL g341 ( 
.A(n_248),
.B(n_141),
.CI(n_175),
.CON(n_341),
.SN(n_341)
);

A2O1A1Ixp33_ASAP7_75t_L g354 ( 
.A1(n_264),
.A2(n_153),
.B(n_172),
.C(n_174),
.Y(n_354)
);

A2O1A1Ixp33_ASAP7_75t_L g416 ( 
.A1(n_354),
.A2(n_336),
.B(n_334),
.C(n_370),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_356),
.A2(n_245),
.B1(n_312),
.B2(n_310),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_362),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_265),
.B(n_187),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_363),
.B(n_373),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_364),
.Y(n_398)
);

O2A1O1Ixp33_ASAP7_75t_L g370 ( 
.A1(n_255),
.A2(n_189),
.B(n_305),
.C(n_240),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_317),
.A2(n_287),
.B(n_288),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_371),
.A2(n_275),
.B(n_242),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_284),
.B(n_280),
.Y(n_373)
);

OAI32xp33_ASAP7_75t_L g377 ( 
.A1(n_261),
.A2(n_267),
.A3(n_244),
.B1(n_266),
.B2(n_255),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_377),
.B(n_308),
.Y(n_384)
);

MAJx2_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_305),
.C(n_302),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_383),
.B(n_378),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_384),
.Y(n_434)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_362),
.Y(n_385)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_385),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_361),
.B(n_243),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_386),
.B(n_400),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_374),
.A2(n_315),
.B1(n_305),
.B2(n_274),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_387),
.A2(n_392),
.B1(n_404),
.B2(n_406),
.Y(n_436)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_359),
.Y(n_388)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_388),
.Y(n_437)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_333),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_390),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_352),
.B(n_271),
.Y(n_391)
);

INVxp33_ASAP7_75t_L g473 ( 
.A(n_391),
.Y(n_473)
);

OAI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_374),
.A2(n_303),
.B1(n_300),
.B2(n_239),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_359),
.Y(n_393)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_393),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_394),
.A2(n_410),
.B(n_321),
.Y(n_453)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_345),
.Y(n_395)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_395),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_323),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_396),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_397),
.A2(n_415),
.B1(n_360),
.B2(n_325),
.Y(n_440)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_319),
.A2(n_249),
.B1(n_268),
.B2(n_282),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_SL g454 ( 
.A1(n_399),
.A2(n_348),
.B1(n_347),
.B2(n_322),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_338),
.B(n_314),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_363),
.B(n_237),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_401),
.B(n_407),
.Y(n_441)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_333),
.Y(n_402)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_402),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_337),
.B(n_238),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_403),
.B(n_428),
.C(n_358),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_374),
.A2(n_297),
.B1(n_270),
.B2(n_277),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_376),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_405),
.B(n_408),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_374),
.A2(n_307),
.B1(n_281),
.B2(n_258),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_373),
.B(n_278),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_372),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_377),
.B(n_313),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_409),
.B(n_411),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_341),
.B(n_304),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_345),
.Y(n_412)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_412),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_413),
.A2(n_416),
.B1(n_417),
.B2(n_424),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_374),
.A2(n_245),
.B1(n_260),
.B2(n_371),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_319),
.A2(n_353),
.B1(n_368),
.B2(n_344),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_338),
.B(n_355),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_418),
.B(n_419),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_350),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_341),
.B(n_339),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_420),
.B(n_328),
.Y(n_468)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_379),
.Y(n_421)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_421),
.Y(n_451)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_335),
.Y(n_422)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_422),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_353),
.A2(n_337),
.B1(n_365),
.B2(n_320),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_342),
.A2(n_320),
.B1(n_364),
.B2(n_354),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_425),
.A2(n_430),
.B1(n_324),
.B2(n_369),
.Y(n_472)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_379),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_426),
.B(n_427),
.Y(n_459)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_335),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_342),
.B(n_340),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_340),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_429),
.B(n_395),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_330),
.A2(n_381),
.B1(n_327),
.B2(n_349),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_375),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_431),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_411),
.B(n_332),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_433),
.A2(n_462),
.B(n_441),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_409),
.A2(n_343),
.B1(n_381),
.B2(n_329),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_438),
.A2(n_455),
.B1(n_458),
.B2(n_416),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_440),
.A2(n_443),
.B1(n_463),
.B2(n_472),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_415),
.A2(n_329),
.B1(n_350),
.B2(n_375),
.Y(n_443)
);

XOR2x2_ASAP7_75t_L g444 ( 
.A(n_389),
.B(n_357),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_444),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_394),
.A2(n_321),
.B(n_326),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_449),
.A2(n_453),
.B(n_410),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_452),
.B(n_466),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_454),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_384),
.A2(n_331),
.B1(n_346),
.B2(n_378),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_367),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_456),
.B(n_469),
.C(n_383),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_420),
.A2(n_331),
.B1(n_346),
.B2(n_322),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_414),
.A2(n_358),
.B(n_347),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_406),
.A2(n_351),
.B1(n_323),
.B2(n_366),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_464),
.B(n_471),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_465),
.B(n_456),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_389),
.B(n_380),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_468),
.B(n_470),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_403),
.B(n_328),
.C(n_380),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_385),
.B(n_366),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_474),
.A2(n_491),
.B1(n_506),
.B2(n_432),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_475),
.B(n_494),
.Y(n_522)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_459),
.Y(n_477)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_477),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_445),
.B(n_423),
.Y(n_478)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_478),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_459),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_480),
.B(n_508),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_481),
.A2(n_489),
.B(n_462),
.Y(n_526)
);

INVx13_ASAP7_75t_L g482 ( 
.A(n_435),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_482),
.Y(n_534)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_464),
.Y(n_483)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_483),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_445),
.B(n_473),
.Y(n_484)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_484),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_467),
.A2(n_413),
.B1(n_398),
.B2(n_387),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_485),
.A2(n_492),
.B1(n_496),
.B2(n_511),
.Y(n_528)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_437),
.Y(n_486)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_486),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_471),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_487),
.B(n_500),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_453),
.A2(n_414),
.B(n_425),
.Y(n_489)
);

CKINVDCx14_ASAP7_75t_R g529 ( 
.A(n_490),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_436),
.A2(n_382),
.B1(n_423),
.B2(n_391),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_467),
.A2(n_424),
.B1(n_416),
.B2(n_404),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_436),
.A2(n_383),
.B1(n_386),
.B2(n_382),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_444),
.B(n_407),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_497),
.B(n_503),
.C(n_466),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_442),
.B(n_418),
.Y(n_498)
);

NAND3xp33_ASAP7_75t_L g531 ( 
.A(n_498),
.B(n_451),
.C(n_450),
.Y(n_531)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_437),
.Y(n_499)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_499),
.Y(n_551)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_439),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_461),
.Y(n_501)
);

OAI21xp33_ASAP7_75t_SL g546 ( 
.A1(n_501),
.A2(n_504),
.B(n_506),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_502),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_465),
.B(n_417),
.C(n_401),
.Y(n_503)
);

OA22x2_ASAP7_75t_L g504 ( 
.A1(n_472),
.A2(n_430),
.B1(n_412),
.B2(n_431),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_439),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_505),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_455),
.A2(n_429),
.B1(n_427),
.B2(n_393),
.Y(n_506)
);

MAJx2_ASAP7_75t_L g507 ( 
.A(n_444),
.B(n_388),
.C(n_421),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_507),
.B(n_452),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_442),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_466),
.B(n_426),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_509),
.B(n_495),
.Y(n_530)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_447),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_510),
.B(n_446),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_434),
.A2(n_390),
.B1(n_402),
.B2(n_422),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_432),
.B(n_441),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_512),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_460),
.A2(n_400),
.B1(n_396),
.B2(n_324),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_513),
.A2(n_463),
.B1(n_461),
.B2(n_457),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_474),
.A2(n_460),
.B1(n_449),
.B2(n_433),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_515),
.A2(n_538),
.B1(n_545),
.B2(n_535),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_SL g578 ( 
.A(n_516),
.B(n_348),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_517),
.B(n_530),
.Y(n_554)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_518),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_519),
.A2(n_523),
.B1(n_531),
.B2(n_540),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_475),
.B(n_468),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_521),
.B(n_537),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_479),
.A2(n_433),
.B1(n_440),
.B2(n_443),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_SL g524 ( 
.A(n_496),
.B(n_489),
.C(n_485),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_524),
.B(n_527),
.C(n_549),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_526),
.A2(n_513),
.B(n_488),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_494),
.B(n_469),
.C(n_470),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_484),
.B(n_458),
.Y(n_532)
);

CKINVDCx14_ASAP7_75t_R g559 ( 
.A(n_532),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_477),
.B(n_438),
.Y(n_533)
);

INVxp33_ASAP7_75t_SL g581 ( 
.A(n_533),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_495),
.B(n_451),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_481),
.A2(n_450),
.B1(n_447),
.B2(n_454),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_483),
.B(n_396),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g574 ( 
.A(n_543),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_492),
.A2(n_435),
.B1(n_461),
.B2(n_448),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_544),
.B(n_546),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_487),
.A2(n_512),
.B1(n_502),
.B2(n_478),
.Y(n_548)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_548),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_503),
.B(n_448),
.C(n_457),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_509),
.B(n_369),
.C(n_351),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_550),
.B(n_511),
.C(n_500),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_521),
.Y(n_552)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_552),
.Y(n_586)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_541),
.Y(n_553)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_553),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_555),
.A2(n_568),
.B(n_565),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_L g558 ( 
.A1(n_514),
.A2(n_526),
.B(n_515),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_558),
.Y(n_594)
);

XOR2x2_ASAP7_75t_L g561 ( 
.A(n_516),
.B(n_497),
.Y(n_561)
);

MAJx2_ASAP7_75t_L g587 ( 
.A(n_561),
.B(n_578),
.C(n_530),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_520),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_563),
.B(n_567),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_564),
.B(n_573),
.C(n_580),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_528),
.A2(n_493),
.B1(n_488),
.B2(n_476),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_565),
.A2(n_566),
.B1(n_575),
.B2(n_545),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_528),
.A2(n_493),
.B1(n_476),
.B2(n_504),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_520),
.Y(n_567)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_567),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_522),
.B(n_507),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_569),
.B(n_571),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_SL g570 ( 
.A1(n_538),
.A2(n_501),
.B1(n_510),
.B2(n_486),
.Y(n_570)
);

OAI22xp33_ASAP7_75t_SL g584 ( 
.A1(n_570),
.A2(n_540),
.B1(n_544),
.B2(n_534),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_522),
.B(n_504),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_525),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_572),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_549),
.B(n_504),
.C(n_499),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_535),
.A2(n_505),
.B1(n_501),
.B2(n_482),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_525),
.Y(n_576)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_576),
.Y(n_607)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_542),
.Y(n_577)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_577),
.Y(n_595)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_542),
.Y(n_579)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_579),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_582),
.A2(n_539),
.B1(n_529),
.B2(n_536),
.Y(n_593)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_547),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_583),
.B(n_551),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_584),
.Y(n_628)
);

FAx1_ASAP7_75t_L g585 ( 
.A(n_558),
.B(n_524),
.CI(n_539),
.CON(n_585),
.SN(n_585)
);

A2O1A1Ixp33_ASAP7_75t_SL g616 ( 
.A1(n_585),
.A2(n_562),
.B(n_578),
.C(n_569),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_587),
.B(n_589),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_SL g614 ( 
.A1(n_588),
.A2(n_599),
.B1(n_555),
.B2(n_568),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_562),
.B(n_527),
.C(n_517),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_590),
.B(n_606),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_592),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_593),
.A2(n_585),
.B1(n_594),
.B2(n_602),
.Y(n_626)
);

AOI211xp5_ASAP7_75t_SL g596 ( 
.A1(n_582),
.A2(n_550),
.B(n_534),
.C(n_537),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_596),
.A2(n_573),
.B(n_568),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_557),
.A2(n_547),
.B1(n_551),
.B2(n_560),
.Y(n_599)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_600),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_L g617 ( 
.A1(n_601),
.A2(n_553),
.B(n_583),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_556),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_603),
.B(n_574),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_564),
.Y(n_604)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_604),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_572),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g608 ( 
.A(n_554),
.B(n_571),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_608),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_575),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_609),
.B(n_595),
.Y(n_631)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_610),
.B(n_626),
.Y(n_639)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_613),
.Y(n_633)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_614),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_SL g615 ( 
.A1(n_588),
.A2(n_581),
.B1(n_559),
.B2(n_566),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_615),
.A2(n_629),
.B1(n_605),
.B2(n_607),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_616),
.B(n_622),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_617),
.A2(n_630),
.B(n_613),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_604),
.B(n_554),
.C(n_580),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_621),
.Y(n_637)
);

FAx1_ASAP7_75t_SL g622 ( 
.A(n_585),
.B(n_561),
.CI(n_587),
.CON(n_622),
.SN(n_622)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_589),
.B(n_590),
.C(n_608),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_623),
.B(n_627),
.C(n_591),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_593),
.B(n_592),
.Y(n_624)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_624),
.Y(n_634)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_626),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_598),
.B(n_594),
.C(n_586),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_599),
.A2(n_601),
.B1(n_597),
.B2(n_596),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_598),
.A2(n_595),
.B(n_605),
.Y(n_630)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_631),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_632),
.B(n_635),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_623),
.B(n_625),
.C(n_611),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_638),
.B(n_642),
.Y(n_663)
);

XNOR2xp5_ASAP7_75t_SL g662 ( 
.A(n_639),
.B(n_643),
.Y(n_662)
);

CKINVDCx14_ASAP7_75t_R g640 ( 
.A(n_620),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_640),
.B(n_616),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_SL g641 ( 
.A1(n_628),
.A2(n_614),
.B1(n_615),
.B2(n_624),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_641),
.B(n_616),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_625),
.B(n_627),
.Y(n_642)
);

XOR2xp5_ASAP7_75t_L g643 ( 
.A(n_610),
.B(n_629),
.Y(n_643)
);

XOR2xp5_ASAP7_75t_L g653 ( 
.A(n_643),
.B(n_647),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_628),
.A2(n_612),
.B1(n_617),
.B2(n_618),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_SL g655 ( 
.A1(n_645),
.A2(n_622),
.B1(n_616),
.B2(n_619),
.Y(n_655)
);

XOR2xp5_ASAP7_75t_L g647 ( 
.A(n_630),
.B(n_619),
.Y(n_647)
);

AOI21x1_ASAP7_75t_L g654 ( 
.A1(n_649),
.A2(n_612),
.B(n_622),
.Y(n_654)
);

INVxp67_ASAP7_75t_SL g651 ( 
.A(n_635),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_651),
.B(n_652),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_637),
.B(n_618),
.Y(n_652)
);

INVxp67_ASAP7_75t_SL g666 ( 
.A(n_654),
.Y(n_666)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_655),
.B(n_656),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_648),
.B(n_621),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_657),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_SL g658 ( 
.A(n_638),
.B(n_616),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_658),
.B(n_660),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_659),
.B(n_656),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g660 ( 
.A(n_647),
.B(n_636),
.C(n_639),
.Y(n_660)
);

INVx11_ASAP7_75t_L g661 ( 
.A(n_649),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g667 ( 
.A1(n_661),
.A2(n_646),
.B1(n_641),
.B2(n_644),
.Y(n_667)
);

XOR2xp5_ASAP7_75t_L g674 ( 
.A(n_662),
.B(n_653),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_645),
.B(n_633),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_664),
.B(n_634),
.Y(n_665)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_665),
.Y(n_677)
);

AOI21x1_ASAP7_75t_L g678 ( 
.A1(n_667),
.A2(n_660),
.B(n_650),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_661),
.A2(n_636),
.B1(n_632),
.B2(n_646),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_670),
.B(n_672),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_674),
.A2(n_654),
.B(n_653),
.Y(n_681)
);

OAI21xp5_ASAP7_75t_SL g675 ( 
.A1(n_671),
.A2(n_673),
.B(n_669),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_SL g685 ( 
.A(n_675),
.B(n_655),
.Y(n_685)
);

OAI21x1_ASAP7_75t_SL g683 ( 
.A1(n_678),
.A2(n_679),
.B(n_681),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_666),
.B(n_663),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_666),
.B(n_657),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_680),
.B(n_668),
.Y(n_682)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_682),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_L g684 ( 
.A1(n_679),
.A2(n_668),
.B(n_672),
.Y(n_684)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_684),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_686),
.B(n_677),
.Y(n_688)
);

BUFx24_ASAP7_75t_SL g689 ( 
.A(n_688),
.Y(n_689)
);

O2A1O1Ixp33_ASAP7_75t_SL g690 ( 
.A1(n_689),
.A2(n_687),
.B(n_683),
.C(n_685),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_690),
.A2(n_676),
.B(n_662),
.Y(n_691)
);


endmodule