module fake_jpeg_20714_n_48 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_48);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_48;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx5_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx4f_ASAP7_75t_SL g11 ( 
.A(n_1),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_22),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_17),
.A2(n_3),
.B1(n_4),
.B2(n_13),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g18 ( 
.A(n_15),
.B(n_2),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_20),
.C(n_9),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_7),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_19)
);

AO22x1_ASAP7_75t_L g32 ( 
.A1(n_19),
.A2(n_21),
.B1(n_8),
.B2(n_11),
.Y(n_32)
);

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_8),
.B(n_3),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_18),
.B(n_14),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_32),
.B1(n_30),
.B2(n_27),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_19),
.A2(n_21),
.B1(n_20),
.B2(n_23),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_19),
.B1(n_24),
.B2(n_25),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_13),
.B(n_32),
.C(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_11),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_18),
.C(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_37),
.Y(n_41)
);

AO21x1_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_37),
.B(n_35),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_36),
.A2(n_26),
.B1(n_33),
.B2(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_35),
.B(n_27),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_44),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_SL g46 ( 
.A1(n_45),
.A2(n_36),
.B(n_39),
.C(n_42),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_40),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_41),
.C(n_43),
.Y(n_48)
);


endmodule