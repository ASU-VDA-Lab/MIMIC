module fake_jpeg_17358_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx24_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_7),
.Y(n_39)
);

NAND3xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_24),
.C(n_30),
.Y(n_49)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_25),
.B1(n_27),
.B2(n_21),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_41),
.A2(n_56),
.B1(n_34),
.B2(n_20),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_42),
.A2(n_52),
.B1(n_54),
.B2(n_57),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_30),
.CON(n_43),
.SN(n_43)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_43),
.A2(n_49),
.B(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_29),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_50),
.Y(n_82)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_29),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_25),
.B1(n_28),
.B2(n_24),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_54)
);

NAND2x1p5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_16),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_34),
.A2(n_27),
.B1(n_31),
.B2(n_21),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_63),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_39),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_66),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_52),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_71),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_38),
.C(n_36),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_36),
.C(n_35),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_53),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_76),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_53),
.B(n_32),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_48),
.A2(n_20),
.B1(n_40),
.B2(n_17),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_88),
.B1(n_16),
.B2(n_23),
.Y(n_100)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_19),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_84),
.Y(n_97)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

CKINVDCx9p33_ASAP7_75t_R g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_35),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

AOI32xp33_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_42),
.A3(n_54),
.B1(n_36),
.B2(n_40),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_89),
.A2(n_95),
.B(n_82),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_35),
.B1(n_17),
.B2(n_23),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_92),
.A2(n_98),
.B1(n_106),
.B2(n_114),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_96),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_35),
.Y(n_96)
);

AO22x2_ASAP7_75t_L g98 ( 
.A1(n_69),
.A2(n_36),
.B1(n_23),
.B2(n_17),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

AO22x2_ASAP7_75t_SL g106 ( 
.A1(n_72),
.A2(n_23),
.B1(n_18),
.B2(n_16),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_18),
.B1(n_26),
.B2(n_16),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_SL g116 ( 
.A1(n_98),
.A2(n_106),
.B(n_94),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_98),
.C(n_106),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_113),
.A2(n_75),
.B1(n_82),
.B2(n_70),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_117),
.A2(n_132),
.B1(n_106),
.B2(n_105),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_65),
.Y(n_119)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_77),
.B(n_75),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_97),
.B(n_109),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_91),
.Y(n_156)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_66),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_128),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_129),
.Y(n_159)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_68),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_101),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_133),
.Y(n_169)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_110),
.A2(n_76),
.B1(n_73),
.B2(n_74),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_101),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_78),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_138),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_85),
.Y(n_135)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_83),
.Y(n_136)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_90),
.B(n_79),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_139),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_59),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_141),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_93),
.B(n_26),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_59),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_143),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_144),
.B(n_156),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_126),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_102),
.B1(n_97),
.B2(n_114),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_SL g182 ( 
.A1(n_146),
.A2(n_157),
.B(n_163),
.C(n_137),
.Y(n_182)
);

NOR2xp67_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_102),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_149),
.A2(n_151),
.B(n_118),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_109),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_158),
.C(n_117),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_91),
.A3(n_26),
.B1(n_115),
.B2(n_18),
.C1(n_61),
.C2(n_19),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_119),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_61),
.B1(n_62),
.B2(n_112),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_112),
.C(n_19),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_167),
.Y(n_186)
);

AO22x1_ASAP7_75t_L g163 ( 
.A1(n_116),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_129),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_133),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_174),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_117),
.C(n_124),
.Y(n_174)
);

NAND2xp33_ASAP7_75t_SL g175 ( 
.A(n_151),
.B(n_120),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_176),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_131),
.C(n_140),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_178),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_180),
.A2(n_182),
.B1(n_188),
.B2(n_189),
.Y(n_206)
);

BUFx12f_ASAP7_75t_SL g181 ( 
.A(n_163),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_181),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_138),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_183),
.B(n_184),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_132),
.C(n_136),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_132),
.C(n_128),
.Y(n_187)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_165),
.A2(n_126),
.B1(n_142),
.B2(n_141),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_190),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_135),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_191),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_192),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_134),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_146),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_148),
.B(n_126),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_148),
.B(n_19),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_166),
.B1(n_144),
.B2(n_172),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_197),
.A2(n_200),
.B1(n_204),
.B2(n_212),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_181),
.A2(n_172),
.B1(n_147),
.B2(n_155),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_187),
.A2(n_160),
.B1(n_145),
.B2(n_155),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_207),
.B(n_193),
.Y(n_220)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_201),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_174),
.A2(n_160),
.B1(n_164),
.B2(n_163),
.Y(n_212)
);

XOR2x2_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_164),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_213),
.B(n_196),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_219),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_173),
.C(n_177),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_222),
.C(n_226),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_184),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_220),
.B(n_221),
.Y(n_233)
);

AOI21xp33_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_182),
.B(n_178),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_182),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_210),
.A2(n_182),
.B1(n_167),
.B2(n_170),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_223),
.B(n_228),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_211),
.B(n_161),
.Y(n_224)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

AOI321xp33_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_162),
.A3(n_8),
.B1(n_9),
.B2(n_4),
.C(n_5),
.Y(n_225)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_7),
.Y(n_226)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_203),
.B(n_7),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_210),
.A2(n_8),
.B(n_14),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_229),
.B(n_230),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_215),
.B(n_6),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_214),
.C(n_198),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_242),
.C(n_232),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_198),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_239),
.B(n_240),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_212),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_208),
.C(n_200),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_222),
.B(n_226),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_249),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_209),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_248),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_250),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_197),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_251),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_231),
.B(n_202),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_229),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_235),
.B(n_205),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_205),
.B(n_10),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_0),
.C(n_2),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_3),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_246),
.A2(n_236),
.B1(n_241),
.B2(n_5),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_259),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_3),
.Y(n_261)
);

NOR2x1_ASAP7_75t_SL g259 ( 
.A(n_252),
.B(n_241),
.Y(n_259)
);

AOI322xp5_ASAP7_75t_L g267 ( 
.A1(n_261),
.A2(n_264),
.A3(n_6),
.B1(n_10),
.B2(n_11),
.C1(n_13),
.C2(n_14),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_247),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_6),
.B(n_10),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_245),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_253),
.C(n_256),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_4),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_265),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_266),
.A2(n_267),
.B1(n_260),
.B2(n_15),
.Y(n_269)
);

OAI21x1_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_262),
.B(n_13),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_270),
.B(n_15),
.Y(n_271)
);

NAND2x1p5_ASAP7_75t_SL g272 ( 
.A(n_271),
.B(n_268),
.Y(n_272)
);


endmodule