module real_jpeg_6891_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_1),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_1),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_1),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_1),
.Y(n_206)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_1),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_1),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_2),
.Y(n_83)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_2),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_3),
.A2(n_96),
.B1(n_98),
.B2(n_102),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_3),
.Y(n_102)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_5),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_5),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_5),
.Y(n_156)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_5),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_6),
.A2(n_119),
.B1(n_130),
.B2(n_133),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_6),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_6),
.A2(n_133),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_6),
.A2(n_133),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_7),
.A2(n_189),
.B1(n_192),
.B2(n_193),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_7),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_8),
.Y(n_79)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_8),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_8),
.Y(n_209)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_10),
.A2(n_36),
.B1(n_40),
.B2(n_43),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_10),
.A2(n_43),
.B1(n_136),
.B2(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_10),
.A2(n_43),
.B1(n_282),
.B2(n_284),
.Y(n_281)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_11),
.B(n_146),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_11),
.A2(n_71),
.B1(n_247),
.B2(n_249),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_11),
.B(n_122),
.C(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_11),
.B(n_24),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_11),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_11),
.B(n_138),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_12),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_12),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_12),
.A2(n_84),
.B1(n_232),
.B2(n_235),
.Y(n_231)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_13),
.Y(n_114)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_13),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_13),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_14),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_14),
.A2(n_50),
.B1(n_120),
.B2(n_136),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_14),
.A2(n_50),
.B1(n_92),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_14),
.A2(n_50),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_240),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_238),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_160),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_19),
.B(n_160),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_105),
.C(n_139),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_20),
.A2(n_21),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_69),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_22),
.B(n_70),
.C(n_80),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_35),
.B(n_44),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_23),
.A2(n_35),
.B1(n_55),
.B2(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_23),
.B(n_46),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_24),
.B(n_56),
.Y(n_55)
);

AO22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B1(n_30),
.B2(n_32),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_26),
.Y(n_153)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_28),
.Y(n_235)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_29),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_29),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_31),
.Y(n_137)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_31),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_31),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_31),
.Y(n_253)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g224 ( 
.A(n_37),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_38),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g312 ( 
.A(n_38),
.Y(n_312)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_39),
.Y(n_176)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_54),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_49),
.Y(n_141)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_54),
.A2(n_311),
.B(n_314),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_60),
.B1(n_63),
.B2(n_65),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_59),
.Y(n_144)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_62),
.Y(n_228)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_80),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_71),
.B(n_178),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_SL g210 ( 
.A1(n_71),
.A2(n_177),
.B(n_211),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_71),
.A2(n_181),
.B(n_263),
.Y(n_278)
);

OAI21xp33_ASAP7_75t_SL g311 ( 
.A1(n_71),
.A2(n_312),
.B(n_313),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_72),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_72),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_78),
.Y(n_72)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_73),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g164 ( 
.A1(n_75),
.A2(n_165),
.A3(n_169),
.B1(n_171),
.B2(n_177),
.Y(n_164)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_79),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_90),
.B1(n_95),
.B2(n_103),
.Y(n_80)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_81),
.Y(n_155)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_83),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_83),
.Y(n_255)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_83),
.Y(n_286)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_88),
.Y(n_262)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_88),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_90),
.B(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_90),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_90),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_91),
.Y(n_298)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_95),
.Y(n_182)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_122),
.B1(n_124),
.B2(n_127),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_100),
.Y(n_193)
);

BUFx8_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_104),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_105),
.B(n_139),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_129),
.B(n_134),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_106),
.A2(n_134),
.B(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_106),
.A2(n_129),
.B1(n_230),
.B2(n_268),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_107),
.B(n_135),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_121),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_112),
.B1(n_115),
.B2(n_119),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_121),
.A2(n_236),
.B(n_268),
.Y(n_267)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

INVx3_ASAP7_75t_SL g142 ( 
.A(n_136),
.Y(n_142)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_138),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_154),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_140),
.B(n_154),
.Y(n_315)
);

AOI32xp33_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.A3(n_143),
.B1(n_145),
.B2(n_148),
.Y(n_140)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp33_ASAP7_75t_L g313 ( 
.A(n_145),
.Y(n_313)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp33_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B(n_157),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_157),
.A2(n_281),
.B(n_287),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_158),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_159),
.B(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_197),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_161)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_179),
.B2(n_180),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

INVx6_ASAP7_75t_SL g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_187),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_181),
.A2(n_258),
.B(n_263),
.Y(n_257)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_186),
.Y(n_277)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_186),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_194),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_220),
.B2(n_237),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_210),
.B(n_213),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_201)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_211),
.Y(n_218)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_229),
.Y(n_220)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B(n_236),
.Y(n_229)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_235),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

AO21x1_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_317),
.B(n_322),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_303),
.B(n_316),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_272),
.B(n_302),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_256),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_244),
.B(n_256),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_251),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_245),
.A2(n_251),
.B1(n_252),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_245),
.Y(n_300)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_265),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_257),
.B(n_266),
.C(n_271),
.Y(n_304)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_258),
.Y(n_295)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_270),
.B2(n_271),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_292),
.B(n_301),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_279),
.B(n_291),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_290),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_290),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_299),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_299),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_297),
.Y(n_296)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_305),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_315),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_309),
.C(n_315),
.Y(n_318)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_318),
.B(n_319),
.Y(n_322)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);


endmodule