module fake_netlist_1_4520_n_498 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_498);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_498;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_486;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g66 ( .A(n_64), .Y(n_66) );
INVx1_ASAP7_75t_L g67 ( .A(n_60), .Y(n_67) );
CKINVDCx5p33_ASAP7_75t_R g68 ( .A(n_12), .Y(n_68) );
INVx1_ASAP7_75t_L g69 ( .A(n_5), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_13), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_22), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_26), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_28), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_34), .Y(n_74) );
INVxp33_ASAP7_75t_L g75 ( .A(n_51), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_52), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_54), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_29), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_61), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_3), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_46), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_25), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_43), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_9), .Y(n_84) );
INVx1_ASAP7_75t_SL g85 ( .A(n_37), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_10), .Y(n_86) );
INVx1_ASAP7_75t_SL g87 ( .A(n_12), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_65), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_38), .Y(n_89) );
INVxp33_ASAP7_75t_L g90 ( .A(n_30), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_15), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_23), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_11), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_8), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_48), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_11), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_17), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_5), .Y(n_98) );
BUFx2_ASAP7_75t_L g99 ( .A(n_6), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_44), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_4), .Y(n_101) );
CKINVDCx14_ASAP7_75t_R g102 ( .A(n_36), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_62), .Y(n_103) );
AND2x2_ASAP7_75t_L g104 ( .A(n_99), .B(n_0), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_89), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_89), .Y(n_106) );
AND2x4_ASAP7_75t_L g107 ( .A(n_69), .B(n_0), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_67), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_67), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_71), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_100), .Y(n_111) );
AND2x4_ASAP7_75t_L g112 ( .A(n_69), .B(n_1), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_71), .Y(n_113) );
INVx3_ASAP7_75t_L g114 ( .A(n_72), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_72), .Y(n_115) );
BUFx3_ASAP7_75t_L g116 ( .A(n_100), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_73), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_73), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_99), .B(n_1), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_66), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_74), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_74), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_76), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_76), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_118), .Y(n_125) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_104), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_120), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_118), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_118), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_104), .B(n_102), .Y(n_130) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_104), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_118), .Y(n_132) );
OR2x2_ASAP7_75t_SL g133 ( .A(n_108), .B(n_80), .Y(n_133) );
INVxp67_ASAP7_75t_L g134 ( .A(n_119), .Y(n_134) );
INVx8_ASAP7_75t_L g135 ( .A(n_107), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_107), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_118), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_118), .Y(n_138) );
AOI22xp33_ASAP7_75t_L g139 ( .A1(n_107), .A2(n_84), .B1(n_101), .B2(n_91), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_107), .B(n_70), .Y(n_140) );
INVx4_ASAP7_75t_L g141 ( .A(n_107), .Y(n_141) );
BUFx10_ASAP7_75t_L g142 ( .A(n_112), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_108), .B(n_75), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_121), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_119), .B(n_90), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_119), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_121), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_137), .Y(n_148) );
INVx4_ASAP7_75t_L g149 ( .A(n_135), .Y(n_149) );
BUFx3_ASAP7_75t_L g150 ( .A(n_135), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_134), .B(n_112), .Y(n_151) );
CKINVDCx6p67_ASAP7_75t_R g152 ( .A(n_126), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_136), .Y(n_153) );
NAND2x1p5_ASAP7_75t_L g154 ( .A(n_141), .B(n_112), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_137), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_141), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_145), .B(n_114), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_136), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_136), .Y(n_159) );
BUFx3_ASAP7_75t_L g160 ( .A(n_135), .Y(n_160) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_135), .A2(n_112), .B1(n_123), .B2(n_122), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_136), .Y(n_162) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_131), .Y(n_163) );
OR2x6_ASAP7_75t_L g164 ( .A(n_135), .B(n_112), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_135), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_145), .B(n_114), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_137), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_141), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_134), .B(n_114), .Y(n_169) );
BUFx4f_ASAP7_75t_L g170 ( .A(n_140), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_130), .B(n_109), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_141), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_137), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_137), .Y(n_174) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_131), .Y(n_175) );
OR2x2_ASAP7_75t_L g176 ( .A(n_126), .B(n_87), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_140), .A2(n_109), .B1(n_123), .B2(n_122), .Y(n_177) );
INVx4_ASAP7_75t_L g178 ( .A(n_142), .Y(n_178) );
NOR2xp67_ASAP7_75t_SL g179 ( .A(n_149), .B(n_142), .Y(n_179) );
INVx2_ASAP7_75t_SL g180 ( .A(n_150), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_168), .Y(n_181) );
INVxp67_ASAP7_75t_SL g182 ( .A(n_150), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_168), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_149), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_177), .B(n_146), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_149), .B(n_146), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_153), .A2(n_140), .B(n_130), .Y(n_187) );
INVx8_ASAP7_75t_L g188 ( .A(n_164), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_149), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_150), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_160), .B(n_140), .Y(n_191) );
CKINVDCx11_ASAP7_75t_R g192 ( .A(n_152), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_172), .Y(n_193) );
INVx5_ASAP7_75t_L g194 ( .A(n_178), .Y(n_194) );
BUFx2_ASAP7_75t_L g195 ( .A(n_160), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_172), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_163), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_178), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_153), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_163), .Y(n_200) );
INVx3_ASAP7_75t_SL g201 ( .A(n_152), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_177), .B(n_143), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_151), .B(n_139), .Y(n_203) );
INVx5_ASAP7_75t_L g204 ( .A(n_178), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_151), .B(n_142), .Y(n_205) );
INVx1_ASAP7_75t_SL g206 ( .A(n_152), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_175), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_151), .B(n_142), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_151), .B(n_110), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_186), .A2(n_170), .B1(n_175), .B2(n_176), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_202), .A2(n_185), .B1(n_161), .B2(n_203), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_199), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_186), .A2(n_170), .B1(n_176), .B2(n_151), .Y(n_213) );
NAND2x1p5_ASAP7_75t_L g214 ( .A(n_194), .B(n_160), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_192), .Y(n_215) );
CKINVDCx6p67_ASAP7_75t_R g216 ( .A(n_201), .Y(n_216) );
OAI22xp5_ASAP7_75t_SL g217 ( .A1(n_201), .A2(n_133), .B1(n_127), .B2(n_176), .Y(n_217) );
XNOR2x1_ASAP7_75t_L g218 ( .A(n_186), .B(n_154), .Y(n_218) );
HB1xp67_ASAP7_75t_L g219 ( .A(n_206), .Y(n_219) );
OAI22xp5_ASAP7_75t_SL g220 ( .A1(n_197), .A2(n_133), .B1(n_96), .B2(n_86), .Y(n_220) );
BUFx2_ASAP7_75t_L g221 ( .A(n_188), .Y(n_221) );
AOI22xp33_ASAP7_75t_SL g222 ( .A1(n_188), .A2(n_170), .B1(n_165), .B2(n_166), .Y(n_222) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_209), .A2(n_161), .B1(n_170), .B2(n_164), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_199), .Y(n_224) );
AOI21xp33_ASAP7_75t_L g225 ( .A1(n_180), .A2(n_157), .B(n_166), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_184), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_184), .Y(n_227) );
OAI21x1_ASAP7_75t_L g228 ( .A1(n_187), .A2(n_148), .B(n_174), .Y(n_228) );
AOI222xp33_ASAP7_75t_L g229 ( .A1(n_200), .A2(n_171), .B1(n_157), .B2(n_169), .C1(n_70), .C2(n_91), .Y(n_229) );
OAI21x1_ASAP7_75t_L g230 ( .A1(n_198), .A2(n_167), .B(n_174), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_181), .Y(n_231) );
OAI222xp33_ASAP7_75t_L g232 ( .A1(n_207), .A2(n_68), .B1(n_164), .B2(n_101), .C1(n_84), .C2(n_93), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_184), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_183), .B(n_169), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_193), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_217), .A2(n_192), .B1(n_188), .B2(n_191), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_224), .Y(n_237) );
OAI21xp33_ASAP7_75t_L g238 ( .A1(n_218), .A2(n_116), .B(n_117), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_218), .B(n_164), .Y(n_239) );
AOI22xp33_ASAP7_75t_SL g240 ( .A1(n_218), .A2(n_188), .B1(n_195), .B2(n_204), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_229), .B(n_196), .Y(n_241) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_228), .A2(n_111), .B(n_105), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_224), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_217), .A2(n_191), .B1(n_195), .B2(n_190), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_223), .A2(n_191), .B1(n_190), .B2(n_164), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_224), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_212), .Y(n_247) );
BUFx6f_ASAP7_75t_SL g248 ( .A(n_216), .Y(n_248) );
NAND3xp33_ASAP7_75t_L g249 ( .A(n_223), .B(n_121), .C(n_124), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_222), .A2(n_164), .B1(n_182), .B2(n_154), .Y(n_250) );
OAI21xp33_ASAP7_75t_L g251 ( .A1(n_213), .A2(n_116), .B(n_117), .Y(n_251) );
INVxp67_ASAP7_75t_L g252 ( .A(n_219), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_212), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_230), .Y(n_254) );
INVx2_ASAP7_75t_SL g255 ( .A(n_214), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_230), .Y(n_256) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_254), .Y(n_257) );
AOI221xp5_ASAP7_75t_L g258 ( .A1(n_241), .A2(n_220), .B1(n_211), .B2(n_232), .C(n_210), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_246), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_246), .B(n_228), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_246), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_237), .Y(n_262) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_237), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_243), .B(n_226), .Y(n_264) );
NOR3xp33_ASAP7_75t_L g265 ( .A(n_238), .B(n_220), .C(n_225), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_243), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_254), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_254), .Y(n_268) );
OA21x2_ASAP7_75t_L g269 ( .A1(n_256), .A2(n_228), .B(n_230), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_247), .Y(n_270) );
AO21x2_ASAP7_75t_L g271 ( .A1(n_249), .A2(n_225), .B(n_233), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_247), .B(n_231), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_256), .A2(n_226), .B(n_227), .Y(n_273) );
OAI33xp33_ASAP7_75t_L g274 ( .A1(n_252), .A2(n_77), .A3(n_79), .B1(n_81), .B2(n_82), .B3(n_83), .Y(n_274) );
AOI21x1_ASAP7_75t_L g275 ( .A1(n_256), .A2(n_233), .B(n_226), .Y(n_275) );
AOI31xp33_ASAP7_75t_L g276 ( .A1(n_240), .A2(n_215), .A3(n_214), .B(n_216), .Y(n_276) );
NOR2x1_ASAP7_75t_L g277 ( .A(n_276), .B(n_249), .Y(n_277) );
OAI31xp33_ASAP7_75t_SL g278 ( .A1(n_258), .A2(n_238), .A3(n_250), .B(n_239), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_263), .Y(n_279) );
OAI33xp33_ASAP7_75t_L g280 ( .A1(n_270), .A2(n_97), .A3(n_94), .B1(n_98), .B2(n_77), .B3(n_79), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_261), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_270), .Y(n_282) );
INVx4_ASAP7_75t_L g283 ( .A(n_259), .Y(n_283) );
OAI33xp33_ASAP7_75t_L g284 ( .A1(n_272), .A2(n_103), .A3(n_82), .B1(n_83), .B2(n_92), .B3(n_81), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_258), .A2(n_239), .B1(n_245), .B2(n_236), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_272), .B(n_253), .Y(n_286) );
OAI33xp33_ASAP7_75t_L g287 ( .A1(n_262), .A2(n_103), .A3(n_92), .B1(n_95), .B2(n_115), .B3(n_110), .Y(n_287) );
NAND3xp33_ASAP7_75t_L g288 ( .A(n_265), .B(n_244), .C(n_124), .Y(n_288) );
OAI21xp33_ASAP7_75t_L g289 ( .A1(n_276), .A2(n_116), .B(n_105), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_265), .A2(n_253), .B1(n_248), .B2(n_251), .Y(n_290) );
AOI21xp5_ASAP7_75t_SL g291 ( .A1(n_260), .A2(n_255), .B(n_248), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_274), .A2(n_235), .B1(n_231), .B2(n_255), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_262), .B(n_242), .Y(n_293) );
NAND4xp25_ASAP7_75t_SL g294 ( .A(n_266), .B(n_229), .C(n_85), .D(n_115), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_274), .A2(n_221), .B1(n_234), .B2(n_235), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_266), .B(n_113), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_264), .Y(n_297) );
OAI31xp33_ASAP7_75t_L g298 ( .A1(n_260), .A2(n_214), .A3(n_154), .B(n_113), .Y(n_298) );
AND2x4_ASAP7_75t_SL g299 ( .A(n_264), .B(n_227), .Y(n_299) );
NOR2x1_ASAP7_75t_L g300 ( .A(n_261), .B(n_242), .Y(n_300) );
INVx1_ASAP7_75t_SL g301 ( .A(n_264), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_261), .B(n_242), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_257), .B(n_242), .Y(n_303) );
INVxp67_ASAP7_75t_SL g304 ( .A(n_257), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_279), .B(n_267), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_297), .B(n_260), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_300), .B(n_302), .Y(n_307) );
AOI22xp5_ASAP7_75t_L g308 ( .A1(n_294), .A2(n_260), .B1(n_271), .B2(n_234), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_302), .B(n_260), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_285), .B(n_2), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_282), .Y(n_311) );
AND2x2_ASAP7_75t_SL g312 ( .A(n_283), .B(n_291), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_293), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_301), .B(n_267), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_286), .B(n_267), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_281), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_281), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_303), .Y(n_318) );
NAND3xp33_ASAP7_75t_L g319 ( .A(n_290), .B(n_121), .C(n_124), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_283), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_283), .B(n_268), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_304), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_299), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_291), .B(n_268), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_278), .B(n_268), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_299), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_277), .B(n_269), .Y(n_327) );
NOR2x1_ASAP7_75t_L g328 ( .A(n_288), .B(n_271), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_296), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_280), .B(n_2), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_292), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_290), .B(n_269), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_295), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_292), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_298), .B(n_269), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_289), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_287), .B(n_269), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_284), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_282), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_279), .B(n_269), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_279), .B(n_271), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_302), .B(n_273), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_281), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_282), .Y(n_344) );
INVxp67_ASAP7_75t_L g345 ( .A(n_279), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_302), .B(n_273), .Y(n_346) );
OAI21xp5_ASAP7_75t_L g347 ( .A1(n_310), .A2(n_106), .B(n_111), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_345), .B(n_3), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_338), .B(n_4), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_313), .B(n_273), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_305), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_312), .A2(n_233), .B1(n_227), .B2(n_275), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_339), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_311), .B(n_121), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_305), .B(n_105), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_339), .B(n_121), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_344), .B(n_121), .Y(n_357) );
AO22x1_ASAP7_75t_L g358 ( .A1(n_327), .A2(n_204), .B1(n_194), .B2(n_111), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_344), .Y(n_359) );
CKINVDCx14_ASAP7_75t_R g360 ( .A(n_323), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_322), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_340), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_340), .Y(n_363) );
NAND2x1_ASAP7_75t_SL g364 ( .A(n_327), .B(n_106), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_322), .Y(n_365) );
NAND4xp25_ASAP7_75t_L g366 ( .A(n_325), .B(n_114), .C(n_106), .D(n_8), .Y(n_366) );
INVx2_ASAP7_75t_SL g367 ( .A(n_321), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_321), .B(n_194), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_330), .A2(n_124), .B1(n_114), .B2(n_78), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_333), .A2(n_124), .B1(n_88), .B2(n_198), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_306), .B(n_124), .Y(n_371) );
INVx1_ASAP7_75t_SL g372 ( .A(n_321), .Y(n_372) );
NOR4xp25_ASAP7_75t_SL g373 ( .A(n_320), .B(n_6), .C(n_7), .D(n_9), .Y(n_373) );
NOR2x1_ASAP7_75t_L g374 ( .A(n_319), .B(n_198), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_329), .B(n_7), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_331), .A2(n_184), .B1(n_189), .B2(n_204), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_320), .Y(n_377) );
INVx1_ASAP7_75t_SL g378 ( .A(n_326), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_336), .A2(n_204), .B1(n_194), .B2(n_189), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_334), .B(n_10), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_336), .A2(n_204), .B1(n_194), .B2(n_189), .Y(n_381) );
NAND4xp25_ASAP7_75t_L g382 ( .A(n_341), .B(n_13), .C(n_14), .D(n_15), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_314), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_309), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_315), .Y(n_385) );
OAI211xp5_ASAP7_75t_L g386 ( .A1(n_332), .A2(n_189), .B(n_16), .C(n_17), .Y(n_386) );
INVxp67_ASAP7_75t_L g387 ( .A(n_332), .Y(n_387) );
AOI221xp5_ASAP7_75t_L g388 ( .A1(n_318), .A2(n_125), .B1(n_128), .B2(n_129), .C(n_132), .Y(n_388) );
INVx1_ASAP7_75t_SL g389 ( .A(n_326), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_318), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_342), .B(n_14), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_342), .B(n_16), .Y(n_392) );
OAI21xp5_ASAP7_75t_L g393 ( .A1(n_337), .A2(n_179), .B(n_144), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_383), .Y(n_394) );
NOR3xp33_ASAP7_75t_SL g395 ( .A(n_382), .B(n_316), .C(n_19), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_362), .B(n_346), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_363), .B(n_346), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_383), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_353), .Y(n_399) );
INVx1_ASAP7_75t_SL g400 ( .A(n_378), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_359), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_377), .Y(n_402) );
OAI211xp5_ASAP7_75t_L g403 ( .A1(n_360), .A2(n_324), .B(n_308), .C(n_335), .Y(n_403) );
NAND3xp33_ASAP7_75t_L g404 ( .A(n_349), .B(n_328), .C(n_337), .Y(n_404) );
NOR3xp33_ASAP7_75t_L g405 ( .A(n_349), .B(n_335), .C(n_324), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_385), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_368), .A2(n_389), .B1(n_372), .B2(n_367), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_392), .B(n_307), .Y(n_408) );
A2O1A1Ixp33_ASAP7_75t_L g409 ( .A1(n_366), .A2(n_307), .B(n_316), .C(n_343), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_365), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_387), .B(n_307), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_387), .B(n_343), .Y(n_412) );
XNOR2x1_ASAP7_75t_L g413 ( .A(n_358), .B(n_18), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_365), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_371), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_390), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_351), .Y(n_417) );
OAI21xp5_ASAP7_75t_L g418 ( .A1(n_386), .A2(n_317), .B(n_179), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_391), .B(n_317), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_384), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_355), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_361), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_368), .Y(n_423) );
NOR3xp33_ASAP7_75t_L g424 ( .A(n_348), .B(n_18), .C(n_19), .Y(n_424) );
NAND3xp33_ASAP7_75t_SL g425 ( .A(n_348), .B(n_178), .C(n_208), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_375), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_356), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_350), .B(n_144), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_380), .A2(n_147), .B1(n_137), .B2(n_189), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_380), .B(n_20), .Y(n_430) );
NAND3xp33_ASAP7_75t_L g431 ( .A(n_370), .B(n_147), .C(n_144), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_357), .B(n_147), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_374), .A2(n_205), .B(n_165), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g434 ( .A1(n_352), .A2(n_165), .B(n_138), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_394), .B(n_354), .Y(n_435) );
AOI21xp33_ASAP7_75t_L g436 ( .A1(n_413), .A2(n_347), .B(n_369), .Y(n_436) );
OAI211xp5_ASAP7_75t_L g437 ( .A1(n_403), .A2(n_364), .B(n_373), .C(n_393), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_398), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_406), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_416), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_422), .Y(n_441) );
XNOR2xp5_ASAP7_75t_L g442 ( .A(n_426), .B(n_376), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_405), .B(n_381), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_422), .Y(n_444) );
AOI21xp33_ASAP7_75t_SL g445 ( .A1(n_407), .A2(n_379), .B(n_24), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_396), .B(n_388), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_415), .B(n_147), .Y(n_447) );
NAND3xp33_ASAP7_75t_L g448 ( .A(n_395), .B(n_147), .C(n_159), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_399), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_410), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_400), .B(n_21), .Y(n_451) );
NAND3x2_ASAP7_75t_L g452 ( .A(n_421), .B(n_27), .C(n_31), .Y(n_452) );
XNOR2x1_ASAP7_75t_L g453 ( .A(n_408), .B(n_32), .Y(n_453) );
AOI32xp33_ASAP7_75t_L g454 ( .A1(n_424), .A2(n_156), .A3(n_162), .B1(n_158), .B2(n_35), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_397), .B(n_33), .Y(n_455) );
NOR2x1_ASAP7_75t_SL g456 ( .A(n_423), .B(n_39), .Y(n_456) );
INVxp67_ASAP7_75t_L g457 ( .A(n_414), .Y(n_457) );
INVx2_ASAP7_75t_SL g458 ( .A(n_417), .Y(n_458) );
OAI21xp33_ASAP7_75t_SL g459 ( .A1(n_411), .A2(n_40), .B(n_41), .Y(n_459) );
XNOR2x1_ASAP7_75t_L g460 ( .A(n_395), .B(n_419), .Y(n_460) );
NOR3xp33_ASAP7_75t_SL g461 ( .A(n_459), .B(n_409), .C(n_425), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_444), .B(n_412), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_446), .B(n_404), .Y(n_463) );
INVx3_ASAP7_75t_SL g464 ( .A(n_453), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g465 ( .A(n_448), .B(n_424), .C(n_425), .Y(n_465) );
INVx1_ASAP7_75t_SL g466 ( .A(n_453), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_460), .A2(n_443), .B1(n_446), .B2(n_442), .Y(n_467) );
XNOR2x1_ASAP7_75t_L g468 ( .A(n_460), .B(n_420), .Y(n_468) );
CKINVDCx16_ASAP7_75t_R g469 ( .A(n_455), .Y(n_469) );
INVx4_ASAP7_75t_L g470 ( .A(n_444), .Y(n_470) );
NAND2x1p5_ASAP7_75t_L g471 ( .A(n_451), .B(n_430), .Y(n_471) );
AOI322xp5_ASAP7_75t_L g472 ( .A1(n_458), .A2(n_402), .A3(n_401), .B1(n_429), .B2(n_427), .C1(n_428), .C2(n_418), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_439), .B(n_429), .Y(n_473) );
OAI221xp5_ASAP7_75t_SL g474 ( .A1(n_454), .A2(n_434), .B1(n_432), .B2(n_433), .C(n_431), .Y(n_474) );
INVxp67_ASAP7_75t_SL g475 ( .A(n_441), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_457), .B(n_42), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_445), .A2(n_156), .B(n_47), .C(n_49), .Y(n_477) );
OAI221xp5_ASAP7_75t_L g478 ( .A1(n_437), .A2(n_156), .B1(n_50), .B2(n_53), .C(n_55), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_436), .A2(n_174), .B1(n_173), .B2(n_167), .Y(n_479) );
AOI32xp33_ASAP7_75t_L g480 ( .A1(n_458), .A2(n_45), .A3(n_56), .B1(n_57), .B2(n_58), .Y(n_480) );
OAI22xp33_ASAP7_75t_L g481 ( .A1(n_441), .A2(n_435), .B1(n_440), .B2(n_438), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_449), .B(n_59), .Y(n_482) );
AOI211xp5_ASAP7_75t_L g483 ( .A1(n_455), .A2(n_63), .B(n_148), .C(n_155), .Y(n_483) );
OA22x2_ASAP7_75t_L g484 ( .A1(n_450), .A2(n_148), .B1(n_155), .B2(n_167), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_450), .B(n_155), .Y(n_485) );
BUFx12f_ASAP7_75t_L g486 ( .A(n_470), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_467), .A2(n_464), .B1(n_469), .B2(n_463), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_470), .B(n_462), .Y(n_488) );
OAI21x1_ASAP7_75t_SL g489 ( .A1(n_468), .A2(n_477), .B(n_456), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_473), .Y(n_490) );
AOI31xp33_ASAP7_75t_L g491 ( .A1(n_487), .A2(n_466), .A3(n_478), .B(n_471), .Y(n_491) );
XNOR2xp5_ASAP7_75t_L g492 ( .A(n_490), .B(n_461), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_486), .A2(n_465), .B1(n_481), .B2(n_475), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_492), .Y(n_494) );
OAI221xp5_ASAP7_75t_L g495 ( .A1(n_491), .A2(n_488), .B1(n_472), .B2(n_489), .C(n_474), .Y(n_495) );
OAI322xp33_ASAP7_75t_L g496 ( .A1(n_494), .A2(n_493), .A3(n_476), .B1(n_482), .B2(n_447), .C1(n_484), .C2(n_485), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_496), .A2(n_495), .B1(n_452), .B2(n_479), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_497), .A2(n_480), .B(n_483), .Y(n_498) );
endmodule