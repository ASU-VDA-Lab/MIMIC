module fake_jpeg_7819_n_75 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_75);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_75;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_73;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_72;
wire n_49;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_74;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_32;
wire n_70;
wire n_66;

BUFx5_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_9),
.B(n_11),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_37),
.Y(n_47)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_28),
.B(n_26),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_48),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_51),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_16),
.B1(n_21),
.B2(n_2),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_57)
);

NOR2x1_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_50),
.Y(n_59)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_8),
.B(n_10),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_1),
.C(n_3),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_12),
.C(n_14),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_62),
.Y(n_67)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_48),
.B1(n_59),
.B2(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_67),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_60),
.C(n_63),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_47),
.C(n_58),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_55),
.B1(n_42),
.B2(n_58),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_45),
.B(n_65),
.Y(n_74)
);

XNOR2x2_ASAP7_75t_SL g75 ( 
.A(n_74),
.B(n_64),
.Y(n_75)
);


endmodule