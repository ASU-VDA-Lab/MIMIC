module fake_netlist_6_1796_n_1824 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1824);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1824;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_39),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_130),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_24),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_129),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_53),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_176),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_120),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_79),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_65),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_121),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_106),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_74),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_98),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_168),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_5),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_37),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_26),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_163),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_118),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_67),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_97),
.Y(n_200)
);

BUFx8_ASAP7_75t_SL g201 ( 
.A(n_162),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_43),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_111),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_34),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_109),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_107),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_8),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_75),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_11),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_11),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_17),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_58),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_45),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_166),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_25),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_0),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g217 ( 
.A(n_34),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_178),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_54),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_175),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_24),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_154),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_28),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_156),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_31),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_167),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_160),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_28),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_159),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_23),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_93),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_155),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_32),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_71),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_45),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_73),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_19),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_134),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_150),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_19),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_147),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_102),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_91),
.Y(n_243)
);

BUFx2_ASAP7_75t_SL g244 ( 
.A(n_44),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_85),
.Y(n_245)
);

INVxp33_ASAP7_75t_SL g246 ( 
.A(n_100),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_94),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_47),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_31),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_143),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_137),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_123),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_20),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_1),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_144),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_177),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_59),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_52),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_149),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_39),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_128),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_113),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_1),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_40),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_81),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_133),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_33),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_32),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_96),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_136),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_82),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_114),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_66),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_104),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_53),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_18),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_43),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_47),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_42),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_27),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_145),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_157),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_63),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_16),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_14),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_10),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_103),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_48),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_23),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_88),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_135),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_92),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_117),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_72),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_112),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_161),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_6),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_87),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_36),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_174),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_108),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_2),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_83),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_17),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_84),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_70),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_99),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_115),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_18),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_55),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_125),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_148),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_3),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_35),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_15),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_86),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_132),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_9),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_64),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_76),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_35),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_37),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_126),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_78),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_25),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_2),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_46),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_60),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_89),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_4),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_49),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_171),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_38),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_122),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_142),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_46),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_30),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_105),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_62),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_152),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_36),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_51),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_164),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_54),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_110),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_173),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_29),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_21),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_14),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_56),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_140),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_49),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_12),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_6),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_15),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_131),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_226),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_189),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_191),
.B(n_0),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_179),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_210),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_205),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_191),
.B(n_3),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_243),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_189),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_195),
.B(n_263),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_181),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_193),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_193),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_212),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_212),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_227),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_251),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_197),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_262),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_211),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_246),
.B(n_4),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_227),
.B(n_231),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_290),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_183),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_214),
.B(n_5),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_211),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_226),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_194),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_316),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_202),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_219),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_231),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_343),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_308),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_196),
.B(n_7),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_232),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_201),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_232),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_238),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_221),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_238),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_242),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_242),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_308),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_223),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_210),
.B(n_7),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_278),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_230),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_245),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_197),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_245),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_295),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_214),
.B(n_8),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_259),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_295),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_211),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_235),
.Y(n_413)
);

INVxp33_ASAP7_75t_SL g414 ( 
.A(n_330),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_338),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_259),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_265),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_217),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_180),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_240),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_265),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_211),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_229),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_249),
.Y(n_424)
);

INVxp33_ASAP7_75t_SL g425 ( 
.A(n_278),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_182),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_217),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_338),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_273),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_258),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_273),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_281),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_211),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_264),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_267),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_336),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_336),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_268),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_276),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_279),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_280),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_284),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_281),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_285),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_287),
.B(n_9),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_287),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_422),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_393),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_423),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_376),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_423),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_L g452 ( 
.A(n_376),
.B(n_257),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_419),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_382),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_383),
.B(n_350),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_423),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_360),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_426),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_357),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_357),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_390),
.B(n_257),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_366),
.B(n_275),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_382),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_412),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_422),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_412),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_423),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_360),
.Y(n_468)
);

CKINVDCx11_ASAP7_75t_R g469 ( 
.A(n_406),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_433),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_367),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_367),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_380),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_400),
.B(n_296),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_423),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_362),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_433),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_436),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_415),
.B(n_296),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_364),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_380),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_436),
.Y(n_482)
);

OR2x6_ASAP7_75t_L g483 ( 
.A(n_363),
.B(n_350),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_384),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_384),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_437),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_437),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_358),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_365),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_368),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_369),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_370),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_386),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_371),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_372),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_373),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_388),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_386),
.Y(n_498)
);

BUFx8_ASAP7_75t_L g499 ( 
.A(n_402),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_392),
.Y(n_500)
);

BUFx8_ASAP7_75t_L g501 ( 
.A(n_402),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_394),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_375),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_395),
.Y(n_504)
);

AND2x6_ASAP7_75t_L g505 ( 
.A(n_378),
.B(n_229),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_397),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_398),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_R g508 ( 
.A(n_387),
.B(n_184),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_387),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_446),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_428),
.B(n_353),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_399),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_405),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_396),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_407),
.B(n_320),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_396),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_401),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_401),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_410),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_416),
.B(n_320),
.Y(n_520)
);

AND3x2_ASAP7_75t_L g521 ( 
.A(n_359),
.B(n_353),
.C(n_216),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_404),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_417),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_421),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_482),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_505),
.B(n_429),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_451),
.Y(n_527)
);

NAND2xp33_ASAP7_75t_SL g528 ( 
.A(n_455),
.B(n_233),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_455),
.B(n_374),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_511),
.B(n_404),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_510),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_461),
.B(n_414),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_510),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_505),
.A2(n_445),
.B1(n_391),
.B2(n_381),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_459),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_474),
.B(n_425),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_459),
.B(n_460),
.Y(n_537)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_483),
.B(n_244),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_510),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_L g540 ( 
.A(n_505),
.B(n_229),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_459),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_476),
.B(n_379),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_451),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_482),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_482),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_505),
.A2(n_391),
.B1(n_409),
.B2(n_260),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_499),
.B(n_377),
.Y(n_547)
);

OR2x6_ASAP7_75t_L g548 ( 
.A(n_483),
.B(n_244),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_451),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_511),
.B(n_413),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_505),
.B(n_431),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_479),
.B(n_413),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_510),
.Y(n_553)
);

CKINVDCx6p67_ASAP7_75t_R g554 ( 
.A(n_469),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_460),
.B(n_420),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_451),
.Y(n_556)
);

OR2x6_ASAP7_75t_L g557 ( 
.A(n_483),
.B(n_361),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_488),
.Y(n_558)
);

AND2x6_ASAP7_75t_L g559 ( 
.A(n_520),
.B(n_291),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_505),
.B(n_460),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_487),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_505),
.A2(n_260),
.B1(n_209),
.B2(n_322),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_488),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_L g564 ( 
.A(n_505),
.B(n_229),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_508),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_491),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_478),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_478),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_500),
.B(n_420),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_483),
.A2(n_302),
.B1(n_216),
.B2(n_209),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_491),
.Y(n_571)
);

NOR3xp33_ASAP7_75t_L g572 ( 
.A(n_473),
.B(n_427),
.C(n_418),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_500),
.B(n_424),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_473),
.B(n_424),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_480),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_492),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_483),
.A2(n_302),
.B1(n_297),
.B2(n_322),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_457),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_500),
.B(n_430),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_451),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_492),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_472),
.B(n_430),
.Y(n_582)
);

NAND2x1p5_ASAP7_75t_L g583 ( 
.A(n_520),
.B(n_269),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_472),
.B(n_434),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_495),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_485),
.B(n_403),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_499),
.B(n_324),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_499),
.B(n_324),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_L g589 ( 
.A(n_493),
.B(n_435),
.C(n_434),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_447),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_490),
.B(n_432),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_522),
.B(n_435),
.Y(n_592)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_496),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_490),
.B(n_438),
.Y(n_594)
);

AND2x6_ASAP7_75t_L g595 ( 
.A(n_520),
.B(n_291),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_490),
.B(n_443),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_510),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_520),
.A2(n_297),
.B1(n_321),
.B2(n_349),
.Y(n_598)
);

NOR3xp33_ASAP7_75t_L g599 ( 
.A(n_468),
.B(n_439),
.C(n_438),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_521),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_490),
.B(n_439),
.Y(n_601)
);

CKINVDCx6p67_ASAP7_75t_R g602 ( 
.A(n_503),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_447),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_SL g604 ( 
.A(n_471),
.B(n_233),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_510),
.B(n_440),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_495),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_453),
.Y(n_607)
);

BUFx10_ASAP7_75t_L g608 ( 
.A(n_481),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_447),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_465),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_497),
.B(n_440),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_465),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_497),
.Y(n_613)
);

INVx5_ASAP7_75t_L g614 ( 
.A(n_451),
.Y(n_614)
);

INVx5_ASAP7_75t_L g615 ( 
.A(n_456),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_513),
.B(n_441),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_458),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_502),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_502),
.B(n_441),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_456),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_504),
.Y(n_621)
);

INVx5_ASAP7_75t_L g622 ( 
.A(n_456),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_513),
.B(n_442),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_456),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_456),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_484),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_465),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_456),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_498),
.B(n_442),
.Y(n_629)
);

INVx4_ASAP7_75t_SL g630 ( 
.A(n_475),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_509),
.A2(n_444),
.B1(n_411),
.B2(n_408),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_504),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_513),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_513),
.B(n_444),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_462),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_486),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_486),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_507),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_507),
.Y(n_639)
);

INVx5_ASAP7_75t_L g640 ( 
.A(n_475),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_512),
.B(n_321),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_512),
.B(n_366),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_513),
.B(n_282),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g644 ( 
.A(n_514),
.B(n_385),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_499),
.B(n_229),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_SL g646 ( 
.A(n_516),
.B(n_389),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_513),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_517),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_519),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_519),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_489),
.B(n_292),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_486),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_524),
.Y(n_653)
);

NOR2x1p5_ASAP7_75t_L g654 ( 
.A(n_518),
.B(n_288),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_519),
.B(n_349),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_462),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_501),
.B(n_292),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_475),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_519),
.B(n_356),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_489),
.B(n_300),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_487),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_450),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_519),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_519),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_450),
.Y(n_665)
);

OR2x6_ASAP7_75t_L g666 ( 
.A(n_494),
.B(n_196),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_501),
.B(n_300),
.Y(n_667)
);

AND2x6_ASAP7_75t_L g668 ( 
.A(n_494),
.B(n_303),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_501),
.B(n_523),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_506),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_501),
.B(n_303),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_448),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_523),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_523),
.B(n_185),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_454),
.Y(n_675)
);

AND2x6_ASAP7_75t_L g676 ( 
.A(n_506),
.B(n_312),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_523),
.B(n_187),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_662),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_537),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_552),
.B(n_523),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_552),
.B(n_523),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_555),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_574),
.B(n_188),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_672),
.Y(n_684)
);

BUFx6f_ASAP7_75t_SL g685 ( 
.A(n_608),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_530),
.B(n_190),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_594),
.A2(n_252),
.B1(n_198),
.B2(n_351),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_670),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_586),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_537),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_594),
.B(n_524),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_586),
.Y(n_692)
);

OR2x6_ASAP7_75t_L g693 ( 
.A(n_538),
.B(n_204),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_529),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_550),
.B(n_192),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_536),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_536),
.B(n_524),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_532),
.A2(n_271),
.B1(n_307),
.B2(n_270),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_532),
.B(n_524),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_673),
.A2(n_515),
.B(n_475),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_537),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_665),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_665),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_L g704 ( 
.A1(n_538),
.A2(n_312),
.B1(n_340),
.B2(n_346),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_546),
.B(n_524),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_546),
.B(n_524),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_558),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_611),
.B(n_289),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_611),
.B(n_299),
.Y(n_709)
);

BUFx6f_ASAP7_75t_SL g710 ( 
.A(n_608),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_563),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_619),
.B(n_309),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_565),
.B(n_199),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_569),
.B(n_200),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_619),
.B(n_310),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_675),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_675),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_601),
.B(n_313),
.Y(n_718)
);

OR2x6_ASAP7_75t_L g719 ( 
.A(n_538),
.B(n_204),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_567),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_582),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_525),
.B(n_454),
.Y(n_722)
);

AND2x6_ASAP7_75t_SL g723 ( 
.A(n_586),
.B(n_207),
.Y(n_723)
);

INVx4_ASAP7_75t_L g724 ( 
.A(n_535),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_544),
.B(n_463),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_566),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_569),
.B(n_206),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_590),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_534),
.A2(n_331),
.B1(n_207),
.B2(n_213),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_571),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_545),
.B(n_463),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_576),
.Y(n_732)
);

AND2x4_ASAP7_75t_SL g733 ( 
.A(n_602),
.B(n_186),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_659),
.B(n_464),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_573),
.B(n_208),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_573),
.B(n_579),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_579),
.B(n_314),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_R g738 ( 
.A(n_672),
.B(n_218),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_528),
.A2(n_247),
.B1(n_220),
.B2(n_345),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_673),
.A2(n_475),
.B(n_467),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_567),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_659),
.B(n_464),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_656),
.B(n_315),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_528),
.A2(n_239),
.B1(n_222),
.B2(n_224),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_534),
.B(n_466),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_L g746 ( 
.A(n_559),
.B(n_234),
.Y(n_746)
);

INVx8_ASAP7_75t_L g747 ( 
.A(n_548),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_581),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_570),
.B(n_236),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_570),
.B(n_241),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_605),
.B(n_466),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_585),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_616),
.B(n_470),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_623),
.B(n_318),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_535),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_634),
.B(n_470),
.Y(n_756)
);

NOR3xp33_ASAP7_75t_L g757 ( 
.A(n_631),
.B(n_333),
.C(n_325),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_584),
.Y(n_758)
);

OR2x6_ASAP7_75t_L g759 ( 
.A(n_548),
.B(n_213),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_606),
.A2(n_613),
.B(n_621),
.C(n_618),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_632),
.B(n_638),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_568),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_639),
.B(n_643),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_655),
.B(n_477),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_577),
.B(n_250),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_589),
.B(n_326),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_557),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_541),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_655),
.B(n_477),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_629),
.B(n_506),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_541),
.B(n_327),
.Y(n_771)
);

OAI21xp5_ASAP7_75t_L g772 ( 
.A1(n_560),
.A2(n_551),
.B(n_526),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_651),
.B(n_340),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_583),
.B(n_337),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_583),
.B(n_449),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_590),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_591),
.B(n_449),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_577),
.B(n_578),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_603),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_592),
.B(n_255),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_596),
.B(n_449),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_674),
.B(n_449),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_651),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_599),
.B(n_256),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_626),
.B(n_217),
.Y(n_785)
);

NAND2x1_ASAP7_75t_L g786 ( 
.A(n_527),
.B(n_475),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_648),
.B(n_217),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_677),
.B(n_487),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_604),
.B(n_261),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_604),
.B(n_266),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_587),
.B(n_272),
.Y(n_791)
);

A2O1A1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_641),
.A2(n_346),
.B(n_452),
.C(n_237),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_603),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_609),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_669),
.A2(n_317),
.B1(n_274),
.B2(n_323),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_609),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_587),
.B(n_283),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_548),
.B(n_341),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_588),
.B(n_293),
.Y(n_799)
);

NOR3xp33_ASAP7_75t_L g800 ( 
.A(n_642),
.B(n_347),
.C(n_354),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_597),
.B(n_487),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_557),
.B(n_575),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_610),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_562),
.A2(n_311),
.B1(n_294),
.B2(n_298),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_660),
.Y(n_805)
);

NOR3xp33_ASAP7_75t_L g806 ( 
.A(n_547),
.B(n_352),
.C(n_342),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_597),
.B(n_487),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_660),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_633),
.B(n_487),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_588),
.B(n_657),
.Y(n_810)
);

NOR2xp67_ASAP7_75t_L g811 ( 
.A(n_669),
.B(n_301),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_657),
.B(n_305),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_610),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_660),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_612),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_666),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_666),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_633),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_600),
.B(n_344),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_667),
.B(n_671),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_667),
.B(n_306),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_647),
.B(n_467),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_671),
.B(n_319),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_647),
.B(n_467),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_612),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_627),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_645),
.B(n_328),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_557),
.B(n_329),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_645),
.B(n_332),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_598),
.B(n_572),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_627),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_598),
.B(n_334),
.Y(n_832)
);

NAND2xp33_ASAP7_75t_SL g833 ( 
.A(n_654),
.B(n_277),
.Y(n_833)
);

AO221x1_ASAP7_75t_L g834 ( 
.A1(n_527),
.A2(n_336),
.B1(n_355),
.B2(n_215),
.C(n_225),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_562),
.A2(n_254),
.B1(n_355),
.B2(n_348),
.Y(n_835)
);

O2A1O1Ixp5_ASAP7_75t_L g836 ( 
.A1(n_641),
.A2(n_254),
.B(n_348),
.C(n_215),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_666),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_636),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_636),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_SL g840 ( 
.A(n_547),
.B(n_339),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_608),
.B(n_335),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_649),
.B(n_653),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_637),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_637),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_663),
.B(n_452),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_652),
.Y(n_846)
);

NOR2xp67_ASAP7_75t_L g847 ( 
.A(n_721),
.B(n_652),
.Y(n_847)
);

O2A1O1Ixp5_ASAP7_75t_L g848 ( 
.A1(n_820),
.A2(n_553),
.B(n_531),
.C(n_664),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_768),
.B(n_593),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_691),
.A2(n_540),
.B(n_564),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_788),
.A2(n_540),
.B(n_564),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_696),
.B(n_644),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_679),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_680),
.A2(n_539),
.B(n_531),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_678),
.Y(n_855)
);

NAND2x1p5_ASAP7_75t_L g856 ( 
.A(n_679),
.B(n_533),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_681),
.A2(n_650),
.B(n_533),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_758),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_678),
.Y(n_859)
);

OAI21xp33_ASAP7_75t_L g860 ( 
.A1(n_708),
.A2(n_646),
.B(n_228),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_699),
.B(n_559),
.Y(n_861)
);

O2A1O1Ixp5_ASAP7_75t_L g862 ( 
.A1(n_820),
.A2(n_553),
.B(n_539),
.C(n_664),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_679),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_720),
.Y(n_864)
);

NOR3xp33_ASAP7_75t_L g865 ( 
.A(n_708),
.B(n_607),
.C(n_617),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_763),
.A2(n_650),
.B(n_561),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_720),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_782),
.A2(n_561),
.B(n_661),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_768),
.B(n_701),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_736),
.B(n_542),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_705),
.A2(n_595),
.B(n_559),
.Y(n_871)
);

INVx5_ASAP7_75t_L g872 ( 
.A(n_679),
.Y(n_872)
);

AOI21x1_ASAP7_75t_L g873 ( 
.A1(n_740),
.A2(n_630),
.B(n_561),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_706),
.A2(n_661),
.B(n_620),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_772),
.A2(n_661),
.B(n_620),
.Y(n_875)
);

AOI21x1_ASAP7_75t_L g876 ( 
.A1(n_700),
.A2(n_630),
.B(n_543),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_709),
.A2(n_595),
.B1(n_668),
.B2(n_676),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_709),
.A2(n_595),
.B1(n_668),
.B2(n_676),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_751),
.A2(n_756),
.B(n_753),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_770),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_741),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_697),
.B(n_595),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_818),
.A2(n_580),
.B(n_620),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_754),
.B(n_595),
.Y(n_884)
);

NAND2x1_ASAP7_75t_L g885 ( 
.A(n_818),
.B(n_543),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_702),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_801),
.A2(n_625),
.B(n_620),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_702),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_703),
.Y(n_889)
);

AOI21x1_ASAP7_75t_L g890 ( 
.A1(n_786),
.A2(n_630),
.B(n_549),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_712),
.A2(n_715),
.B(n_737),
.C(n_821),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_729),
.B(n_549),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_754),
.B(n_556),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_694),
.B(n_580),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_712),
.B(n_556),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_807),
.A2(n_628),
.B(n_580),
.Y(n_896)
);

INVx11_ASAP7_75t_L g897 ( 
.A(n_685),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_715),
.B(n_635),
.Y(n_898)
);

NAND2x1p5_ASAP7_75t_L g899 ( 
.A(n_690),
.B(n_624),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_809),
.A2(n_628),
.B(n_625),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_718),
.B(n_624),
.Y(n_901)
);

AND2x6_ASAP7_75t_L g902 ( 
.A(n_745),
.B(n_225),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_729),
.A2(n_658),
.B(n_676),
.Y(n_903)
);

BUFx12f_ASAP7_75t_L g904 ( 
.A(n_723),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_718),
.B(n_625),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_755),
.B(n_625),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_822),
.A2(n_628),
.B(n_658),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_783),
.B(n_668),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_835),
.A2(n_228),
.B1(n_237),
.B2(n_248),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_835),
.A2(n_248),
.B1(n_253),
.B2(n_304),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_701),
.B(n_668),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_783),
.B(n_668),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_716),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_824),
.A2(n_628),
.B(n_640),
.Y(n_914)
);

INVx4_ASAP7_75t_L g915 ( 
.A(n_755),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_707),
.B(n_676),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_743),
.B(n_635),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_716),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_711),
.B(n_676),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_778),
.A2(n_186),
.B(n_203),
.C(n_286),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_734),
.B(n_622),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_726),
.B(n_730),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_732),
.B(n_622),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_777),
.A2(n_781),
.B(n_775),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_810),
.A2(n_186),
.B1(n_203),
.B2(n_554),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_742),
.B(n_640),
.Y(n_926)
);

NOR2xp67_ASAP7_75t_L g927 ( 
.A(n_821),
.B(n_77),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_690),
.A2(n_761),
.B(n_764),
.Y(n_928)
);

BUFx4f_ASAP7_75t_L g929 ( 
.A(n_747),
.Y(n_929)
);

BUFx8_ASAP7_75t_L g930 ( 
.A(n_685),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_717),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_748),
.B(n_622),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_752),
.B(n_622),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_769),
.A2(n_640),
.B(n_615),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_845),
.A2(n_640),
.B(n_615),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_830),
.B(n_286),
.Y(n_936)
);

CKINVDCx10_ASAP7_75t_R g937 ( 
.A(n_710),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_755),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_689),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_762),
.Y(n_940)
);

AOI21x1_ASAP7_75t_L g941 ( 
.A1(n_722),
.A2(n_731),
.B(n_725),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_805),
.B(n_614),
.Y(n_942)
);

INVx1_ASAP7_75t_SL g943 ( 
.A(n_684),
.Y(n_943)
);

AOI21x1_ASAP7_75t_L g944 ( 
.A1(n_838),
.A2(n_615),
.B(n_614),
.Y(n_944)
);

INVxp67_ASAP7_75t_L g945 ( 
.A(n_785),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_766),
.B(n_286),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_823),
.A2(n_203),
.B1(n_186),
.B2(n_336),
.Y(n_947)
);

INVxp67_ASAP7_75t_L g948 ( 
.A(n_771),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_808),
.B(n_615),
.Y(n_949)
);

AO21x1_ASAP7_75t_L g950 ( 
.A1(n_823),
.A2(n_203),
.B(n_12),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_814),
.B(n_614),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_766),
.A2(n_336),
.B(n_286),
.C(n_16),
.Y(n_952)
);

NAND3xp33_ASAP7_75t_L g953 ( 
.A(n_819),
.B(n_10),
.C(n_13),
.Y(n_953)
);

NOR2x1p5_ASAP7_75t_SL g954 ( 
.A(n_846),
.B(n_61),
.Y(n_954)
);

AO21x1_ASAP7_75t_L g955 ( 
.A1(n_840),
.A2(n_13),
.B(n_20),
.Y(n_955)
);

AOI21x1_ASAP7_75t_L g956 ( 
.A1(n_839),
.A2(n_68),
.B(n_170),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_842),
.A2(n_760),
.B(n_746),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_755),
.B(n_172),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_774),
.A2(n_22),
.B(n_26),
.C(n_27),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_806),
.A2(n_834),
.B1(n_773),
.B2(n_765),
.Y(n_960)
);

AOI21xp33_ASAP7_75t_L g961 ( 
.A1(n_749),
.A2(n_22),
.B(n_29),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_774),
.A2(n_80),
.B1(n_165),
.B2(n_153),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_773),
.B(n_688),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_771),
.B(n_30),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_819),
.A2(n_33),
.B(n_38),
.C(n_40),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_714),
.B(n_41),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_776),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_842),
.A2(n_95),
.B(n_151),
.Y(n_968)
);

INVx4_ASAP7_75t_L g969 ( 
.A(n_724),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_836),
.A2(n_90),
.B(n_146),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_846),
.A2(n_69),
.B(n_141),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_827),
.A2(n_169),
.B(n_139),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_724),
.B(n_138),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_776),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_811),
.A2(n_41),
.B(n_42),
.C(n_44),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_727),
.B(n_48),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_735),
.B(n_50),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_779),
.Y(n_978)
);

INVx11_ASAP7_75t_L g979 ( 
.A(n_710),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_802),
.B(n_50),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_SL g981 ( 
.A(n_747),
.B(n_51),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_798),
.A2(n_812),
.B(n_816),
.C(n_837),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_829),
.A2(n_101),
.B(n_124),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_SL g984 ( 
.A(n_747),
.B(n_52),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_787),
.B(n_55),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_843),
.A2(n_116),
.B(n_119),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_844),
.A2(n_127),
.B(n_57),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_698),
.B(n_57),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_793),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_728),
.A2(n_815),
.B(n_831),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_687),
.B(n_739),
.Y(n_991)
);

AND2x6_ASAP7_75t_L g992 ( 
.A(n_817),
.B(n_825),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_793),
.B(n_803),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_794),
.A2(n_813),
.B(n_803),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_796),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_692),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_738),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_683),
.B(n_686),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_798),
.A2(n_750),
.B(n_797),
.C(n_799),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_695),
.B(n_733),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_733),
.B(n_757),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_704),
.A2(n_693),
.B1(n_719),
.B2(n_759),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_828),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_796),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_813),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_825),
.A2(n_831),
.B(n_826),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_826),
.A2(n_791),
.B(n_713),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_780),
.A2(n_790),
.B(n_789),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_792),
.A2(n_832),
.B(n_804),
.C(n_784),
.Y(n_1009)
);

INVxp67_ASAP7_75t_L g1010 ( 
.A(n_828),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_841),
.A2(n_693),
.B(n_719),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_693),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_719),
.A2(n_759),
.B(n_795),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_759),
.A2(n_767),
.B(n_800),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_744),
.B(n_833),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_738),
.A2(n_673),
.B(n_691),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_699),
.B(n_697),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_696),
.B(n_736),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_SL g1019 ( 
.A1(n_810),
.A2(n_745),
.B(n_706),
.C(n_705),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_696),
.B(n_682),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_696),
.B(n_736),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_696),
.B(n_682),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_679),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_691),
.A2(n_673),
.B(n_788),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_678),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_1017),
.A2(n_891),
.B(n_1024),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_967),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_849),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_SL g1029 ( 
.A1(n_971),
.A2(n_1008),
.B(n_955),
.Y(n_1029)
);

AOI21xp33_ASAP7_75t_L g1030 ( 
.A1(n_946),
.A2(n_898),
.B(n_936),
.Y(n_1030)
);

AOI21x1_ASAP7_75t_L g1031 ( 
.A1(n_905),
.A2(n_893),
.B(n_875),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_994),
.A2(n_1006),
.B(n_896),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_880),
.B(n_1018),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_887),
.A2(n_900),
.B(n_944),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_880),
.B(n_1021),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_853),
.Y(n_1036)
);

AOI21xp33_ASAP7_75t_L g1037 ( 
.A1(n_991),
.A2(n_860),
.B(n_988),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_890),
.A2(n_868),
.B(n_907),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_882),
.A2(n_861),
.B(n_1019),
.Y(n_1039)
);

AOI21x1_ASAP7_75t_L g1040 ( 
.A1(n_901),
.A2(n_895),
.B(n_861),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_974),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_849),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_978),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_957),
.A2(n_928),
.B(n_884),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_855),
.Y(n_1045)
);

AOI21x1_ASAP7_75t_SL g1046 ( 
.A1(n_964),
.A2(n_976),
.B(n_966),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_854),
.A2(n_857),
.B(n_924),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_892),
.A2(n_850),
.B(n_903),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_859),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_869),
.B(n_1012),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_892),
.A2(n_903),
.B(n_871),
.Y(n_1051)
);

AOI21x1_ASAP7_75t_SL g1052 ( 
.A1(n_977),
.A2(n_912),
.B(n_908),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_851),
.A2(n_871),
.B(n_921),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_914),
.A2(n_990),
.B(n_883),
.Y(n_1054)
);

AOI22x1_ASAP7_75t_L g1055 ( 
.A1(n_1007),
.A2(n_1016),
.B1(n_866),
.B2(n_995),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_864),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_993),
.A2(n_848),
.B(n_862),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_921),
.A2(n_926),
.B(n_927),
.Y(n_1058)
);

AND2x6_ASAP7_75t_L g1059 ( 
.A(n_911),
.B(n_853),
.Y(n_1059)
);

AO21x1_ASAP7_75t_L g1060 ( 
.A1(n_1009),
.A2(n_970),
.B(n_971),
.Y(n_1060)
);

AO21x2_ASAP7_75t_L g1061 ( 
.A1(n_926),
.A2(n_878),
.B(n_877),
.Y(n_1061)
);

NOR2x1_ASAP7_75t_L g1062 ( 
.A(n_969),
.B(n_915),
.Y(n_1062)
);

O2A1O1Ixp5_ASAP7_75t_L g1063 ( 
.A1(n_970),
.A2(n_950),
.B(n_941),
.C(n_999),
.Y(n_1063)
);

OA22x2_ASAP7_75t_L g1064 ( 
.A1(n_925),
.A2(n_852),
.B1(n_945),
.B2(n_1003),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_948),
.B(n_922),
.Y(n_1065)
);

BUFx4f_ASAP7_75t_L g1066 ( 
.A(n_1015),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_867),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_847),
.B(n_902),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_993),
.A2(n_935),
.B(n_885),
.Y(n_1069)
);

AOI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_1010),
.A2(n_870),
.B1(n_998),
.B2(n_865),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_916),
.A2(n_919),
.B(n_872),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_872),
.A2(n_982),
.B(n_951),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_872),
.A2(n_949),
.B(n_942),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_886),
.A2(n_1025),
.B(n_931),
.Y(n_1074)
);

AO22x1_ASAP7_75t_L g1075 ( 
.A1(n_917),
.A2(n_997),
.B1(n_1015),
.B2(n_943),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_961),
.A2(n_902),
.B1(n_953),
.B2(n_909),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_888),
.A2(n_918),
.B(n_913),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_902),
.B(n_985),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_872),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_961),
.A2(n_959),
.B(n_965),
.C(n_952),
.Y(n_1080)
);

INVx2_ASAP7_75t_SL g1081 ( 
.A(n_996),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_902),
.B(n_963),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_1001),
.A2(n_869),
.B1(n_1000),
.B2(n_1002),
.Y(n_1083)
);

NOR2xp67_ASAP7_75t_SL g1084 ( 
.A(n_863),
.B(n_969),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_863),
.B(n_960),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_856),
.A2(n_899),
.B(n_934),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_889),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_938),
.B(n_1023),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_939),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_906),
.A2(n_1013),
.B(n_973),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_938),
.B(n_1023),
.Y(n_1091)
);

OAI22x1_ASAP7_75t_L g1092 ( 
.A1(n_947),
.A2(n_943),
.B1(n_858),
.B2(n_980),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_881),
.B(n_940),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_911),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_923),
.A2(n_933),
.B(n_932),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_930),
.Y(n_1096)
);

OAI22x1_ASAP7_75t_L g1097 ( 
.A1(n_1020),
.A2(n_1022),
.B1(n_984),
.B2(n_981),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1011),
.A2(n_968),
.B(n_894),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_989),
.A2(n_1005),
.B(n_1004),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_992),
.B(n_1014),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_SL g1101 ( 
.A1(n_972),
.A2(n_983),
.B(n_956),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_986),
.A2(n_958),
.B(n_987),
.Y(n_1102)
);

OAI21xp33_ASAP7_75t_L g1103 ( 
.A1(n_981),
.A2(n_984),
.B(n_909),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_962),
.A2(n_920),
.B(n_1002),
.Y(n_1104)
);

AOI21x1_ASAP7_75t_L g1105 ( 
.A1(n_910),
.A2(n_954),
.B(n_992),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_992),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_975),
.A2(n_929),
.B(n_910),
.Y(n_1107)
);

AOI21x1_ASAP7_75t_L g1108 ( 
.A1(n_992),
.A2(n_929),
.B(n_897),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_979),
.A2(n_930),
.B(n_937),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_904),
.B(n_1017),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1017),
.A2(n_891),
.B(n_1024),
.Y(n_1111)
);

OA21x2_ASAP7_75t_L g1112 ( 
.A1(n_1017),
.A2(n_1024),
.B(n_957),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_880),
.B(n_696),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_855),
.Y(n_1114)
);

OA22x2_ASAP7_75t_L g1115 ( 
.A1(n_925),
.A2(n_696),
.B1(n_483),
.B2(n_721),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_891),
.A2(n_1017),
.B(n_879),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1017),
.B(n_696),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1017),
.A2(n_891),
.B(n_1024),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1017),
.A2(n_891),
.B(n_1024),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_988),
.A2(n_729),
.B1(n_820),
.B2(n_961),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1017),
.B(n_696),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_872),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_880),
.B(n_696),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1017),
.A2(n_891),
.B(n_1024),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_858),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_967),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_880),
.B(n_696),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_876),
.A2(n_874),
.B(n_873),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1017),
.B(n_696),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1017),
.B(n_696),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_891),
.A2(n_1017),
.B(n_879),
.Y(n_1131)
);

AND3x4_ASAP7_75t_L g1132 ( 
.A(n_865),
.B(n_599),
.C(n_800),
.Y(n_1132)
);

NAND2xp33_ASAP7_75t_L g1133 ( 
.A(n_891),
.B(n_729),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1017),
.A2(n_891),
.B(n_1024),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_891),
.A2(n_1017),
.B(n_879),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_880),
.B(n_696),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_891),
.A2(n_1017),
.B(n_879),
.Y(n_1137)
);

NOR2x1_ASAP7_75t_L g1138 ( 
.A(n_969),
.B(n_915),
.Y(n_1138)
);

OAI22x1_ASAP7_75t_L g1139 ( 
.A1(n_898),
.A2(n_366),
.B1(n_462),
.B2(n_696),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_1018),
.B(n_696),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_872),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_849),
.Y(n_1142)
);

NOR2xp67_ASAP7_75t_L g1143 ( 
.A(n_997),
.B(n_565),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1017),
.A2(n_891),
.B(n_1024),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_880),
.B(n_696),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_SL g1146 ( 
.A(n_849),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1017),
.B(n_696),
.Y(n_1147)
);

AOI21xp33_ASAP7_75t_L g1148 ( 
.A1(n_946),
.A2(n_891),
.B(n_696),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_891),
.A2(n_1017),
.B(n_879),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1017),
.B(n_696),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_876),
.A2(n_874),
.B(n_873),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_849),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_853),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_SL g1154 ( 
.A1(n_971),
.A2(n_1008),
.B(n_955),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_891),
.A2(n_1017),
.B(n_879),
.Y(n_1155)
);

AO31x2_ASAP7_75t_L g1156 ( 
.A1(n_891),
.A2(n_1017),
.A3(n_950),
.B(n_820),
.Y(n_1156)
);

NAND2x1p5_ASAP7_75t_L g1157 ( 
.A(n_872),
.B(n_853),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_869),
.B(n_768),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_880),
.B(n_696),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_967),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_SL g1161 ( 
.A1(n_891),
.A2(n_861),
.B(n_871),
.Y(n_1161)
);

AO31x2_ASAP7_75t_L g1162 ( 
.A1(n_891),
.A2(n_1017),
.A3(n_950),
.B(n_820),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1017),
.B(n_696),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1017),
.B(n_696),
.Y(n_1164)
);

AO31x2_ASAP7_75t_L g1165 ( 
.A1(n_891),
.A2(n_1017),
.A3(n_950),
.B(n_820),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_849),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1017),
.A2(n_891),
.B(n_1024),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1017),
.A2(n_891),
.B(n_1024),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1117),
.B(n_1121),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1148),
.B(n_1030),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1027),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1120),
.A2(n_1066),
.B1(n_1163),
.B2(n_1164),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1133),
.A2(n_1120),
.B(n_1103),
.C(n_1037),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1079),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1045),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1129),
.B(n_1130),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1049),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1133),
.A2(n_1155),
.B(n_1116),
.C(n_1149),
.Y(n_1178)
);

O2A1O1Ixp5_ASAP7_75t_L g1179 ( 
.A1(n_1060),
.A2(n_1063),
.B(n_1135),
.C(n_1131),
.Y(n_1179)
);

OAI21xp33_ASAP7_75t_L g1180 ( 
.A1(n_1140),
.A2(n_1150),
.B(n_1147),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1076),
.A2(n_1115),
.B1(n_1064),
.B2(n_1097),
.Y(n_1181)
);

NAND2x1p5_ASAP7_75t_L g1182 ( 
.A(n_1084),
.B(n_1079),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1140),
.B(n_1065),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_1028),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1076),
.A2(n_1115),
.B1(n_1064),
.B2(n_1066),
.Y(n_1185)
);

BUFx12f_ASAP7_75t_L g1186 ( 
.A(n_1089),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1137),
.A2(n_1080),
.B(n_1063),
.C(n_1051),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1158),
.B(n_1050),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1087),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1033),
.B(n_1113),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1035),
.B(n_1123),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_1079),
.Y(n_1192)
);

BUFx12f_ASAP7_75t_L g1193 ( 
.A(n_1142),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_1042),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_SL g1195 ( 
.A1(n_1044),
.A2(n_1026),
.B(n_1167),
.C(n_1144),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1110),
.B(n_1127),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1136),
.B(n_1145),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1159),
.B(n_1042),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1070),
.B(n_1083),
.Y(n_1199)
);

INVxp67_ASAP7_75t_SL g1200 ( 
.A(n_1157),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1026),
.A2(n_1168),
.B(n_1167),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1158),
.B(n_1094),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1111),
.A2(n_1168),
.B(n_1118),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1100),
.B(n_1068),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1114),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1094),
.B(n_1082),
.Y(n_1206)
);

INVx1_ASAP7_75t_SL g1207 ( 
.A(n_1081),
.Y(n_1207)
);

NOR2x1_ASAP7_75t_SL g1208 ( 
.A(n_1079),
.B(n_1122),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_SL g1209 ( 
.A(n_1166),
.Y(n_1209)
);

INVx1_ASAP7_75t_SL g1210 ( 
.A(n_1166),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1041),
.Y(n_1211)
);

BUFx4_ASAP7_75t_R g1212 ( 
.A(n_1146),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1075),
.B(n_1080),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1122),
.Y(n_1214)
);

CKINVDCx8_ASAP7_75t_R g1215 ( 
.A(n_1050),
.Y(n_1215)
);

OR2x2_ASAP7_75t_L g1216 ( 
.A(n_1125),
.B(n_1152),
.Y(n_1216)
);

INVx5_ASAP7_75t_L g1217 ( 
.A(n_1122),
.Y(n_1217)
);

AO21x1_ASAP7_75t_L g1218 ( 
.A1(n_1085),
.A2(n_1090),
.B(n_1072),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1132),
.A2(n_1139),
.B1(n_1146),
.B2(n_1092),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1111),
.A2(n_1134),
.B(n_1144),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1043),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_1059),
.Y(n_1222)
);

OR2x6_ASAP7_75t_L g1223 ( 
.A(n_1122),
.B(n_1141),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1125),
.B(n_1078),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1056),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1118),
.B(n_1119),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1143),
.B(n_1067),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1108),
.B(n_1062),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1161),
.A2(n_1085),
.B1(n_1134),
.B2(n_1124),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1141),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1132),
.A2(n_1107),
.B1(n_1029),
.B2(n_1154),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1119),
.B(n_1124),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1090),
.A2(n_1107),
.B1(n_1077),
.B2(n_1074),
.Y(n_1233)
);

OA21x2_ASAP7_75t_L g1234 ( 
.A1(n_1057),
.A2(n_1053),
.B(n_1039),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1126),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1160),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1141),
.Y(n_1237)
);

INVx1_ASAP7_75t_SL g1238 ( 
.A(n_1096),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1156),
.B(n_1165),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1157),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1099),
.A2(n_1048),
.B1(n_1058),
.B2(n_1098),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1036),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1138),
.B(n_1153),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1106),
.A2(n_1091),
.B1(n_1088),
.B2(n_1093),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1156),
.B(n_1165),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1071),
.A2(n_1104),
.B(n_1095),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1156),
.B(n_1165),
.Y(n_1247)
);

INVxp67_ASAP7_75t_L g1248 ( 
.A(n_1036),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1071),
.A2(n_1095),
.B(n_1073),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1059),
.A2(n_1061),
.B1(n_1096),
.B2(n_1112),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1112),
.A2(n_1040),
.B1(n_1105),
.B2(n_1055),
.Y(n_1251)
);

INVx2_ASAP7_75t_SL g1252 ( 
.A(n_1059),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1156),
.B(n_1165),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1162),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1162),
.B(n_1059),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1162),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1059),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1032),
.Y(n_1258)
);

INVxp67_ASAP7_75t_L g1259 ( 
.A(n_1061),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1162),
.B(n_1109),
.Y(n_1260)
);

OAI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1031),
.A2(n_1046),
.B1(n_1052),
.B2(n_1102),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1047),
.A2(n_1101),
.B(n_1038),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1086),
.B(n_1069),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1054),
.B(n_1034),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1128),
.Y(n_1265)
);

AOI21xp33_ASAP7_75t_SL g1266 ( 
.A1(n_1046),
.A2(n_1151),
.B(n_1052),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_SL g1267 ( 
.A1(n_1030),
.A2(n_946),
.B(n_1148),
.C(n_820),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1117),
.B(n_1121),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1042),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1030),
.A2(n_891),
.B(n_1148),
.C(n_946),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1033),
.B(n_1113),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1117),
.B(n_1121),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1045),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1033),
.B(n_1113),
.Y(n_1274)
);

BUFx2_ASAP7_75t_SL g1275 ( 
.A(n_1146),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1028),
.Y(n_1276)
);

INVxp67_ASAP7_75t_L g1277 ( 
.A(n_1113),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1148),
.B(n_891),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1117),
.B(n_1121),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1028),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1117),
.B(n_1121),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1113),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1158),
.B(n_1050),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1116),
.A2(n_1135),
.B(n_1131),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1033),
.B(n_1113),
.Y(n_1285)
);

INVx2_ASAP7_75t_SL g1286 ( 
.A(n_1089),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_SL g1287 ( 
.A1(n_1132),
.A2(n_898),
.B1(n_635),
.B2(n_462),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_1096),
.Y(n_1288)
);

AOI221x1_ASAP7_75t_L g1289 ( 
.A1(n_1030),
.A2(n_891),
.B1(n_1148),
.B2(n_1037),
.C(n_1161),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1158),
.B(n_1050),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1117),
.B(n_1121),
.Y(n_1291)
);

AOI21xp33_ASAP7_75t_SL g1292 ( 
.A1(n_1030),
.A2(n_462),
.B(n_898),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1033),
.B(n_1113),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1117),
.B(n_1121),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1028),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1045),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1117),
.B(n_1121),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1148),
.A2(n_891),
.B(n_1120),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1117),
.B(n_1121),
.Y(n_1299)
);

AO21x2_ASAP7_75t_L g1300 ( 
.A1(n_1029),
.A2(n_1154),
.B(n_891),
.Y(n_1300)
);

BUFx3_ASAP7_75t_L g1301 ( 
.A(n_1042),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1120),
.A2(n_891),
.B1(n_1030),
.B2(n_1066),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1033),
.B(n_1113),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1033),
.B(n_1113),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_1079),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1030),
.B(n_696),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_1079),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1116),
.A2(n_1135),
.B(n_1131),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1030),
.B(n_696),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1120),
.A2(n_1133),
.B1(n_1030),
.B2(n_1037),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1117),
.B(n_1121),
.Y(n_1311)
);

O2A1O1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1030),
.A2(n_891),
.B(n_1148),
.C(n_946),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_1096),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_1028),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1045),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1033),
.B(n_1113),
.Y(n_1316)
);

AO21x2_ASAP7_75t_L g1317 ( 
.A1(n_1262),
.A2(n_1298),
.B(n_1249),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1310),
.A2(n_1183),
.B1(n_1268),
.B2(n_1306),
.Y(n_1318)
);

NOR2x1_ASAP7_75t_R g1319 ( 
.A(n_1288),
.B(n_1275),
.Y(n_1319)
);

INVxp67_ASAP7_75t_L g1320 ( 
.A(n_1196),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1207),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1287),
.A2(n_1306),
.B1(n_1309),
.B2(n_1302),
.Y(n_1322)
);

NAND2x1p5_ASAP7_75t_L g1323 ( 
.A(n_1217),
.B(n_1228),
.Y(n_1323)
);

BUFx12f_ASAP7_75t_L g1324 ( 
.A(n_1186),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_SL g1325 ( 
.A1(n_1309),
.A2(n_1199),
.B1(n_1172),
.B2(n_1213),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1194),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1177),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1212),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1189),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1169),
.B(n_1176),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_SL g1331 ( 
.A(n_1194),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1201),
.A2(n_1220),
.B(n_1203),
.Y(n_1332)
);

OAI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1292),
.A2(n_1294),
.B1(n_1281),
.B2(n_1311),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1205),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_1313),
.Y(n_1335)
);

AOI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1219),
.A2(n_1180),
.B1(n_1310),
.B2(n_1170),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1273),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1296),
.Y(n_1338)
);

AO21x1_ASAP7_75t_SL g1339 ( 
.A1(n_1185),
.A2(n_1181),
.B(n_1256),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1173),
.B(n_1185),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1257),
.Y(n_1341)
);

CKINVDCx6p67_ASAP7_75t_R g1342 ( 
.A(n_1209),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1246),
.A2(n_1263),
.B(n_1251),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1315),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1272),
.A2(n_1279),
.B1(n_1291),
.B2(n_1297),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1170),
.A2(n_1278),
.B1(n_1181),
.B2(n_1284),
.Y(n_1346)
);

BUFx2_ASAP7_75t_R g1347 ( 
.A(n_1215),
.Y(n_1347)
);

INVx3_ASAP7_75t_L g1348 ( 
.A(n_1257),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1299),
.B(n_1191),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1217),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1173),
.B(n_1245),
.Y(n_1351)
);

CKINVDCx11_ASAP7_75t_R g1352 ( 
.A(n_1238),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1175),
.Y(n_1353)
);

NAND2x1p5_ASAP7_75t_L g1354 ( 
.A(n_1217),
.B(n_1228),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_SL g1355 ( 
.A1(n_1229),
.A2(n_1282),
.B1(n_1233),
.B2(n_1308),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1269),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_1184),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1198),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1269),
.Y(n_1359)
);

INVx1_ASAP7_75t_SL g1360 ( 
.A(n_1190),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_SL g1361 ( 
.A1(n_1270),
.A2(n_1312),
.B(n_1250),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1282),
.A2(n_1260),
.B1(n_1285),
.B2(n_1316),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1265),
.A2(n_1232),
.B(n_1226),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1276),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1258),
.A2(n_1241),
.B(n_1179),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1301),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1231),
.B(n_1271),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1258),
.A2(n_1179),
.B(n_1218),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1236),
.Y(n_1369)
);

OR2x6_ASAP7_75t_L g1370 ( 
.A(n_1178),
.B(n_1204),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1221),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1225),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1235),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1231),
.B(n_1304),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1234),
.A2(n_1204),
.B(n_1244),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1274),
.A2(n_1303),
.B1(n_1293),
.B2(n_1209),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1171),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1211),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1230),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_1230),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_SL g1381 ( 
.A1(n_1224),
.A2(n_1197),
.B1(n_1227),
.B2(n_1210),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1224),
.A2(n_1295),
.B1(n_1280),
.B2(n_1300),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1188),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_SL g1384 ( 
.A1(n_1300),
.A2(n_1314),
.B1(n_1277),
.B2(n_1193),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_SL g1385 ( 
.A1(n_1289),
.A2(n_1283),
.B1(n_1290),
.B2(n_1188),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_1286),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1230),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1206),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1248),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1283),
.B(n_1290),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1248),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1254),
.A2(n_1239),
.B1(n_1247),
.B2(n_1253),
.Y(n_1392)
);

INVx4_ASAP7_75t_L g1393 ( 
.A(n_1223),
.Y(n_1393)
);

AO21x1_ASAP7_75t_L g1394 ( 
.A1(n_1255),
.A2(n_1261),
.B(n_1266),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1259),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1240),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1240),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1259),
.Y(n_1398)
);

INVx2_ASAP7_75t_SL g1399 ( 
.A(n_1237),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1178),
.B(n_1187),
.Y(n_1400)
);

AO21x1_ASAP7_75t_SL g1401 ( 
.A1(n_1202),
.A2(n_1216),
.B(n_1267),
.Y(n_1401)
);

INVx1_ASAP7_75t_SL g1402 ( 
.A(n_1212),
.Y(n_1402)
);

AO21x2_ASAP7_75t_L g1403 ( 
.A1(n_1261),
.A2(n_1195),
.B(n_1267),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1242),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1187),
.A2(n_1182),
.B(n_1243),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1223),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1174),
.Y(n_1407)
);

INVx6_ASAP7_75t_L g1408 ( 
.A(n_1305),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1305),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1182),
.A2(n_1200),
.B1(n_1252),
.B2(n_1192),
.Y(n_1410)
);

AO21x1_ASAP7_75t_SL g1411 ( 
.A1(n_1208),
.A2(n_1195),
.B(n_1200),
.Y(n_1411)
);

OAI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1214),
.A2(n_1030),
.B1(n_981),
.B2(n_984),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1307),
.B(n_1264),
.Y(n_1413)
);

CKINVDCx20_ASAP7_75t_R g1414 ( 
.A(n_1307),
.Y(n_1414)
);

INVx5_ASAP7_75t_L g1415 ( 
.A(n_1257),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1270),
.A2(n_891),
.B(n_1030),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1298),
.A2(n_1030),
.B1(n_1120),
.B2(n_1133),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1282),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1298),
.A2(n_1030),
.B1(n_1120),
.B2(n_1133),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1222),
.B(n_1228),
.Y(n_1420)
);

INVx3_ASAP7_75t_SL g1421 ( 
.A(n_1288),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1177),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1310),
.A2(n_1120),
.B1(n_891),
.B2(n_898),
.Y(n_1423)
);

INVxp67_ASAP7_75t_SL g1424 ( 
.A(n_1282),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1198),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1395),
.B(n_1398),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1395),
.B(n_1398),
.Y(n_1427)
);

AOI222xp33_ASAP7_75t_L g1428 ( 
.A1(n_1423),
.A2(n_1416),
.B1(n_1419),
.B2(n_1417),
.C1(n_1318),
.C2(n_1340),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1386),
.Y(n_1429)
);

AO21x2_ASAP7_75t_L g1430 ( 
.A1(n_1361),
.A2(n_1403),
.B(n_1343),
.Y(n_1430)
);

BUFx4_ASAP7_75t_R g1431 ( 
.A(n_1383),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1386),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1353),
.Y(n_1433)
);

OA21x2_ASAP7_75t_L g1434 ( 
.A1(n_1375),
.A2(n_1332),
.B(n_1368),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1351),
.B(n_1400),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1418),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1351),
.B(n_1400),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1367),
.B(n_1374),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1345),
.B(n_1349),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1326),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1392),
.B(n_1370),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1417),
.A2(n_1419),
.B(n_1322),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1321),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1363),
.A2(n_1365),
.B(n_1394),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1392),
.B(n_1370),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1367),
.B(n_1374),
.Y(n_1446)
);

INVxp67_ASAP7_75t_L g1447 ( 
.A(n_1364),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1340),
.B(n_1355),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1333),
.A2(n_1325),
.B(n_1336),
.Y(n_1449)
);

INVx1_ASAP7_75t_SL g1450 ( 
.A(n_1360),
.Y(n_1450)
);

INVx1_ASAP7_75t_SL g1451 ( 
.A(n_1357),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1327),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1329),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1370),
.B(n_1346),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1420),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1334),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1424),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1420),
.B(n_1413),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1330),
.B(n_1320),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1388),
.B(n_1381),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1420),
.Y(n_1461)
);

INVxp67_ASAP7_75t_L g1462 ( 
.A(n_1358),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1390),
.B(n_1425),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1377),
.B(n_1378),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1366),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1337),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1338),
.Y(n_1467)
);

AO21x2_ASAP7_75t_L g1468 ( 
.A1(n_1403),
.A2(n_1317),
.B(n_1405),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1317),
.B(n_1362),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1396),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1344),
.B(n_1422),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1373),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1323),
.Y(n_1473)
);

BUFx8_ASAP7_75t_L g1474 ( 
.A(n_1331),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1373),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1371),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1372),
.Y(n_1477)
);

INVxp67_ASAP7_75t_L g1478 ( 
.A(n_1404),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1366),
.Y(n_1479)
);

AO21x2_ASAP7_75t_L g1480 ( 
.A1(n_1412),
.A2(n_1410),
.B(n_1406),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1414),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1339),
.B(n_1369),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_SL g1483 ( 
.A(n_1347),
.B(n_1328),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1323),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1397),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_1415),
.Y(n_1486)
);

AOI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1407),
.A2(n_1409),
.B(n_1389),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1391),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1354),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1356),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1382),
.B(n_1384),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1414),
.Y(n_1492)
);

INVxp67_ASAP7_75t_SL g1493 ( 
.A(n_1356),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1357),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1341),
.Y(n_1495)
);

INVxp67_ASAP7_75t_SL g1496 ( 
.A(n_1359),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1415),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1341),
.Y(n_1498)
);

OR2x2_ASAP7_75t_SL g1499 ( 
.A(n_1350),
.B(n_1408),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1469),
.B(n_1359),
.Y(n_1500)
);

INVxp67_ASAP7_75t_L g1501 ( 
.A(n_1470),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1430),
.B(n_1401),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1457),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1430),
.B(n_1411),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1430),
.B(n_1385),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1443),
.B(n_1421),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1435),
.B(n_1437),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1457),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1437),
.B(n_1376),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1426),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1427),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1427),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_1470),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1441),
.B(n_1402),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1433),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1468),
.B(n_1348),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1439),
.B(n_1393),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1468),
.B(n_1348),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1438),
.B(n_1393),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1445),
.B(n_1444),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1449),
.A2(n_1352),
.B1(n_1383),
.B2(n_1421),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1499),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1487),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1434),
.B(n_1387),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1446),
.B(n_1428),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1490),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1454),
.B(n_1399),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_L g1528 ( 
.A(n_1486),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1434),
.B(n_1387),
.Y(n_1529)
);

NOR2x1_ASAP7_75t_SL g1530 ( 
.A(n_1487),
.B(n_1415),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1499),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1434),
.B(n_1379),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1485),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1436),
.B(n_1342),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1434),
.B(n_1380),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1448),
.B(n_1380),
.Y(n_1536)
);

OAI221xp5_ASAP7_75t_L g1537 ( 
.A1(n_1521),
.A2(n_1442),
.B1(n_1460),
.B2(n_1491),
.C(n_1459),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1533),
.Y(n_1538)
);

OAI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1525),
.A2(n_1491),
.B1(n_1451),
.B2(n_1447),
.C(n_1462),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1526),
.B(n_1488),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1526),
.B(n_1488),
.Y(n_1541)
);

NAND2xp33_ASAP7_75t_L g1542 ( 
.A(n_1525),
.B(n_1328),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1507),
.B(n_1480),
.Y(n_1543)
);

OA211x2_ASAP7_75t_L g1544 ( 
.A1(n_1506),
.A2(n_1483),
.B(n_1478),
.C(n_1474),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1507),
.B(n_1480),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_SL g1546 ( 
.A1(n_1530),
.A2(n_1486),
.B(n_1497),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1517),
.B(n_1476),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1508),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1507),
.B(n_1480),
.Y(n_1549)
);

NAND3xp33_ASAP7_75t_L g1550 ( 
.A(n_1517),
.B(n_1474),
.C(n_1477),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1510),
.B(n_1450),
.Y(n_1551)
);

OAI221xp5_ASAP7_75t_SL g1552 ( 
.A1(n_1509),
.A2(n_1342),
.B1(n_1463),
.B2(n_1481),
.C(n_1492),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_SL g1553 ( 
.A1(n_1522),
.A2(n_1481),
.B1(n_1492),
.B2(n_1494),
.Y(n_1553)
);

AND2x2_ASAP7_75t_SL g1554 ( 
.A(n_1505),
.B(n_1431),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1527),
.B(n_1458),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1508),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1527),
.B(n_1458),
.Y(n_1557)
);

OAI221xp5_ASAP7_75t_SL g1558 ( 
.A1(n_1509),
.A2(n_1494),
.B1(n_1482),
.B2(n_1429),
.C(n_1432),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1534),
.B(n_1455),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1509),
.A2(n_1458),
.B1(n_1455),
.B2(n_1461),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1511),
.B(n_1512),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1527),
.B(n_1482),
.Y(n_1562)
);

NAND3xp33_ASAP7_75t_L g1563 ( 
.A(n_1523),
.B(n_1489),
.C(n_1474),
.Y(n_1563)
);

NAND3xp33_ASAP7_75t_L g1564 ( 
.A(n_1523),
.B(n_1489),
.C(n_1472),
.Y(n_1564)
);

INVxp67_ASAP7_75t_L g1565 ( 
.A(n_1534),
.Y(n_1565)
);

OAI221xp5_ASAP7_75t_SL g1566 ( 
.A1(n_1505),
.A2(n_1429),
.B1(n_1432),
.B2(n_1464),
.C(n_1496),
.Y(n_1566)
);

OAI221xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1505),
.A2(n_1493),
.B1(n_1471),
.B2(n_1453),
.C(n_1467),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1522),
.A2(n_1331),
.B1(n_1484),
.B2(n_1473),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1512),
.B(n_1475),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1519),
.B(n_1515),
.Y(n_1570)
);

NAND3xp33_ASAP7_75t_L g1571 ( 
.A(n_1514),
.B(n_1452),
.C(n_1456),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1515),
.B(n_1466),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1533),
.Y(n_1573)
);

NAND3xp33_ASAP7_75t_L g1574 ( 
.A(n_1514),
.B(n_1471),
.C(n_1495),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1531),
.A2(n_1455),
.B1(n_1461),
.B2(n_1352),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1531),
.A2(n_1331),
.B1(n_1484),
.B2(n_1473),
.Y(n_1576)
);

NAND3xp33_ASAP7_75t_L g1577 ( 
.A(n_1520),
.B(n_1498),
.C(n_1495),
.Y(n_1577)
);

OAI21xp5_ASAP7_75t_SL g1578 ( 
.A1(n_1502),
.A2(n_1473),
.B(n_1484),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1531),
.B(n_1455),
.Y(n_1579)
);

NAND2x1p5_ASAP7_75t_L g1580 ( 
.A(n_1554),
.B(n_1503),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1543),
.B(n_1516),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1538),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1545),
.B(n_1501),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1538),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1573),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1545),
.B(n_1520),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1549),
.B(n_1501),
.Y(n_1587)
);

INVx3_ASAP7_75t_L g1588 ( 
.A(n_1573),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1548),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1549),
.B(n_1503),
.Y(n_1590)
);

NOR2xp67_ASAP7_75t_L g1591 ( 
.A(n_1577),
.B(n_1520),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1556),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1577),
.B(n_1529),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1570),
.B(n_1500),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1554),
.B(n_1461),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1572),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1564),
.Y(n_1597)
);

AND2x4_ASAP7_75t_SL g1598 ( 
.A(n_1562),
.B(n_1528),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1555),
.B(n_1518),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1561),
.B(n_1547),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1555),
.B(n_1518),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1557),
.B(n_1565),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1569),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1540),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1554),
.B(n_1504),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1541),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1574),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1578),
.B(n_1504),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1574),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1571),
.Y(n_1610)
);

BUFx2_ASAP7_75t_L g1611 ( 
.A(n_1580),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1593),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1584),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1593),
.Y(n_1614)
);

INVx3_ASAP7_75t_L g1615 ( 
.A(n_1593),
.Y(n_1615)
);

INVxp67_ASAP7_75t_SL g1616 ( 
.A(n_1610),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1598),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1593),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1581),
.B(n_1504),
.Y(n_1619)
);

NOR2x1p5_ASAP7_75t_L g1620 ( 
.A(n_1605),
.B(n_1550),
.Y(n_1620)
);

INVx2_ASAP7_75t_SL g1621 ( 
.A(n_1598),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1608),
.B(n_1532),
.Y(n_1622)
);

OAI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1580),
.A2(n_1537),
.B1(n_1539),
.B2(n_1550),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1582),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1584),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1607),
.B(n_1571),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1607),
.B(n_1524),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1607),
.B(n_1609),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1608),
.B(n_1535),
.Y(n_1629)
);

OAI221xp5_ASAP7_75t_SL g1630 ( 
.A1(n_1597),
.A2(n_1575),
.B1(n_1563),
.B2(n_1560),
.C(n_1536),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1609),
.B(n_1551),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1588),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1588),
.Y(n_1633)
);

AOI211xp5_ASAP7_75t_L g1634 ( 
.A1(n_1597),
.A2(n_1542),
.B(n_1552),
.C(n_1566),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1582),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1588),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1603),
.B(n_1513),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1586),
.B(n_1524),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1585),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1600),
.B(n_1542),
.Y(n_1640)
);

AND2x2_ASAP7_75t_SL g1641 ( 
.A(n_1605),
.B(n_1513),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1584),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1624),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1641),
.B(n_1599),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1624),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1641),
.B(n_1601),
.Y(n_1646)
);

OAI21xp33_ASAP7_75t_L g1647 ( 
.A1(n_1616),
.A2(n_1580),
.B(n_1595),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1611),
.B(n_1591),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1635),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1640),
.B(n_1606),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1640),
.B(n_1606),
.Y(n_1651)
);

INVx1_ASAP7_75t_SL g1652 ( 
.A(n_1641),
.Y(n_1652)
);

OAI32xp33_ASAP7_75t_L g1653 ( 
.A1(n_1626),
.A2(n_1590),
.A3(n_1583),
.B1(n_1587),
.B2(n_1604),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1635),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1631),
.B(n_1324),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1639),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1639),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1637),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1626),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1631),
.B(n_1604),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1626),
.B(n_1583),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1616),
.B(n_1602),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1628),
.B(n_1587),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1632),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1632),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1634),
.B(n_1602),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1628),
.B(n_1590),
.Y(n_1667)
);

OAI21xp33_ASAP7_75t_L g1668 ( 
.A1(n_1634),
.A2(n_1558),
.B(n_1600),
.Y(n_1668)
);

BUFx2_ASAP7_75t_L g1669 ( 
.A(n_1641),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1628),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1611),
.B(n_1591),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1632),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1637),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1632),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1633),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1627),
.B(n_1612),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1633),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1627),
.B(n_1594),
.Y(n_1678)
);

OAI21xp33_ASAP7_75t_L g1679 ( 
.A1(n_1630),
.A2(n_1567),
.B(n_1596),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1611),
.B(n_1601),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1613),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1613),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1613),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1633),
.Y(n_1684)
);

INVxp67_ASAP7_75t_L g1685 ( 
.A(n_1620),
.Y(n_1685)
);

INVxp67_ASAP7_75t_SL g1686 ( 
.A(n_1669),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1669),
.B(n_1644),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1676),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1655),
.B(n_1324),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1643),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1659),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1643),
.Y(n_1692)
);

BUFx12f_ASAP7_75t_L g1693 ( 
.A(n_1648),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1654),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1652),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1661),
.B(n_1627),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1654),
.Y(n_1697)
);

INVx1_ASAP7_75t_SL g1698 ( 
.A(n_1650),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1656),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1644),
.B(n_1615),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1668),
.B(n_1620),
.Y(n_1701)
);

BUFx2_ASAP7_75t_L g1702 ( 
.A(n_1685),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1656),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1666),
.B(n_1622),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1647),
.B(n_1623),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1657),
.Y(n_1706)
);

AOI22x1_ASAP7_75t_L g1707 ( 
.A1(n_1648),
.A2(n_1615),
.B1(n_1623),
.B2(n_1612),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1646),
.B(n_1615),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1679),
.A2(n_1630),
.B1(n_1553),
.B2(n_1544),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1676),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1651),
.A2(n_1553),
.B1(n_1544),
.B2(n_1568),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1646),
.B(n_1680),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1680),
.B(n_1615),
.Y(n_1713)
);

INVx4_ASAP7_75t_L g1714 ( 
.A(n_1648),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1657),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1671),
.B(n_1615),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_1662),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1658),
.B(n_1622),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1645),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_SL g1720 ( 
.A1(n_1653),
.A2(n_1614),
.B1(n_1618),
.B2(n_1612),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1664),
.Y(n_1721)
);

AOI21xp33_ASAP7_75t_L g1722 ( 
.A1(n_1701),
.A2(n_1670),
.B(n_1661),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1709),
.B(n_1711),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1695),
.B(n_1673),
.Y(n_1724)
);

INVxp67_ASAP7_75t_L g1725 ( 
.A(n_1691),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1690),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1705),
.A2(n_1671),
.B1(n_1660),
.B2(n_1618),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1714),
.B(n_1671),
.Y(n_1728)
);

NAND4xp25_ASAP7_75t_L g1729 ( 
.A(n_1702),
.B(n_1653),
.C(n_1667),
.D(n_1663),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1711),
.A2(n_1693),
.B1(n_1687),
.B2(n_1695),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1702),
.B(n_1663),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1714),
.Y(n_1732)
);

OAI21xp33_ASAP7_75t_L g1733 ( 
.A1(n_1687),
.A2(n_1667),
.B(n_1614),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1689),
.B(n_1335),
.Y(n_1734)
);

NOR2x1p5_ASAP7_75t_SL g1735 ( 
.A(n_1688),
.B(n_1664),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1712),
.B(n_1619),
.Y(n_1736)
);

INVxp67_ASAP7_75t_L g1737 ( 
.A(n_1686),
.Y(n_1737)
);

O2A1O1Ixp33_ASAP7_75t_L g1738 ( 
.A1(n_1698),
.A2(n_1612),
.B(n_1614),
.C(n_1618),
.Y(n_1738)
);

OAI21xp33_ASAP7_75t_L g1739 ( 
.A1(n_1720),
.A2(n_1618),
.B(n_1614),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1712),
.B(n_1619),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1717),
.B(n_1622),
.Y(n_1741)
);

NAND2x1_ASAP7_75t_L g1742 ( 
.A(n_1714),
.B(n_1617),
.Y(n_1742)
);

AOI22x1_ASAP7_75t_L g1743 ( 
.A1(n_1693),
.A2(n_1621),
.B1(n_1617),
.B2(n_1678),
.Y(n_1743)
);

INVx1_ASAP7_75t_SL g1744 ( 
.A(n_1693),
.Y(n_1744)
);

OAI221xp5_ASAP7_75t_L g1745 ( 
.A1(n_1707),
.A2(n_1617),
.B1(n_1621),
.B2(n_1678),
.C(n_1649),
.Y(n_1745)
);

OAI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1707),
.A2(n_1621),
.B1(n_1576),
.B2(n_1638),
.Y(n_1746)
);

AOI222xp33_ASAP7_75t_L g1747 ( 
.A1(n_1717),
.A2(n_1704),
.B1(n_1708),
.B2(n_1700),
.C1(n_1718),
.C2(n_1719),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1728),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1726),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1737),
.B(n_1719),
.Y(n_1750)
);

NOR2x1p5_ASAP7_75t_L g1751 ( 
.A(n_1731),
.B(n_1742),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1744),
.B(n_1714),
.Y(n_1752)
);

OAI21xp33_ASAP7_75t_SL g1753 ( 
.A1(n_1729),
.A2(n_1708),
.B(n_1700),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1724),
.B(n_1696),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1725),
.B(n_1744),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1729),
.B(n_1696),
.Y(n_1756)
);

INVxp67_ASAP7_75t_SL g1757 ( 
.A(n_1728),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1732),
.Y(n_1758)
);

INVxp67_ASAP7_75t_L g1759 ( 
.A(n_1743),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1730),
.A2(n_1713),
.B1(n_1716),
.B2(n_1710),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1736),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1740),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1747),
.B(n_1688),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1741),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1722),
.B(n_1688),
.Y(n_1765)
);

NAND2x1_ASAP7_75t_L g1766 ( 
.A(n_1727),
.B(n_1716),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1723),
.B(n_1733),
.Y(n_1767)
);

NOR3x1_ASAP7_75t_L g1768 ( 
.A(n_1757),
.B(n_1745),
.C(n_1692),
.Y(n_1768)
);

BUFx6f_ASAP7_75t_SL g1769 ( 
.A(n_1758),
.Y(n_1769)
);

OAI221xp5_ASAP7_75t_SL g1770 ( 
.A1(n_1759),
.A2(n_1746),
.B1(n_1739),
.B2(n_1738),
.C(n_1710),
.Y(n_1770)
);

NAND2xp67_ASAP7_75t_SL g1771 ( 
.A(n_1752),
.B(n_1713),
.Y(n_1771)
);

NAND2xp33_ASAP7_75t_R g1772 ( 
.A(n_1755),
.B(n_1734),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1767),
.B(n_1710),
.Y(n_1773)
);

NAND3xp33_ASAP7_75t_L g1774 ( 
.A(n_1760),
.B(n_1692),
.C(n_1690),
.Y(n_1774)
);

AOI21xp5_ASAP7_75t_L g1775 ( 
.A1(n_1763),
.A2(n_1766),
.B(n_1765),
.Y(n_1775)
);

AOI221xp5_ASAP7_75t_L g1776 ( 
.A1(n_1760),
.A2(n_1706),
.B1(n_1697),
.B2(n_1699),
.C(n_1715),
.Y(n_1776)
);

XNOR2x1_ASAP7_75t_L g1777 ( 
.A(n_1756),
.B(n_1735),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1754),
.Y(n_1778)
);

O2A1O1Ixp33_ASAP7_75t_L g1779 ( 
.A1(n_1765),
.A2(n_1694),
.B(n_1715),
.C(n_1706),
.Y(n_1779)
);

NOR3xp33_ASAP7_75t_L g1780 ( 
.A(n_1775),
.B(n_1773),
.C(n_1778),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1769),
.Y(n_1781)
);

NOR3xp33_ASAP7_75t_L g1782 ( 
.A(n_1770),
.B(n_1748),
.C(n_1750),
.Y(n_1782)
);

NOR3x1_ASAP7_75t_L g1783 ( 
.A(n_1774),
.B(n_1750),
.C(n_1764),
.Y(n_1783)
);

NAND3xp33_ASAP7_75t_L g1784 ( 
.A(n_1777),
.B(n_1753),
.C(n_1749),
.Y(n_1784)
);

NAND2xp33_ASAP7_75t_SL g1785 ( 
.A(n_1769),
.B(n_1751),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1779),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1768),
.B(n_1761),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1776),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1771),
.B(n_1762),
.Y(n_1789)
);

AND5x1_ASAP7_75t_L g1790 ( 
.A(n_1772),
.B(n_1721),
.C(n_1703),
.D(n_1699),
.E(n_1697),
.Y(n_1790)
);

NAND3xp33_ASAP7_75t_L g1791 ( 
.A(n_1780),
.B(n_1703),
.C(n_1694),
.Y(n_1791)
);

NAND3xp33_ASAP7_75t_SL g1792 ( 
.A(n_1785),
.B(n_1335),
.C(n_1721),
.Y(n_1792)
);

OAI222xp33_ASAP7_75t_L g1793 ( 
.A1(n_1788),
.A2(n_1721),
.B1(n_1684),
.B2(n_1672),
.C1(n_1674),
.C2(n_1675),
.Y(n_1793)
);

A2O1A1Ixp33_ASAP7_75t_L g1794 ( 
.A1(n_1784),
.A2(n_1681),
.B(n_1682),
.C(n_1683),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1781),
.B(n_1629),
.Y(n_1795)
);

O2A1O1Ixp33_ASAP7_75t_L g1796 ( 
.A1(n_1786),
.A2(n_1683),
.B(n_1684),
.C(n_1677),
.Y(n_1796)
);

NOR4xp75_ASAP7_75t_L g1797 ( 
.A(n_1787),
.B(n_1579),
.C(n_1559),
.D(n_1319),
.Y(n_1797)
);

NOR2xp67_ASAP7_75t_L g1798 ( 
.A(n_1792),
.B(n_1789),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1795),
.A2(n_1782),
.B1(n_1783),
.B2(n_1790),
.Y(n_1799)
);

AOI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1791),
.A2(n_1794),
.B1(n_1797),
.B2(n_1672),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1796),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1793),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1795),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1795),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1802),
.B(n_1677),
.Y(n_1805)
);

OAI211xp5_ASAP7_75t_L g1806 ( 
.A1(n_1799),
.A2(n_1675),
.B(n_1674),
.C(n_1665),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1801),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1803),
.B(n_1665),
.Y(n_1808)
);

NOR2xp67_ASAP7_75t_SL g1809 ( 
.A(n_1804),
.B(n_1440),
.Y(n_1809)
);

AOI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1807),
.A2(n_1798),
.B1(n_1800),
.B2(n_1629),
.Y(n_1810)
);

NOR2xp67_ASAP7_75t_SL g1811 ( 
.A(n_1805),
.B(n_1440),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1808),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1810),
.Y(n_1813)
);

AOI211xp5_ASAP7_75t_L g1814 ( 
.A1(n_1813),
.A2(n_1812),
.B(n_1811),
.C(n_1809),
.Y(n_1814)
);

AOI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1814),
.A2(n_1806),
.B(n_1636),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1814),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1816),
.A2(n_1633),
.B1(n_1636),
.B2(n_1589),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1815),
.B(n_1636),
.Y(n_1818)
);

AOI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1817),
.A2(n_1818),
.B1(n_1636),
.B2(n_1629),
.Y(n_1819)
);

OAI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1818),
.A2(n_1592),
.B(n_1619),
.Y(n_1820)
);

OAI21xp5_ASAP7_75t_SL g1821 ( 
.A1(n_1819),
.A2(n_1350),
.B(n_1592),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1821),
.A2(n_1820),
.B1(n_1589),
.B2(n_1625),
.Y(n_1822)
);

AOI221xp5_ASAP7_75t_L g1823 ( 
.A1(n_1822),
.A2(n_1642),
.B1(n_1625),
.B2(n_1585),
.C(n_1588),
.Y(n_1823)
);

AOI211xp5_ASAP7_75t_L g1824 ( 
.A1(n_1823),
.A2(n_1546),
.B(n_1479),
.C(n_1465),
.Y(n_1824)
);


endmodule