module fake_netlist_1_8168_n_31 (n_1, n_2, n_4, n_3, n_0, n_31);
input n_1;
input n_2;
input n_4;
input n_3;
input n_0;
output n_31;
wire n_20;
wire n_5;
wire n_23;
wire n_8;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_6;
wire n_29;
wire n_7;
wire n_27;
CKINVDCx20_ASAP7_75t_R g5 ( .A(n_1), .Y(n_5) );
BUFx3_ASAP7_75t_L g6 ( .A(n_4), .Y(n_6) );
INVx2_ASAP7_75t_L g7 ( .A(n_0), .Y(n_7) );
HB1xp67_ASAP7_75t_L g8 ( .A(n_2), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_3), .Y(n_9) );
NAND2xp5_ASAP7_75t_SL g10 ( .A(n_8), .B(n_0), .Y(n_10) );
AOI21xp5_ASAP7_75t_L g11 ( .A1(n_7), .A2(n_0), .B(n_1), .Y(n_11) );
AOI22xp5_ASAP7_75t_L g12 ( .A1(n_5), .A2(n_4), .B1(n_1), .B2(n_2), .Y(n_12) );
INVx1_ASAP7_75t_SL g13 ( .A(n_6), .Y(n_13) );
OAI22xp5_ASAP7_75t_L g14 ( .A1(n_6), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_11), .Y(n_15) );
AOI22xp33_ASAP7_75t_SL g16 ( .A1(n_14), .A2(n_7), .B1(n_9), .B2(n_4), .Y(n_16) );
NOR2xp33_ASAP7_75t_R g17 ( .A(n_13), .B(n_0), .Y(n_17) );
BUFx2_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_15), .B(n_10), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_15), .Y(n_20) );
OR2x2_ASAP7_75t_L g21 ( .A(n_18), .B(n_12), .Y(n_21) );
AOI222xp33_ASAP7_75t_L g22 ( .A1(n_20), .A2(n_18), .B1(n_9), .B2(n_16), .C1(n_17), .C2(n_2), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_19), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_21), .B(n_17), .Y(n_24) );
AOI221x1_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_16), .B1(n_4), .B2(n_3), .C(n_2), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
AOI21xp5_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_21), .B(n_18), .Y(n_27) );
NOR2x1_ASAP7_75t_L g28 ( .A(n_26), .B(n_27), .Y(n_28) );
HB1xp67_ASAP7_75t_L g29 ( .A(n_25), .Y(n_29) );
AOI22xp5_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_3), .B1(n_22), .B2(n_29), .Y(n_30) );
AOI22xp5_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_3), .B1(n_28), .B2(n_24), .Y(n_31) );
endmodule