module fake_netlist_6_4386_n_1877 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1877);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1877;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_20),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_58),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_115),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_40),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_4),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_5),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_92),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_120),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_42),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_159),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_100),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_140),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_168),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_28),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_107),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_122),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_131),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_45),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_87),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_53),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_53),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_156),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_134),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_93),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_19),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_104),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_137),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_83),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_73),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_89),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_60),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_16),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_39),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_44),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_103),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_88),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_117),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_148),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_160),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_116),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_158),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_102),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_109),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_46),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_20),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_144),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_57),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_129),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_29),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_37),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_170),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_44),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_3),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_48),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_147),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_59),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_18),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_9),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_47),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_17),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_141),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_121),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_45),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_94),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_32),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_74),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_78),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_46),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_99),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_27),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_58),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_146),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_56),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_155),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_138),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_139),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_172),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_166),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_23),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_55),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_28),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_63),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_9),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_95),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_27),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_114),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_6),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_18),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_22),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_66),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_164),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_0),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_124),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_80),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_22),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_37),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_97),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_167),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_106),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_135),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_40),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_2),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_136),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_130),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_47),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_108),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_61),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_151),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_38),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_52),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_149),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_142),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_65),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_56),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_125),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_111),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_62),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_75),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_38),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_86),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_30),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_50),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_59),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_67),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_112),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_98),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_82),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_84),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_12),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_79),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_174),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_6),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_127),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_96),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_91),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_54),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_64),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_90),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_55),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_54),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_152),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_35),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_35),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_157),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_77),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_15),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_17),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_15),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_0),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_169),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_101),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_69),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_50),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_7),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_31),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_12),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_21),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_118),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_123),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_49),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_57),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_39),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_41),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_11),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_8),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_16),
.Y(n_344)
);

BUFx10_ASAP7_75t_L g345 ( 
.A(n_49),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_41),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_14),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_182),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_300),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_187),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_R g351 ( 
.A(n_195),
.B(n_173),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_232),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_209),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_238),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_175),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_277),
.B(n_1),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_225),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_210),
.B(n_1),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_210),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_274),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_304),
.B(n_2),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_227),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_210),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_230),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_234),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_237),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_253),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_210),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_241),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_210),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_242),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_210),
.B(n_304),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_208),
.B(n_3),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_303),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_180),
.B(n_4),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_255),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_210),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_210),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_262),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_297),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_289),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_243),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_201),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_251),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_297),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_231),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_231),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_338),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_338),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_274),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_298),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_231),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_231),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_258),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_265),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_231),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_266),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_308),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_267),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_330),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_213),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_236),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_328),
.B(n_7),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_280),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_175),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_214),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_236),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_236),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_288),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_254),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_236),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_236),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_301),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_215),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_301),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_301),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_292),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_274),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_328),
.B(n_190),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_301),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_301),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_217),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_219),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_345),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_299),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g426 ( 
.A(n_254),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_344),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_307),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_220),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_224),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_229),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_344),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_310),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_347),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_344),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_374),
.Y(n_436)
);

INVx6_ASAP7_75t_L g437 ( 
.A(n_374),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_410),
.B(n_328),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_356),
.B(n_203),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_426),
.B(n_302),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_386),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_411),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_411),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_386),
.Y(n_444)
);

AND2x6_ASAP7_75t_L g445 ( 
.A(n_419),
.B(n_303),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_359),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_403),
.B(n_392),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_363),
.Y(n_448)
);

BUFx12f_ASAP7_75t_L g449 ( 
.A(n_349),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_361),
.B(n_203),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_393),
.B(n_344),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_387),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_387),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_368),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_396),
.B(n_344),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_402),
.Y(n_456)
);

OA21x2_ASAP7_75t_L g457 ( 
.A1(n_358),
.A2(n_342),
.B(n_235),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_407),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_408),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_377),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_373),
.B(n_203),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_412),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_413),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_374),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_355),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_415),
.B(n_302),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_416),
.B(n_177),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_420),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_374),
.Y(n_469)
);

AND2x6_ASAP7_75t_L g470 ( 
.A(n_374),
.B(n_303),
.Y(n_470)
);

OAI21x1_ASAP7_75t_L g471 ( 
.A1(n_372),
.A2(n_191),
.B(n_190),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_370),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_352),
.B(n_193),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_351),
.B(n_244),
.Y(n_474)
);

BUFx8_ASAP7_75t_L g475 ( 
.A(n_418),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_421),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_427),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_432),
.B(n_191),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_370),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_435),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_378),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_380),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_385),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_375),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_388),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_389),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_375),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_371),
.B(n_244),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_418),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_354),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_353),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_353),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_357),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_357),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_405),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_362),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_349),
.Y(n_497)
);

BUFx8_ASAP7_75t_L g498 ( 
.A(n_401),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_362),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_364),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_364),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_365),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_365),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_366),
.B(n_177),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_366),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_SL g506 ( 
.A(n_369),
.B(n_176),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_369),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_382),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_382),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_384),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_360),
.B(n_206),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_384),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_394),
.Y(n_513)
);

OR2x6_ASAP7_75t_L g514 ( 
.A(n_491),
.B(n_206),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_444),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_449),
.B(n_406),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_497),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_441),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_481),
.Y(n_519)
);

AND2x2_ASAP7_75t_SL g520 ( 
.A(n_457),
.B(n_240),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_441),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_436),
.Y(n_522)
);

OAI22xp33_ASAP7_75t_SL g523 ( 
.A1(n_450),
.A2(n_390),
.B1(n_424),
.B2(n_240),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_449),
.B(n_414),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_484),
.B(n_394),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_504),
.B(n_422),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_481),
.Y(n_527)
);

INVx6_ASAP7_75t_L g528 ( 
.A(n_466),
.Y(n_528)
);

NAND2xp33_ASAP7_75t_SL g529 ( 
.A(n_439),
.B(n_395),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g530 ( 
.A(n_472),
.Y(n_530)
);

INVx5_ASAP7_75t_L g531 ( 
.A(n_470),
.Y(n_531)
);

OR2x6_ASAP7_75t_L g532 ( 
.A(n_491),
.B(n_268),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_489),
.B(n_395),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_489),
.B(n_397),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_436),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_466),
.B(n_268),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_484),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_441),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_436),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_466),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_444),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_472),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_441),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_466),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_444),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_504),
.B(n_423),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_489),
.B(n_397),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_446),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_470),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_446),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_446),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_436),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_472),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_472),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_446),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_439),
.B(n_450),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_436),
.Y(n_557)
);

BUFx8_ASAP7_75t_SL g558 ( 
.A(n_449),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_472),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_489),
.B(n_399),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_436),
.Y(n_561)
);

NOR3xp33_ASAP7_75t_L g562 ( 
.A(n_461),
.B(n_383),
.C(n_399),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_448),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_448),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_484),
.B(n_404),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_448),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_484),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_448),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_479),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_454),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_436),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_454),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_489),
.B(n_404),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_473),
.B(n_409),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_438),
.B(n_409),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_454),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_454),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_L g578 ( 
.A(n_484),
.B(n_417),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_473),
.B(n_417),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_436),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_484),
.B(n_425),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_460),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_438),
.B(n_425),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_464),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_479),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_460),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_SL g587 ( 
.A(n_461),
.B(n_428),
.Y(n_587)
);

INVx5_ASAP7_75t_L g588 ( 
.A(n_470),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_438),
.B(n_428),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_506),
.A2(n_325),
.B1(n_211),
.B2(n_273),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_460),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_464),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_479),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_479),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_465),
.B(n_484),
.Y(n_595)
);

AND3x2_ASAP7_75t_L g596 ( 
.A(n_507),
.B(n_271),
.C(n_235),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_464),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_498),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_484),
.B(n_433),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_479),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_460),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_452),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_452),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_464),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_L g605 ( 
.A(n_493),
.B(n_434),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_453),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_466),
.B(n_271),
.Y(n_607)
);

BUFx4f_ASAP7_75t_L g608 ( 
.A(n_457),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_493),
.B(n_433),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_447),
.B(n_434),
.Y(n_610)
);

AND2x6_ASAP7_75t_L g611 ( 
.A(n_491),
.B(n_303),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_464),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_440),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_453),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_451),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_493),
.B(n_429),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_457),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_464),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_507),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_442),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_493),
.B(n_431),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_506),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_487),
.A2(n_430),
.B1(n_207),
.B2(n_245),
.Y(n_623)
);

BUFx4f_ASAP7_75t_L g624 ( 
.A(n_457),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_451),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_455),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_442),
.Y(n_627)
);

BUFx4f_ASAP7_75t_L g628 ( 
.A(n_457),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_447),
.B(n_233),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_498),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_464),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_464),
.Y(n_632)
);

NOR3xp33_ASAP7_75t_L g633 ( 
.A(n_488),
.B(n_261),
.C(n_246),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_L g634 ( 
.A(n_493),
.B(n_303),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_455),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_443),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_443),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_469),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_456),
.Y(n_639)
);

NAND3xp33_ASAP7_75t_L g640 ( 
.A(n_457),
.B(n_199),
.C(n_181),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_456),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_496),
.B(n_400),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_458),
.Y(n_643)
);

NAND3xp33_ASAP7_75t_L g644 ( 
.A(n_440),
.B(n_205),
.C(n_204),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_498),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_465),
.B(n_183),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_458),
.Y(n_647)
);

INVx4_ASAP7_75t_L g648 ( 
.A(n_470),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_493),
.B(n_244),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_437),
.Y(n_650)
);

AND2x6_ASAP7_75t_L g651 ( 
.A(n_491),
.B(n_212),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_459),
.Y(n_652)
);

OR2x6_ASAP7_75t_L g653 ( 
.A(n_492),
.B(n_216),
.Y(n_653)
);

BUFx10_ASAP7_75t_L g654 ( 
.A(n_493),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_459),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_462),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_440),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_495),
.A2(n_327),
.B1(n_279),
.B2(n_196),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_462),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_467),
.B(n_239),
.Y(n_660)
);

INVxp33_ASAP7_75t_L g661 ( 
.A(n_497),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_469),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_463),
.Y(n_663)
);

NAND2xp33_ASAP7_75t_L g664 ( 
.A(n_493),
.B(n_184),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_463),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_468),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_558),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_613),
.B(n_492),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_540),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_540),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_L g671 ( 
.A(n_651),
.B(n_499),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_657),
.B(n_540),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_556),
.B(n_492),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_615),
.B(n_625),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_610),
.B(n_492),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_615),
.B(n_494),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_544),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_625),
.B(n_494),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g679 ( 
.A1(n_640),
.A2(n_471),
.B(n_494),
.Y(n_679)
);

AOI21x1_ASAP7_75t_L g680 ( 
.A1(n_519),
.A2(n_471),
.B(n_467),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_626),
.B(n_494),
.Y(n_681)
);

NAND3xp33_ASAP7_75t_L g682 ( 
.A(n_575),
.B(n_501),
.C(n_496),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_L g683 ( 
.A(n_651),
.B(n_499),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_525),
.A2(n_505),
.B1(n_503),
.B2(n_500),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_626),
.B(n_500),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_515),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_544),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_635),
.B(n_500),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_520),
.A2(n_445),
.B1(n_487),
.B2(n_342),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_515),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_537),
.A2(n_471),
.B(n_500),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_583),
.B(n_503),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_525),
.B(n_499),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_635),
.B(n_503),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_565),
.B(n_499),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_565),
.B(n_499),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_581),
.A2(n_503),
.B1(n_505),
.B2(n_512),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_581),
.A2(n_505),
.B1(n_512),
.B2(n_502),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_515),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_544),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_599),
.B(n_505),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_641),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_599),
.B(n_499),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_523),
.B(n_499),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_537),
.B(n_499),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_523),
.B(n_513),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_567),
.B(n_513),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_567),
.B(n_513),
.Y(n_708)
);

AND2x6_ASAP7_75t_SL g709 ( 
.A(n_642),
.B(n_490),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_641),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_643),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_595),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_520),
.B(n_513),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_541),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_595),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_520),
.A2(n_445),
.B1(n_283),
.B2(n_248),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_589),
.B(n_501),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_619),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_528),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_629),
.B(n_513),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_643),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_652),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_646),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_519),
.B(n_513),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_646),
.Y(n_725)
);

BUFx5_ASAP7_75t_L g726 ( 
.A(n_617),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_L g727 ( 
.A(n_651),
.B(n_513),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_578),
.A2(n_512),
.B1(n_508),
.B2(n_502),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_652),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_654),
.B(n_513),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_527),
.B(n_512),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_527),
.B(n_512),
.Y(n_732)
);

INVxp33_ASAP7_75t_L g733 ( 
.A(n_661),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_596),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_528),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_655),
.B(n_482),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_533),
.Y(n_737)
);

NAND2xp33_ASAP7_75t_L g738 ( 
.A(n_651),
.B(n_508),
.Y(n_738)
);

INVx5_ASAP7_75t_L g739 ( 
.A(n_549),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_654),
.B(n_509),
.Y(n_740)
);

O2A1O1Ixp33_ASAP7_75t_L g741 ( 
.A1(n_664),
.A2(n_605),
.B(n_649),
.C(n_609),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_655),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_534),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_526),
.A2(n_510),
.B1(n_509),
.B2(n_507),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_530),
.B(n_510),
.Y(n_745)
);

OAI22xp33_ASAP7_75t_L g746 ( 
.A1(n_658),
.A2(n_495),
.B1(n_490),
.B2(n_270),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_663),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_546),
.B(n_511),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_663),
.B(n_482),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_654),
.B(n_475),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_665),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_562),
.B(n_475),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_633),
.B(n_475),
.Y(n_753)
);

BUFx6f_ASAP7_75t_SL g754 ( 
.A(n_651),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_665),
.Y(n_755)
);

AND2x4_ASAP7_75t_SL g756 ( 
.A(n_653),
.B(n_348),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_547),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_666),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_660),
.B(n_475),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_654),
.B(n_475),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_608),
.B(n_474),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_574),
.B(n_488),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_517),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_579),
.B(n_511),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_517),
.B(n_511),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_541),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_560),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_541),
.Y(n_768)
);

OR2x6_ASAP7_75t_L g769 ( 
.A(n_616),
.B(n_474),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_545),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_666),
.Y(n_771)
);

INVx4_ASAP7_75t_L g772 ( 
.A(n_528),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_636),
.B(n_637),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_545),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_622),
.B(n_483),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_636),
.B(n_637),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_623),
.B(n_483),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_573),
.B(n_486),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_639),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_598),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_639),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_587),
.A2(n_350),
.B1(n_367),
.B2(n_376),
.Y(n_782)
);

OR2x6_ASAP7_75t_L g783 ( 
.A(n_621),
.B(n_486),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_576),
.Y(n_784)
);

INVx4_ASAP7_75t_L g785 ( 
.A(n_528),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_608),
.B(n_218),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_647),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_644),
.B(n_184),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_542),
.B(n_445),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_608),
.B(n_221),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_644),
.B(n_529),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_658),
.B(n_379),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_542),
.B(n_445),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_576),
.Y(n_794)
);

AO221x1_ASAP7_75t_L g795 ( 
.A1(n_638),
.A2(n_257),
.B1(n_222),
.B2(n_223),
.C(n_228),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_624),
.B(n_226),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_536),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_653),
.B(n_185),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_656),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_653),
.A2(n_532),
.B1(n_514),
.B2(n_624),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_624),
.B(n_247),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_656),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_650),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_659),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_659),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_628),
.B(n_260),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_653),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_620),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_653),
.B(n_185),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_638),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_553),
.B(n_445),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_553),
.B(n_445),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_620),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_617),
.A2(n_445),
.B1(n_263),
.B2(n_259),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_536),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_554),
.B(n_445),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_630),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_640),
.A2(n_478),
.B(n_312),
.C(n_309),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_554),
.B(n_445),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_627),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_536),
.A2(n_381),
.B1(n_391),
.B2(n_398),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_628),
.B(n_264),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_559),
.B(n_445),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_514),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_536),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_627),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_577),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_559),
.B(n_569),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_602),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_603),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_675),
.B(n_516),
.Y(n_831)
);

NAND3xp33_ASAP7_75t_L g832 ( 
.A(n_762),
.B(n_498),
.C(n_524),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_693),
.A2(n_628),
.B(n_695),
.Y(n_833)
);

AND2x6_ASAP7_75t_L g834 ( 
.A(n_701),
.B(n_617),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_679),
.A2(n_585),
.B(n_569),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_693),
.A2(n_532),
.B(n_514),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_675),
.B(n_607),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_672),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_672),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_692),
.A2(n_607),
.B(n_585),
.C(n_593),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_692),
.B(n_607),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_701),
.B(n_549),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_765),
.Y(n_843)
);

NOR2x1_ASAP7_75t_L g844 ( 
.A(n_682),
.B(n_514),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_758),
.B(n_607),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_695),
.A2(n_532),
.B(n_514),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_673),
.A2(n_532),
.B1(n_600),
.B2(n_594),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_808),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_718),
.B(n_498),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_813),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_820),
.Y(n_851)
);

AOI21x1_ASAP7_75t_L g852 ( 
.A1(n_707),
.A2(n_594),
.B(n_593),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_668),
.B(n_651),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_810),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_748),
.B(n_651),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_696),
.A2(n_532),
.B(n_521),
.Y(n_856)
);

A2O1A1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_762),
.A2(n_600),
.B(n_518),
.C(n_521),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_696),
.A2(n_538),
.B(n_518),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_703),
.A2(n_543),
.B(n_538),
.Y(n_859)
);

NAND3xp33_ASAP7_75t_L g860 ( 
.A(n_717),
.B(n_645),
.C(n_634),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_717),
.B(n_549),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_826),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_723),
.B(n_485),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_669),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_730),
.A2(n_543),
.B(n_549),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_810),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_725),
.B(n_485),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_674),
.B(n_638),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_676),
.B(n_638),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_718),
.B(n_733),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_678),
.B(n_662),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_739),
.A2(n_648),
.B(n_552),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_739),
.A2(n_648),
.B(n_552),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_730),
.A2(n_648),
.B(n_550),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_712),
.A2(n_614),
.B(n_606),
.C(n_603),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_791),
.A2(n_662),
.B1(n_611),
.B2(n_648),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_725),
.B(n_485),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_681),
.B(n_662),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_786),
.A2(n_550),
.B(n_548),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_691),
.A2(n_790),
.B(n_786),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_685),
.B(n_601),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_790),
.A2(n_551),
.B(n_548),
.Y(n_882)
);

OAI21xp33_ASAP7_75t_L g883 ( 
.A1(n_777),
.A2(n_178),
.B(n_176),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_669),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_744),
.B(n_186),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_829),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_684),
.B(n_531),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_745),
.B(n_186),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_688),
.B(n_601),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_694),
.B(n_551),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_697),
.A2(n_269),
.B1(n_322),
.B2(n_319),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_763),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_698),
.B(n_531),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_SL g894 ( 
.A(n_780),
.B(n_281),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_716),
.A2(n_284),
.B1(n_305),
.B2(n_313),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_796),
.A2(n_563),
.B(n_555),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_712),
.B(n_555),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_830),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_791),
.A2(n_606),
.B(n_614),
.C(n_566),
.Y(n_899)
);

BUFx8_ASAP7_75t_SL g900 ( 
.A(n_667),
.Y(n_900)
);

BUFx4f_ASAP7_75t_L g901 ( 
.A(n_769),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_796),
.A2(n_564),
.B(n_563),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_801),
.A2(n_566),
.B(n_564),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_821),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_770),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_715),
.B(n_568),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_715),
.B(n_702),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_797),
.A2(n_611),
.B1(n_572),
.B2(n_568),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_779),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_710),
.B(n_570),
.Y(n_910)
);

BUFx2_ASAP7_75t_SL g911 ( 
.A(n_775),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_781),
.Y(n_912)
);

OAI321xp33_ASAP7_75t_L g913 ( 
.A1(n_746),
.A2(n_287),
.A3(n_249),
.B1(n_314),
.B2(n_318),
.C(n_320),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_711),
.B(n_570),
.Y(n_914)
);

A2O1A1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_788),
.A2(n_572),
.B(n_582),
.C(n_586),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_801),
.A2(n_582),
.B(n_586),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_721),
.B(n_591),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_769),
.B(n_189),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_737),
.B(n_189),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_774),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_743),
.B(n_192),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_788),
.A2(n_591),
.B(n_577),
.C(n_631),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_777),
.A2(n_631),
.B(n_632),
.C(n_580),
.Y(n_923)
);

O2A1O1Ixp5_ASAP7_75t_L g924 ( 
.A1(n_704),
.A2(n_631),
.B(n_632),
.C(n_561),
.Y(n_924)
);

NOR3xp33_ASAP7_75t_L g925 ( 
.A(n_746),
.B(n_329),
.C(n_202),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_806),
.A2(n_632),
.B(n_580),
.Y(n_926)
);

CKINVDCx20_ASAP7_75t_R g927 ( 
.A(n_817),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_686),
.Y(n_928)
);

BUFx12f_ASAP7_75t_L g929 ( 
.A(n_734),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_716),
.A2(n_329),
.B1(n_336),
.B2(n_323),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_764),
.B(n_345),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_736),
.Y(n_932)
);

OAI21xp33_ASAP7_75t_L g933 ( 
.A1(n_778),
.A2(n_324),
.B(n_339),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_736),
.B(n_331),
.Y(n_934)
);

AO21x1_ASAP7_75t_L g935 ( 
.A1(n_806),
.A2(n_478),
.B(n_333),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_728),
.B(n_531),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_739),
.A2(n_539),
.B(n_552),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_787),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_669),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_739),
.A2(n_708),
.B(n_705),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_799),
.Y(n_941)
);

AOI21xp33_ASAP7_75t_L g942 ( 
.A1(n_798),
.A2(n_196),
.B(n_194),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_722),
.B(n_522),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_729),
.B(n_522),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_669),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_706),
.A2(n_341),
.B(n_468),
.C(n_476),
.Y(n_946)
);

INVxp67_ASAP7_75t_SL g947 ( 
.A(n_726),
.Y(n_947)
);

BUFx8_ASAP7_75t_L g948 ( 
.A(n_792),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_742),
.B(n_522),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_689),
.A2(n_202),
.B1(n_336),
.B2(n_323),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_757),
.B(n_531),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_747),
.B(n_522),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_822),
.A2(n_571),
.B(n_618),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_687),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_767),
.B(n_531),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_783),
.B(n_192),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_783),
.B(n_198),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_822),
.A2(n_561),
.B(n_618),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_751),
.B(n_535),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_687),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_690),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_699),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_802),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_713),
.A2(n_561),
.B(n_618),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_749),
.B(n_650),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_749),
.B(n_650),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_713),
.A2(n_561),
.B(n_618),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_761),
.A2(n_724),
.B(n_720),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_805),
.Y(n_969)
);

AO21x1_ASAP7_75t_L g970 ( 
.A1(n_761),
.A2(n_478),
.B(n_480),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_731),
.A2(n_732),
.B(n_707),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_689),
.A2(n_557),
.B(n_612),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_783),
.B(n_198),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_714),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_797),
.A2(n_200),
.B1(n_337),
.B2(n_316),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_755),
.B(n_535),
.Y(n_976)
);

AOI21xp33_ASAP7_75t_L g977 ( 
.A1(n_798),
.A2(n_809),
.B(n_778),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_687),
.B(n_531),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_766),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_814),
.A2(n_557),
.B(n_612),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_814),
.A2(n_557),
.B(n_612),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_687),
.B(n_588),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_726),
.B(n_588),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_709),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_789),
.A2(n_580),
.B(n_612),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_771),
.B(n_535),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_800),
.A2(n_557),
.B(n_604),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_804),
.B(n_773),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_776),
.B(n_535),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_756),
.Y(n_990)
);

BUFx4f_ASAP7_75t_L g991 ( 
.A(n_735),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_809),
.A2(n_571),
.B(n_604),
.C(n_597),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_741),
.A2(n_571),
.B(n_604),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_793),
.A2(n_571),
.B(n_604),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_811),
.A2(n_816),
.B(n_812),
.Y(n_995)
);

NOR2xp67_ASAP7_75t_SL g996 ( 
.A(n_824),
.B(n_588),
.Y(n_996)
);

AND2x2_ASAP7_75t_SL g997 ( 
.A(n_782),
.B(n_807),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_819),
.A2(n_597),
.B(n_592),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_670),
.A2(n_677),
.B(n_700),
.C(n_825),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_807),
.A2(n_316),
.B1(n_200),
.B2(n_337),
.Y(n_1000)
);

AOI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_815),
.A2(n_611),
.B1(n_478),
.B2(n_597),
.Y(n_1001)
);

INVx2_ASAP7_75t_SL g1002 ( 
.A(n_795),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_772),
.B(n_580),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_735),
.Y(n_1004)
);

INVxp67_ASAP7_75t_L g1005 ( 
.A(n_753),
.Y(n_1005)
);

AO21x1_ASAP7_75t_L g1006 ( 
.A1(n_740),
.A2(n_478),
.B(n_480),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_752),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_824),
.B(n_345),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_768),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_823),
.A2(n_584),
.B(n_597),
.Y(n_1010)
);

O2A1O1Ixp5_ASAP7_75t_L g1011 ( 
.A1(n_740),
.A2(n_592),
.B(n_584),
.C(n_476),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_671),
.A2(n_584),
.B(n_592),
.Y(n_1012)
);

NOR3xp33_ASAP7_75t_L g1013 ( 
.A(n_759),
.B(n_188),
.C(n_194),
.Y(n_1013)
);

AOI21x1_ASAP7_75t_L g1014 ( 
.A1(n_680),
.A2(n_477),
.B(n_592),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_772),
.B(n_584),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_735),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_828),
.A2(n_611),
.B(n_588),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_735),
.B(n_179),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_911),
.B(n_726),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_892),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_988),
.B(n_907),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_977),
.B(n_726),
.Y(n_1022)
);

AOI221xp5_ASAP7_75t_L g1023 ( 
.A1(n_883),
.A2(n_317),
.B1(n_197),
.B2(n_188),
.C(n_321),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_SL g1024 ( 
.A1(n_1013),
.A2(n_727),
.B(n_683),
.C(n_738),
.Y(n_1024)
);

AOI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_942),
.A2(n_719),
.B1(n_726),
.B2(n_754),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_841),
.A2(n_785),
.B(n_719),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_837),
.A2(n_785),
.B(n_750),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_885),
.A2(n_818),
.B(n_750),
.C(n_760),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_939),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_867),
.B(n_726),
.Y(n_1030)
);

O2A1O1Ixp5_ASAP7_75t_L g1031 ( 
.A1(n_831),
.A2(n_827),
.B(n_794),
.C(n_784),
.Y(n_1031)
);

NAND2x1_ASAP7_75t_L g1032 ( 
.A(n_834),
.B(n_803),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_888),
.A2(n_315),
.B(n_252),
.C(n_256),
.Y(n_1033)
);

NOR2xp67_ASAP7_75t_L g1034 ( 
.A(n_832),
.B(n_250),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_939),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_848),
.Y(n_1036)
);

NAND3xp33_ASAP7_75t_L g1037 ( 
.A(n_1005),
.B(n_477),
.C(n_275),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_931),
.B(n_281),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_877),
.B(n_838),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_918),
.A2(n_956),
.B(n_973),
.C(n_957),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_928),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_850),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_939),
.Y(n_1043)
);

INVxp67_ASAP7_75t_SL g1044 ( 
.A(n_945),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_961),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_1018),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_913),
.A2(n_469),
.B(n_281),
.C(n_611),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_932),
.B(n_845),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_968),
.A2(n_588),
.B(n_552),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_947),
.A2(n_861),
.B1(n_901),
.B2(n_839),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_872),
.A2(n_539),
.B(n_803),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_925),
.A2(n_754),
.B1(n_611),
.B2(n_803),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_962),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_843),
.B(n_803),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_863),
.B(n_611),
.Y(n_1055)
);

INVx6_ASAP7_75t_SL g1056 ( 
.A(n_934),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_870),
.B(n_317),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_873),
.A2(n_880),
.B(n_842),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_897),
.B(n_272),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_849),
.B(n_321),
.Y(n_1060)
);

O2A1O1Ixp5_ASAP7_75t_L g1061 ( 
.A1(n_970),
.A2(n_469),
.B(n_276),
.C(n_311),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_945),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_904),
.B(n_324),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_940),
.A2(n_868),
.B(n_846),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_836),
.A2(n_539),
.B(n_469),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_851),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_836),
.A2(n_539),
.B(n_650),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_862),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_901),
.A2(n_306),
.B1(n_282),
.B2(n_285),
.Y(n_1069)
);

NAND2x1p5_ASAP7_75t_L g1070 ( 
.A(n_991),
.B(n_650),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_846),
.A2(n_833),
.B(n_1003),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_927),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_906),
.B(n_278),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_833),
.A2(n_539),
.B(n_294),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_919),
.A2(n_286),
.B(n_290),
.C(n_291),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_921),
.B(n_293),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_898),
.B(n_909),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_997),
.B(n_295),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1015),
.A2(n_296),
.B(n_470),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_974),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_933),
.B(n_326),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_855),
.A2(n_332),
.B(n_334),
.C(n_335),
.Y(n_1082)
);

OAI221xp5_ASAP7_75t_L g1083 ( 
.A1(n_894),
.A2(n_332),
.B1(n_334),
.B2(n_335),
.C(n_339),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_912),
.B(n_340),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_934),
.B(n_70),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_869),
.A2(n_470),
.B(n_437),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_R g1087 ( 
.A(n_1007),
.B(n_864),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_871),
.A2(n_470),
.B(n_437),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_900),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_945),
.B(n_340),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_954),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_SL g1092 ( 
.A(n_834),
.B(n_346),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_979),
.Y(n_1093)
);

INVx6_ASAP7_75t_L g1094 ( 
.A(n_948),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_834),
.A2(n_346),
.B1(n_343),
.B2(n_470),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_1009),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_954),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_1002),
.A2(n_343),
.B(n_10),
.C(n_11),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_R g1099 ( 
.A(n_864),
.B(n_68),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_938),
.B(n_8),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_876),
.A2(n_437),
.B1(n_71),
.B2(n_163),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_878),
.A2(n_470),
.B(n_437),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_989),
.A2(n_161),
.B(n_154),
.Y(n_1103)
);

CKINVDCx6p67_ASAP7_75t_R g1104 ( 
.A(n_929),
.Y(n_1104)
);

OR2x6_ASAP7_75t_SL g1105 ( 
.A(n_930),
.B(n_10),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_941),
.B(n_13),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_840),
.A2(n_153),
.B1(n_150),
.B2(n_145),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_853),
.A2(n_143),
.B1(n_133),
.B2(n_132),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_937),
.A2(n_128),
.B(n_126),
.Y(n_1109)
);

OAI21xp33_ASAP7_75t_SL g1110 ( 
.A1(n_844),
.A2(n_13),
.B(n_14),
.Y(n_1110)
);

NOR3xp33_ASAP7_75t_L g1111 ( 
.A(n_984),
.B(n_19),
.C(n_21),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_963),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_856),
.A2(n_119),
.B(n_110),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_1000),
.B(n_23),
.Y(n_1114)
);

NAND2x1p5_ASAP7_75t_L g1115 ( 
.A(n_991),
.B(n_105),
.Y(n_1115)
);

INVx1_ASAP7_75t_SL g1116 ( 
.A(n_1008),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_969),
.B(n_24),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_856),
.A2(n_85),
.B(n_81),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_972),
.A2(n_881),
.B(n_889),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_990),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_972),
.A2(n_76),
.B(n_72),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_834),
.A2(n_52),
.B1(n_25),
.B2(n_26),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_910),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_999),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_1124)
);

NAND2x1p5_ASAP7_75t_L g1125 ( 
.A(n_954),
.B(n_29),
.Y(n_1125)
);

O2A1O1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_895),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_965),
.B(n_33),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_971),
.A2(n_875),
.B(n_924),
.C(n_995),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_960),
.Y(n_1129)
);

OR2x6_ASAP7_75t_L g1130 ( 
.A(n_960),
.B(n_33),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_971),
.A2(n_34),
.B(n_36),
.C(n_42),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_995),
.A2(n_34),
.B(n_36),
.C(n_43),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_914),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_917),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_950),
.A2(n_43),
.B(n_48),
.C(n_51),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_960),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_886),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_890),
.A2(n_51),
.B(n_983),
.Y(n_1138)
);

AO22x1_ASAP7_75t_L g1139 ( 
.A1(n_834),
.A2(n_965),
.B1(n_966),
.B2(n_884),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_905),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_923),
.A2(n_891),
.B(n_992),
.C(n_975),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_920),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_854),
.B(n_866),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_966),
.Y(n_1144)
);

NAND2x1p5_ASAP7_75t_L g1145 ( 
.A(n_884),
.B(n_1016),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_943),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_944),
.Y(n_1147)
);

INVx1_ASAP7_75t_SL g1148 ( 
.A(n_1004),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_852),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_949),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_835),
.A2(n_922),
.B(n_993),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_R g1152 ( 
.A(n_1004),
.B(n_1016),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_857),
.A2(n_899),
.B(n_946),
.C(n_847),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_860),
.B(n_1006),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_952),
.Y(n_1155)
);

O2A1O1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_915),
.A2(n_959),
.B(n_986),
.C(n_976),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_865),
.A2(n_985),
.B(n_981),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_935),
.B(n_1001),
.Y(n_1158)
);

AOI221xp5_ASAP7_75t_L g1159 ( 
.A1(n_987),
.A2(n_951),
.B1(n_955),
.B2(n_980),
.C(n_981),
.Y(n_1159)
);

OR2x6_ASAP7_75t_L g1160 ( 
.A(n_980),
.B(n_987),
.Y(n_1160)
);

OAI21xp33_ASAP7_75t_L g1161 ( 
.A1(n_908),
.A2(n_887),
.B(n_953),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_865),
.A2(n_874),
.B(n_993),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_874),
.A2(n_1012),
.B(n_936),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_893),
.A2(n_1011),
.B(n_902),
.C(n_994),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_978),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_964),
.A2(n_967),
.B1(n_958),
.B2(n_1017),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_SL g1167 ( 
.A(n_996),
.B(n_967),
.Y(n_1167)
);

AOI21x1_ASAP7_75t_L g1168 ( 
.A1(n_858),
.A2(n_859),
.B(n_926),
.Y(n_1168)
);

INVx6_ASAP7_75t_L g1169 ( 
.A(n_982),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_859),
.B(n_1010),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_994),
.B(n_1010),
.Y(n_1171)
);

INVxp67_ASAP7_75t_L g1172 ( 
.A(n_926),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1119),
.A2(n_879),
.B(n_882),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1064),
.A2(n_879),
.B(n_882),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1116),
.B(n_998),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1036),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1040),
.B(n_998),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_SL g1178 ( 
.A1(n_1063),
.A2(n_896),
.B1(n_903),
.B2(n_916),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1060),
.A2(n_896),
.B(n_903),
.C(n_916),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1028),
.A2(n_1081),
.B(n_1141),
.C(n_1057),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_1166),
.A2(n_1128),
.A3(n_1162),
.B(n_1071),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1027),
.A2(n_1157),
.B(n_1058),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_1120),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1163),
.A2(n_1022),
.B(n_1026),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_1029),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1042),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_SL g1187 ( 
.A1(n_1131),
.A2(n_1024),
.B(n_1132),
.C(n_1082),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1123),
.B(n_1133),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1029),
.Y(n_1189)
);

BUFx8_ASAP7_75t_L g1190 ( 
.A(n_1072),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1172),
.A2(n_1138),
.B(n_1161),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1116),
.B(n_1020),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_SL g1193 ( 
.A1(n_1154),
.A2(n_1158),
.B(n_1033),
.C(n_1107),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1067),
.A2(n_1101),
.A3(n_1065),
.B(n_1049),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1114),
.A2(n_1153),
.B(n_1076),
.C(n_1037),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1127),
.Y(n_1196)
);

INVx6_ASAP7_75t_SL g1197 ( 
.A(n_1130),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1066),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1068),
.Y(n_1199)
);

AO22x2_ASAP7_75t_L g1200 ( 
.A1(n_1124),
.A2(n_1078),
.B1(n_1111),
.B2(n_1151),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1134),
.B(n_1039),
.Y(n_1201)
);

NAND3xp33_ASAP7_75t_L g1202 ( 
.A(n_1083),
.B(n_1038),
.C(n_1023),
.Y(n_1202)
);

O2A1O1Ixp5_ASAP7_75t_L g1203 ( 
.A1(n_1061),
.A2(n_1151),
.B(n_1171),
.C(n_1050),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1051),
.A2(n_1164),
.B(n_1156),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1031),
.A2(n_1170),
.B(n_1074),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1146),
.B(n_1147),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1037),
.A2(n_1161),
.B(n_1135),
.C(n_1121),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1159),
.A2(n_1025),
.B(n_1030),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_1129),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1167),
.A2(n_1019),
.B(n_1171),
.Y(n_1210)
);

O2A1O1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1126),
.A2(n_1098),
.B(n_1110),
.C(n_1090),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1167),
.A2(n_1160),
.B(n_1139),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1059),
.B(n_1073),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1113),
.A2(n_1118),
.B(n_1075),
.C(n_1155),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1089),
.Y(n_1215)
);

AO32x2_ASAP7_75t_L g1216 ( 
.A1(n_1108),
.A2(n_1069),
.A3(n_1160),
.B1(n_1035),
.B2(n_1097),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_1087),
.Y(n_1217)
);

O2A1O1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1100),
.A2(n_1106),
.B(n_1117),
.C(n_1084),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1029),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1055),
.A2(n_1150),
.B(n_1143),
.Y(n_1220)
);

OR2x6_ASAP7_75t_L g1221 ( 
.A(n_1094),
.B(n_1130),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1112),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1048),
.B(n_1144),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1086),
.A2(n_1102),
.A3(n_1088),
.B(n_1079),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1160),
.A2(n_1092),
.B(n_1032),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1077),
.B(n_1137),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1142),
.Y(n_1227)
);

CKINVDCx11_ASAP7_75t_R g1228 ( 
.A(n_1104),
.Y(n_1228)
);

CKINVDCx11_ASAP7_75t_R g1229 ( 
.A(n_1105),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1140),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1054),
.B(n_1080),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1041),
.B(n_1053),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1045),
.Y(n_1233)
);

INVx5_ASAP7_75t_L g1234 ( 
.A(n_1062),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1093),
.B(n_1096),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1145),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1092),
.A2(n_1103),
.B(n_1109),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1130),
.B(n_1125),
.Y(n_1238)
);

AO32x2_ASAP7_75t_L g1239 ( 
.A1(n_1035),
.A2(n_1097),
.A3(n_1122),
.B1(n_1034),
.B2(n_1047),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1062),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_1094),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1070),
.A2(n_1145),
.B(n_1115),
.Y(n_1242)
);

OR2x2_ASAP7_75t_L g1243 ( 
.A(n_1148),
.B(n_1043),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_1062),
.Y(n_1244)
);

AO31x2_ASAP7_75t_L g1245 ( 
.A1(n_1052),
.A2(n_1095),
.A3(n_1070),
.B(n_1115),
.Y(n_1245)
);

OAI22x1_ASAP7_75t_L g1246 ( 
.A1(n_1044),
.A2(n_1091),
.B1(n_1056),
.B2(n_1169),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1091),
.A2(n_1136),
.B(n_1165),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1165),
.Y(n_1248)
);

O2A1O1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1056),
.A2(n_1099),
.B(n_1169),
.C(n_1152),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1165),
.A2(n_556),
.B(n_977),
.C(n_762),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1136),
.B(n_1021),
.Y(n_1251)
);

O2A1O1Ixp33_ASAP7_75t_SL g1252 ( 
.A1(n_1136),
.A2(n_977),
.B(n_1028),
.C(n_1131),
.Y(n_1252)
);

NOR2xp67_ASAP7_75t_L g1253 ( 
.A(n_1037),
.B(n_718),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1036),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1040),
.B(n_348),
.Y(n_1255)
);

AO31x2_ASAP7_75t_L g1256 ( 
.A1(n_1166),
.A2(n_1128),
.A3(n_970),
.B(n_1162),
.Y(n_1256)
);

NAND3xp33_ASAP7_75t_SL g1257 ( 
.A(n_1040),
.B(n_556),
.C(n_1060),
.Y(n_1257)
);

NOR3xp33_ASAP7_75t_L g1258 ( 
.A(n_1040),
.B(n_546),
.C(n_526),
.Y(n_1258)
);

O2A1O1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1040),
.A2(n_1060),
.B(n_556),
.C(n_977),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1040),
.A2(n_556),
.B(n_977),
.C(n_762),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1168),
.A2(n_993),
.B(n_1162),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1036),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1119),
.A2(n_739),
.B(n_730),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1036),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1119),
.A2(n_739),
.B(n_730),
.Y(n_1265)
);

AO31x2_ASAP7_75t_L g1266 ( 
.A1(n_1166),
.A2(n_1128),
.A3(n_970),
.B(n_1162),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1119),
.A2(n_739),
.B(n_730),
.Y(n_1267)
);

INVx2_ASAP7_75t_SL g1268 ( 
.A(n_1020),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1040),
.B(n_348),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1168),
.A2(n_993),
.B(n_1162),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1149),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1119),
.A2(n_739),
.B(n_730),
.Y(n_1272)
);

AND2x6_ASAP7_75t_L g1273 ( 
.A(n_1085),
.B(n_1127),
.Y(n_1273)
);

INVx1_ASAP7_75t_SL g1274 ( 
.A(n_1020),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1119),
.A2(n_739),
.B(n_730),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1028),
.A2(n_977),
.B(n_675),
.Y(n_1276)
);

OAI22x1_ASAP7_75t_L g1277 ( 
.A1(n_1114),
.A2(n_762),
.B1(n_1060),
.B2(n_1007),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1120),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1028),
.A2(n_977),
.B(n_675),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1119),
.A2(n_739),
.B(n_730),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1168),
.A2(n_993),
.B(n_1162),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1020),
.Y(n_1282)
);

AOI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1060),
.A2(n_642),
.B1(n_546),
.B2(n_526),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1040),
.B(n_348),
.Y(n_1284)
);

A2O1A1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1040),
.A2(n_556),
.B(n_977),
.C(n_762),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_SL g1286 ( 
.A1(n_1028),
.A2(n_977),
.B(n_1131),
.C(n_1040),
.Y(n_1286)
);

A2O1A1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1040),
.A2(n_556),
.B(n_977),
.C(n_762),
.Y(n_1287)
);

AOI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1154),
.A2(n_1014),
.B(n_1027),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1166),
.A2(n_1128),
.A3(n_970),
.B(n_1162),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1021),
.B(n_675),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1119),
.A2(n_739),
.B(n_730),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1032),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1040),
.A2(n_556),
.B(n_977),
.C(n_762),
.Y(n_1293)
);

INVxp67_ASAP7_75t_L g1294 ( 
.A(n_1020),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1048),
.B(n_1046),
.Y(n_1295)
);

OA21x2_ASAP7_75t_L g1296 ( 
.A1(n_1151),
.A2(n_1071),
.B(n_1064),
.Y(n_1296)
);

AO31x2_ASAP7_75t_L g1297 ( 
.A1(n_1166),
.A2(n_1128),
.A3(n_970),
.B(n_1162),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1021),
.A2(n_556),
.B1(n_911),
.B2(n_977),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1036),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1021),
.A2(n_556),
.B1(n_911),
.B2(n_977),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1119),
.A2(n_739),
.B(n_730),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1028),
.A2(n_977),
.B(n_675),
.Y(n_1302)
);

AO21x1_ASAP7_75t_L g1303 ( 
.A1(n_1154),
.A2(n_977),
.B(n_556),
.Y(n_1303)
);

O2A1O1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1040),
.A2(n_1060),
.B(n_556),
.C(n_977),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1021),
.B(n_675),
.Y(n_1305)
);

OAI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1116),
.A2(n_517),
.B1(n_619),
.B2(n_590),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1036),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1119),
.A2(n_739),
.B(n_730),
.Y(n_1308)
);

AO32x2_ASAP7_75t_L g1309 ( 
.A1(n_1166),
.A2(n_1124),
.A3(n_1002),
.B1(n_895),
.B2(n_891),
.Y(n_1309)
);

O2A1O1Ixp33_ASAP7_75t_L g1310 ( 
.A1(n_1040),
.A2(n_1060),
.B(n_556),
.C(n_977),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1036),
.Y(n_1311)
);

BUFx4_ASAP7_75t_SL g1312 ( 
.A(n_1089),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_1089),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1168),
.A2(n_993),
.B(n_1162),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1119),
.A2(n_739),
.B(n_730),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1028),
.A2(n_977),
.B(n_675),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1021),
.B(n_675),
.Y(n_1317)
);

CKINVDCx16_ASAP7_75t_R g1318 ( 
.A(n_1089),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_1020),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1168),
.A2(n_993),
.B(n_1162),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1168),
.A2(n_993),
.B(n_1162),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1028),
.A2(n_977),
.B(n_675),
.Y(n_1322)
);

AOI31xp67_ASAP7_75t_L g1323 ( 
.A1(n_1154),
.A2(n_1171),
.A3(n_706),
.B(n_704),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1119),
.A2(n_739),
.B(n_730),
.Y(n_1324)
);

AO31x2_ASAP7_75t_L g1325 ( 
.A1(n_1166),
.A2(n_1128),
.A3(n_970),
.B(n_1162),
.Y(n_1325)
);

BUFx4f_ASAP7_75t_SL g1326 ( 
.A(n_1197),
.Y(n_1326)
);

INVx4_ASAP7_75t_L g1327 ( 
.A(n_1234),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1258),
.A2(n_1257),
.B1(n_1283),
.B2(n_1255),
.Y(n_1328)
);

BUFx2_ASAP7_75t_SL g1329 ( 
.A(n_1183),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1181),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_1313),
.Y(n_1331)
);

CKINVDCx14_ASAP7_75t_R g1332 ( 
.A(n_1228),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_SL g1333 ( 
.A1(n_1269),
.A2(n_1284),
.B1(n_1276),
.B2(n_1322),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1312),
.Y(n_1334)
);

INVx6_ASAP7_75t_L g1335 ( 
.A(n_1234),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_SL g1336 ( 
.A1(n_1279),
.A2(n_1302),
.B1(n_1316),
.B2(n_1202),
.Y(n_1336)
);

BUFx8_ASAP7_75t_L g1337 ( 
.A(n_1282),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1176),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_SL g1339 ( 
.A1(n_1259),
.A2(n_1310),
.B(n_1304),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1290),
.B(n_1305),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1222),
.Y(n_1341)
);

OAI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1317),
.A2(n_1277),
.B1(n_1221),
.B2(n_1188),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1180),
.A2(n_1260),
.B1(n_1293),
.B2(n_1285),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1234),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1262),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_SL g1346 ( 
.A1(n_1200),
.A2(n_1273),
.B1(n_1298),
.B2(n_1300),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_SL g1347 ( 
.A1(n_1200),
.A2(n_1273),
.B1(n_1221),
.B2(n_1238),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1274),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_SL g1349 ( 
.A1(n_1273),
.A2(n_1213),
.B1(n_1212),
.B2(n_1229),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1253),
.A2(n_1273),
.B1(n_1287),
.B2(n_1306),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1185),
.Y(n_1351)
);

INVx6_ASAP7_75t_L g1352 ( 
.A(n_1190),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1303),
.A2(n_1191),
.B1(n_1175),
.B2(n_1201),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1195),
.A2(n_1250),
.B1(n_1206),
.B2(n_1196),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1197),
.A2(n_1177),
.B1(n_1299),
.B2(n_1226),
.Y(n_1355)
);

OAI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1251),
.A2(n_1264),
.B1(n_1198),
.B2(n_1186),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1199),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1319),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1218),
.B(n_1192),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1295),
.B(n_1232),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1210),
.A2(n_1208),
.B1(n_1190),
.B2(n_1307),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_1268),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1254),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1227),
.A2(n_1178),
.B1(n_1233),
.B2(n_1230),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1295),
.A2(n_1235),
.B1(n_1223),
.B2(n_1220),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1311),
.Y(n_1366)
);

AOI21xp33_ASAP7_75t_L g1367 ( 
.A1(n_1211),
.A2(n_1207),
.B(n_1203),
.Y(n_1367)
);

BUFx10_ASAP7_75t_L g1368 ( 
.A(n_1215),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_1318),
.Y(n_1369)
);

INVx2_ASAP7_75t_SL g1370 ( 
.A(n_1278),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1294),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_1217),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_1241),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1223),
.B(n_1235),
.Y(n_1374)
);

INVx1_ASAP7_75t_SL g1375 ( 
.A(n_1209),
.Y(n_1375)
);

INVx1_ASAP7_75t_SL g1376 ( 
.A(n_1243),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1271),
.Y(n_1377)
);

INVx6_ASAP7_75t_L g1378 ( 
.A(n_1189),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1248),
.Y(n_1379)
);

INVx1_ASAP7_75t_SL g1380 ( 
.A(n_1248),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1231),
.Y(n_1381)
);

INVx4_ASAP7_75t_L g1382 ( 
.A(n_1189),
.Y(n_1382)
);

BUFx2_ASAP7_75t_SL g1383 ( 
.A(n_1219),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_SL g1384 ( 
.A(n_1219),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1246),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1219),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_SL g1387 ( 
.A1(n_1225),
.A2(n_1247),
.B1(n_1236),
.B2(n_1244),
.Y(n_1387)
);

CKINVDCx11_ASAP7_75t_R g1388 ( 
.A(n_1240),
.Y(n_1388)
);

CKINVDCx11_ASAP7_75t_R g1389 ( 
.A(n_1240),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1214),
.A2(n_1286),
.B(n_1237),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1249),
.A2(n_1292),
.B1(n_1324),
.B2(n_1291),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1296),
.A2(n_1182),
.B1(n_1204),
.B2(n_1292),
.Y(n_1392)
);

BUFx8_ASAP7_75t_L g1393 ( 
.A(n_1240),
.Y(n_1393)
);

BUFx8_ASAP7_75t_SL g1394 ( 
.A(n_1288),
.Y(n_1394)
);

INVx4_ASAP7_75t_L g1395 ( 
.A(n_1296),
.Y(n_1395)
);

BUFx4f_ASAP7_75t_SL g1396 ( 
.A(n_1252),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1263),
.A2(n_1265),
.B1(n_1315),
.B2(n_1267),
.Y(n_1397)
);

CKINVDCx14_ASAP7_75t_R g1398 ( 
.A(n_1187),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1323),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1242),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1193),
.B(n_1266),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_1184),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_SL g1403 ( 
.A1(n_1309),
.A2(n_1275),
.B1(n_1272),
.B2(n_1280),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1173),
.A2(n_1309),
.B1(n_1321),
.B2(n_1320),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1239),
.B(n_1309),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_SL g1406 ( 
.A1(n_1301),
.A2(n_1308),
.B1(n_1239),
.B2(n_1314),
.Y(n_1406)
);

INVx4_ASAP7_75t_L g1407 ( 
.A(n_1216),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_1174),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1179),
.A2(n_1216),
.B1(n_1239),
.B2(n_1245),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1256),
.Y(n_1410)
);

BUFx2_ASAP7_75t_SL g1411 ( 
.A(n_1216),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1261),
.A2(n_1281),
.B1(n_1270),
.B2(n_1205),
.Y(n_1412)
);

BUFx12f_ASAP7_75t_L g1413 ( 
.A(n_1245),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1266),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1245),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1325),
.A2(n_1289),
.B1(n_1297),
.B2(n_1194),
.Y(n_1416)
);

OAI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1289),
.A2(n_1297),
.B1(n_1325),
.B2(n_1194),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1194),
.A2(n_1224),
.B1(n_1283),
.B2(n_1040),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1224),
.A2(n_1258),
.B1(n_1257),
.B2(n_556),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1312),
.Y(n_1420)
);

CKINVDCx11_ASAP7_75t_R g1421 ( 
.A(n_1228),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_SL g1422 ( 
.A1(n_1255),
.A2(n_1269),
.B1(n_1284),
.B2(n_556),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1282),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1258),
.A2(n_1257),
.B1(n_556),
.B2(n_1283),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1181),
.Y(n_1425)
);

CKINVDCx11_ASAP7_75t_R g1426 ( 
.A(n_1228),
.Y(n_1426)
);

BUFx8_ASAP7_75t_L g1427 ( 
.A(n_1282),
.Y(n_1427)
);

OAI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1283),
.A2(n_1105),
.B1(n_1130),
.B2(n_1202),
.Y(n_1428)
);

BUFx4f_ASAP7_75t_SL g1429 ( 
.A(n_1197),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_1313),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1258),
.A2(n_1257),
.B1(n_556),
.B2(n_1283),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1282),
.Y(n_1432)
);

INVx6_ASAP7_75t_L g1433 ( 
.A(n_1234),
.Y(n_1433)
);

NAND2x1p5_ASAP7_75t_L g1434 ( 
.A(n_1234),
.B(n_1242),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1222),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1312),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1276),
.A2(n_1302),
.B(n_1279),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1258),
.A2(n_1257),
.B1(n_556),
.B2(n_1283),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1185),
.Y(n_1439)
);

INVx6_ASAP7_75t_L g1440 ( 
.A(n_1234),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_SL g1441 ( 
.A1(n_1255),
.A2(n_1269),
.B1(n_1284),
.B2(n_556),
.Y(n_1441)
);

INVx6_ASAP7_75t_L g1442 ( 
.A(n_1234),
.Y(n_1442)
);

BUFx2_ASAP7_75t_L g1443 ( 
.A(n_1282),
.Y(n_1443)
);

INVx4_ASAP7_75t_L g1444 ( 
.A(n_1234),
.Y(n_1444)
);

NAND2x1p5_ASAP7_75t_L g1445 ( 
.A(n_1234),
.B(n_1242),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_SL g1446 ( 
.A1(n_1255),
.A2(n_1269),
.B1(n_1284),
.B2(n_556),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1283),
.A2(n_1040),
.B1(n_1180),
.B2(n_556),
.Y(n_1447)
);

CKINVDCx20_ASAP7_75t_R g1448 ( 
.A(n_1313),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1258),
.A2(n_1257),
.B1(n_556),
.B2(n_1283),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1410),
.Y(n_1450)
);

INVx2_ASAP7_75t_SL g1451 ( 
.A(n_1335),
.Y(n_1451)
);

OR2x6_ASAP7_75t_L g1452 ( 
.A(n_1437),
.B(n_1413),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1414),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1330),
.Y(n_1454)
);

OAI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1333),
.A2(n_1447),
.B(n_1336),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1376),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1422),
.A2(n_1446),
.B1(n_1441),
.B2(n_1333),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1330),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1407),
.B(n_1405),
.Y(n_1459)
);

BUFx10_ASAP7_75t_L g1460 ( 
.A(n_1352),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1380),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1400),
.B(n_1408),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1422),
.A2(n_1446),
.B1(n_1441),
.B2(n_1328),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1399),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1395),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1394),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1395),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1425),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_SL g1469 ( 
.A(n_1334),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1407),
.B(n_1409),
.Y(n_1470)
);

OAI222xp33_ASAP7_75t_L g1471 ( 
.A1(n_1328),
.A2(n_1336),
.B1(n_1428),
.B2(n_1438),
.C1(n_1431),
.C2(n_1424),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1411),
.B(n_1353),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1397),
.A2(n_1390),
.B(n_1412),
.Y(n_1473)
);

BUFx12f_ASAP7_75t_L g1474 ( 
.A(n_1421),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1341),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1375),
.Y(n_1476)
);

AO21x2_ASAP7_75t_L g1477 ( 
.A1(n_1367),
.A2(n_1417),
.B(n_1401),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1353),
.B(n_1419),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1381),
.B(n_1340),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1419),
.B(n_1435),
.Y(n_1480)
);

INVx4_ASAP7_75t_L g1481 ( 
.A(n_1344),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1418),
.B(n_1415),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1402),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1331),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1398),
.A2(n_1428),
.B1(n_1424),
.B2(n_1449),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1377),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1357),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1363),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1366),
.Y(n_1489)
);

AND2x2_ASAP7_75t_SL g1490 ( 
.A(n_1431),
.B(n_1449),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1434),
.Y(n_1491)
);

AOI21xp33_ASAP7_75t_L g1492 ( 
.A1(n_1438),
.A2(n_1339),
.B(n_1343),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1417),
.Y(n_1493)
);

OAI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1354),
.A2(n_1364),
.B(n_1359),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1416),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1445),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1416),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1412),
.A2(n_1392),
.B(n_1404),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1356),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1379),
.B(n_1346),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1360),
.B(n_1423),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1356),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1345),
.Y(n_1503)
);

BUFx4f_ASAP7_75t_SL g1504 ( 
.A(n_1448),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1432),
.Y(n_1505)
);

OA21x2_ASAP7_75t_L g1506 ( 
.A1(n_1404),
.A2(n_1392),
.B(n_1364),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1346),
.B(n_1347),
.Y(n_1507)
);

INVxp67_ASAP7_75t_SL g1508 ( 
.A(n_1338),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1391),
.A2(n_1355),
.B(n_1350),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1443),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1396),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1396),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1347),
.B(n_1361),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1327),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1403),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1337),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1387),
.B(n_1355),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1361),
.A2(n_1342),
.B(n_1403),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1406),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1406),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1342),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1337),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1348),
.B(n_1358),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1365),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1349),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1349),
.A2(n_1385),
.B1(n_1374),
.B2(n_1352),
.Y(n_1526)
);

INVx6_ASAP7_75t_L g1527 ( 
.A(n_1393),
.Y(n_1527)
);

INVx8_ASAP7_75t_L g1528 ( 
.A(n_1344),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1327),
.B(n_1444),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1335),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1335),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1352),
.A2(n_1371),
.B1(n_1369),
.B2(n_1362),
.Y(n_1532)
);

A2O1A1Ixp33_ASAP7_75t_L g1533 ( 
.A1(n_1455),
.A2(n_1372),
.B(n_1386),
.C(n_1439),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1471),
.B(n_1427),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1499),
.B(n_1386),
.Y(n_1535)
);

OA21x2_ASAP7_75t_L g1536 ( 
.A1(n_1498),
.A2(n_1370),
.B(n_1384),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1459),
.B(n_1329),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_SL g1538 ( 
.A1(n_1466),
.A2(n_1430),
.B1(n_1332),
.B2(n_1420),
.Y(n_1538)
);

OR2x6_ASAP7_75t_L g1539 ( 
.A(n_1452),
.B(n_1442),
.Y(n_1539)
);

OAI21xp33_ASAP7_75t_L g1540 ( 
.A1(n_1463),
.A2(n_1436),
.B(n_1373),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1505),
.Y(n_1541)
);

AND2x4_ASAP7_75t_SL g1542 ( 
.A(n_1484),
.B(n_1368),
.Y(n_1542)
);

OAI21xp33_ASAP7_75t_L g1543 ( 
.A1(n_1457),
.A2(n_1351),
.B(n_1326),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1475),
.Y(n_1544)
);

AOI221xp5_ASAP7_75t_L g1545 ( 
.A1(n_1455),
.A2(n_1382),
.B1(n_1351),
.B2(n_1383),
.C(n_1429),
.Y(n_1545)
);

CKINVDCx14_ASAP7_75t_R g1546 ( 
.A(n_1474),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1462),
.B(n_1368),
.Y(n_1547)
);

AO32x2_ASAP7_75t_L g1548 ( 
.A1(n_1485),
.A2(n_1388),
.A3(n_1389),
.B1(n_1378),
.B2(n_1326),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1499),
.B(n_1433),
.Y(n_1549)
);

AO32x2_ASAP7_75t_L g1550 ( 
.A1(n_1470),
.A2(n_1378),
.A3(n_1429),
.B1(n_1433),
.B2(n_1440),
.Y(n_1550)
);

OAI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1494),
.A2(n_1433),
.B(n_1440),
.Y(n_1551)
);

AOI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1490),
.A2(n_1426),
.B1(n_1442),
.B2(n_1494),
.Y(n_1552)
);

AOI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1490),
.A2(n_1492),
.B1(n_1526),
.B2(n_1525),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1454),
.Y(n_1554)
);

OAI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1492),
.A2(n_1490),
.B(n_1509),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1460),
.Y(n_1556)
);

O2A1O1Ixp33_ASAP7_75t_SL g1557 ( 
.A1(n_1518),
.A2(n_1526),
.B(n_1512),
.C(n_1511),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1521),
.B(n_1500),
.Y(n_1558)
);

BUFx2_ASAP7_75t_L g1559 ( 
.A(n_1505),
.Y(n_1559)
);

CKINVDCx6p67_ASAP7_75t_R g1560 ( 
.A(n_1474),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1521),
.B(n_1500),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1507),
.A2(n_1479),
.B1(n_1466),
.B2(n_1512),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1469),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1483),
.B(n_1501),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1456),
.B(n_1487),
.Y(n_1565)
);

O2A1O1Ixp5_ASAP7_75t_L g1566 ( 
.A1(n_1518),
.A2(n_1515),
.B(n_1520),
.C(n_1519),
.Y(n_1566)
);

CKINVDCx20_ASAP7_75t_R g1567 ( 
.A(n_1504),
.Y(n_1567)
);

AO32x2_ASAP7_75t_L g1568 ( 
.A1(n_1451),
.A2(n_1481),
.A3(n_1495),
.B1(n_1497),
.B2(n_1515),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1487),
.B(n_1488),
.Y(n_1569)
);

OA21x2_ASAP7_75t_L g1570 ( 
.A1(n_1498),
.A2(n_1473),
.B(n_1509),
.Y(n_1570)
);

AO32x2_ASAP7_75t_L g1571 ( 
.A1(n_1481),
.A2(n_1493),
.A3(n_1480),
.B1(n_1520),
.B2(n_1519),
.Y(n_1571)
);

AO21x1_ASAP7_75t_L g1572 ( 
.A1(n_1507),
.A2(n_1517),
.B(n_1525),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1502),
.B(n_1480),
.Y(n_1573)
);

AOI22x1_ASAP7_75t_L g1574 ( 
.A1(n_1512),
.A2(n_1511),
.B1(n_1483),
.B2(n_1513),
.Y(n_1574)
);

OAI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1478),
.A2(n_1473),
.B(n_1517),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_SL g1576 ( 
.A(n_1466),
.B(n_1474),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1472),
.B(n_1513),
.Y(n_1577)
);

OA21x2_ASAP7_75t_L g1578 ( 
.A1(n_1464),
.A2(n_1493),
.B(n_1453),
.Y(n_1578)
);

NOR2x1_ASAP7_75t_L g1579 ( 
.A(n_1496),
.B(n_1530),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1472),
.B(n_1486),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1486),
.B(n_1510),
.Y(n_1581)
);

OAI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1478),
.A2(n_1517),
.B(n_1524),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1461),
.B(n_1488),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_SL g1584 ( 
.A1(n_1517),
.A2(n_1524),
.B1(n_1477),
.B2(n_1506),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1477),
.A2(n_1452),
.B(n_1506),
.Y(n_1585)
);

AOI221xp5_ASAP7_75t_L g1586 ( 
.A1(n_1476),
.A2(n_1523),
.B1(n_1482),
.B2(n_1477),
.C(n_1503),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_SL g1587 ( 
.A1(n_1527),
.A2(n_1532),
.B1(n_1516),
.B2(n_1522),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1578),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1578),
.Y(n_1589)
);

INVxp67_ASAP7_75t_SL g1590 ( 
.A(n_1554),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1544),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1570),
.B(n_1477),
.Y(n_1592)
);

OR2x2_ASAP7_75t_SL g1593 ( 
.A(n_1536),
.B(n_1527),
.Y(n_1593)
);

NAND3xp33_ASAP7_75t_L g1594 ( 
.A(n_1586),
.B(n_1482),
.C(n_1532),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1554),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1562),
.B(n_1452),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1534),
.A2(n_1512),
.B1(n_1506),
.B2(n_1511),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1575),
.B(n_1467),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1573),
.B(n_1583),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1569),
.Y(n_1600)
);

BUFx3_ASAP7_75t_L g1601 ( 
.A(n_1536),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1553),
.A2(n_1527),
.B1(n_1516),
.B2(n_1522),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1585),
.B(n_1468),
.Y(n_1603)
);

NOR2x1_ASAP7_75t_L g1604 ( 
.A(n_1539),
.B(n_1491),
.Y(n_1604)
);

NOR2xp67_ASAP7_75t_L g1605 ( 
.A(n_1585),
.B(n_1491),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1573),
.B(n_1468),
.Y(n_1606)
);

OAI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1555),
.A2(n_1506),
.B(n_1508),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1571),
.Y(n_1608)
);

BUFx2_ASAP7_75t_L g1609 ( 
.A(n_1550),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1571),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1562),
.B(n_1531),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1565),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1586),
.B(n_1489),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1571),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1580),
.B(n_1458),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1571),
.B(n_1465),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1595),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1609),
.B(n_1584),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1589),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1599),
.B(n_1576),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1589),
.Y(n_1621)
);

NAND4xp25_ASAP7_75t_L g1622 ( 
.A(n_1594),
.B(n_1534),
.C(n_1566),
.D(n_1552),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1589),
.Y(n_1623)
);

AO21x2_ASAP7_75t_L g1624 ( 
.A1(n_1592),
.A2(n_1555),
.B(n_1450),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1609),
.B(n_1584),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1615),
.B(n_1541),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_1589),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1595),
.Y(n_1628)
);

INVx1_ASAP7_75t_SL g1629 ( 
.A(n_1612),
.Y(n_1629)
);

NOR3xp33_ASAP7_75t_L g1630 ( 
.A(n_1594),
.B(n_1540),
.C(n_1557),
.Y(n_1630)
);

AOI221xp5_ASAP7_75t_L g1631 ( 
.A1(n_1594),
.A2(n_1557),
.B1(n_1566),
.B2(n_1582),
.C(n_1572),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1615),
.B(n_1559),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1590),
.Y(n_1633)
);

INVx4_ASAP7_75t_L g1634 ( 
.A(n_1601),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1609),
.B(n_1568),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1590),
.Y(n_1636)
);

NAND4xp25_ASAP7_75t_SL g1637 ( 
.A(n_1597),
.B(n_1533),
.C(n_1545),
.D(n_1582),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1615),
.B(n_1581),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1616),
.B(n_1568),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1599),
.B(n_1576),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1612),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1606),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1589),
.Y(n_1643)
);

OAI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1597),
.A2(n_1543),
.B1(n_1533),
.B2(n_1551),
.C(n_1574),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1591),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1589),
.Y(n_1646)
);

AOI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1613),
.A2(n_1587),
.B1(n_1551),
.B2(n_1577),
.C(n_1558),
.Y(n_1647)
);

NAND3xp33_ASAP7_75t_SL g1648 ( 
.A(n_1602),
.B(n_1545),
.C(n_1563),
.Y(n_1648)
);

OAI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1607),
.A2(n_1549),
.B(n_1579),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1616),
.B(n_1568),
.Y(n_1650)
);

NAND4xp25_ASAP7_75t_L g1651 ( 
.A(n_1607),
.B(n_1549),
.C(n_1538),
.D(n_1535),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1588),
.Y(n_1652)
);

AOI31xp33_ASAP7_75t_SL g1653 ( 
.A1(n_1596),
.A2(n_1537),
.A3(n_1548),
.B(n_1546),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1616),
.B(n_1568),
.Y(n_1654)
);

OAI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1602),
.A2(n_1539),
.B(n_1535),
.Y(n_1655)
);

INVxp67_ASAP7_75t_SL g1656 ( 
.A(n_1588),
.Y(n_1656)
);

INVxp67_ASAP7_75t_SL g1657 ( 
.A(n_1588),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1591),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1588),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_1628),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1639),
.B(n_1608),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1645),
.Y(n_1662)
);

NAND2x1p5_ASAP7_75t_L g1663 ( 
.A(n_1634),
.B(n_1604),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1629),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1645),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1650),
.B(n_1598),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1659),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1650),
.B(n_1598),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1654),
.B(n_1610),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1654),
.B(n_1610),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1654),
.B(n_1635),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1658),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1635),
.B(n_1614),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1629),
.B(n_1606),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1659),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1659),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1620),
.B(n_1560),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1618),
.B(n_1598),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_1641),
.Y(n_1679)
);

NAND4xp25_ASAP7_75t_L g1680 ( 
.A(n_1631),
.B(n_1613),
.C(n_1596),
.D(n_1592),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1658),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_R g1682 ( 
.A(n_1648),
.B(n_1567),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1635),
.B(n_1614),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1642),
.B(n_1606),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1618),
.B(n_1606),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1643),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1633),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1633),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1652),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1636),
.B(n_1614),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1636),
.B(n_1600),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1634),
.B(n_1601),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1617),
.B(n_1600),
.Y(n_1693)
);

NAND2x1p5_ASAP7_75t_L g1694 ( 
.A(n_1634),
.B(n_1604),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1617),
.B(n_1600),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1677),
.B(n_1516),
.Y(n_1696)
);

BUFx2_ASAP7_75t_L g1697 ( 
.A(n_1663),
.Y(n_1697)
);

OAI33xp33_ASAP7_75t_L g1698 ( 
.A1(n_1680),
.A2(n_1651),
.A3(n_1622),
.B1(n_1603),
.B2(n_1626),
.B3(n_1632),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1678),
.B(n_1618),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1662),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1692),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1662),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1686),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1680),
.B(n_1631),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1679),
.B(n_1640),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1678),
.B(n_1625),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1679),
.B(n_1647),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1665),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1664),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1665),
.Y(n_1710)
);

OAI21xp33_ASAP7_75t_L g1711 ( 
.A1(n_1682),
.A2(n_1622),
.B(n_1630),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1671),
.B(n_1625),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1686),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1671),
.B(n_1666),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1686),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1664),
.B(n_1522),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1685),
.B(n_1625),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1672),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1685),
.B(n_1647),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1672),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1692),
.B(n_1671),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1666),
.B(n_1634),
.Y(n_1722)
);

INVxp67_ASAP7_75t_L g1723 ( 
.A(n_1693),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1681),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1674),
.B(n_1651),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1681),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1689),
.Y(n_1727)
);

NOR2x1_ASAP7_75t_L g1728 ( 
.A(n_1692),
.B(n_1648),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_R g1729 ( 
.A(n_1687),
.B(n_1527),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1687),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1688),
.Y(n_1731)
);

BUFx3_ASAP7_75t_L g1732 ( 
.A(n_1692),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1692),
.B(n_1601),
.Y(n_1733)
);

INVxp67_ASAP7_75t_SL g1734 ( 
.A(n_1663),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1674),
.B(n_1564),
.Y(n_1735)
);

AOI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1663),
.A2(n_1630),
.B1(n_1637),
.B2(n_1644),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1693),
.B(n_1638),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1695),
.B(n_1638),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1700),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1717),
.B(n_1660),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1700),
.Y(n_1741)
);

INVx2_ASAP7_75t_SL g1742 ( 
.A(n_1721),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1702),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1712),
.B(n_1668),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1712),
.B(n_1668),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1699),
.B(n_1673),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1704),
.B(n_1660),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1702),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1708),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1711),
.B(n_1649),
.Y(n_1750)
);

AOI211xp5_ASAP7_75t_L g1751 ( 
.A1(n_1736),
.A2(n_1653),
.B(n_1637),
.C(n_1644),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1708),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1709),
.B(n_1649),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1710),
.Y(n_1754)
);

AOI21xp33_ASAP7_75t_L g1755 ( 
.A1(n_1728),
.A2(n_1655),
.B(n_1624),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1714),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1710),
.Y(n_1757)
);

AOI211x1_ASAP7_75t_SL g1758 ( 
.A1(n_1707),
.A2(n_1655),
.B(n_1690),
.C(n_1689),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1699),
.B(n_1673),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1717),
.B(n_1690),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1709),
.B(n_1688),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1719),
.B(n_1695),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1737),
.B(n_1691),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1738),
.B(n_1691),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1706),
.B(n_1684),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1718),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1725),
.B(n_1684),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1718),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_1729),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1705),
.B(n_1561),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1720),
.Y(n_1771)
);

INVxp67_ASAP7_75t_SL g1772 ( 
.A(n_1728),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1706),
.B(n_1624),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1720),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1767),
.B(n_1735),
.Y(n_1775)
);

NAND2xp33_ASAP7_75t_SL g1776 ( 
.A(n_1750),
.B(n_1697),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1742),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1772),
.B(n_1698),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1751),
.B(n_1716),
.Y(n_1779)
);

AOI31xp33_ASAP7_75t_L g1780 ( 
.A1(n_1769),
.A2(n_1696),
.A3(n_1694),
.B(n_1663),
.Y(n_1780)
);

AOI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1747),
.A2(n_1721),
.B1(n_1722),
.B2(n_1701),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1758),
.B(n_1721),
.Y(n_1782)
);

XNOR2x1_ASAP7_75t_L g1783 ( 
.A(n_1753),
.B(n_1547),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1739),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1742),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1741),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1762),
.A2(n_1756),
.B1(n_1755),
.B2(n_1770),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1746),
.B(n_1759),
.Y(n_1788)
);

OAI211xp5_ASAP7_75t_L g1789 ( 
.A1(n_1761),
.A2(n_1734),
.B(n_1697),
.C(n_1701),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1743),
.Y(n_1790)
);

OAI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1756),
.A2(n_1714),
.B1(n_1694),
.B2(n_1593),
.Y(n_1791)
);

INVxp67_ASAP7_75t_SL g1792 ( 
.A(n_1740),
.Y(n_1792)
);

OAI221xp5_ASAP7_75t_SL g1793 ( 
.A1(n_1740),
.A2(n_1723),
.B1(n_1732),
.B2(n_1722),
.C(n_1713),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1748),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1749),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1744),
.B(n_1732),
.Y(n_1796)
);

OAI322xp33_ASAP7_75t_L g1797 ( 
.A1(n_1765),
.A2(n_1773),
.A3(n_1760),
.B1(n_1771),
.B2(n_1768),
.C1(n_1766),
.C2(n_1752),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1744),
.B(n_1703),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1754),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1757),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1792),
.B(n_1765),
.Y(n_1801)
);

OAI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1778),
.A2(n_1694),
.B(n_1774),
.Y(n_1802)
);

INVx1_ASAP7_75t_SL g1803 ( 
.A(n_1776),
.Y(n_1803)
);

OAI311xp33_ASAP7_75t_L g1804 ( 
.A1(n_1779),
.A2(n_1760),
.A3(n_1773),
.B1(n_1763),
.C1(n_1764),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1777),
.Y(n_1805)
);

XNOR2xp5_ASAP7_75t_L g1806 ( 
.A(n_1783),
.B(n_1542),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1778),
.A2(n_1776),
.B1(n_1782),
.B2(n_1783),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1788),
.B(n_1746),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1775),
.B(n_1763),
.Y(n_1809)
);

AND2x4_ASAP7_75t_L g1810 ( 
.A(n_1777),
.B(n_1759),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1793),
.B(n_1764),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1785),
.Y(n_1812)
);

INVx1_ASAP7_75t_SL g1813 ( 
.A(n_1785),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1796),
.Y(n_1814)
);

OAI21xp33_ASAP7_75t_L g1815 ( 
.A1(n_1781),
.A2(n_1789),
.B(n_1798),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1784),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1787),
.B(n_1703),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1786),
.Y(n_1818)
);

INVx1_ASAP7_75t_SL g1819 ( 
.A(n_1788),
.Y(n_1819)
);

INVx2_ASAP7_75t_SL g1820 ( 
.A(n_1790),
.Y(n_1820)
);

INVxp67_ASAP7_75t_SL g1821 ( 
.A(n_1794),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1819),
.B(n_1745),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1810),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1808),
.B(n_1745),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1801),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1805),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1814),
.B(n_1795),
.Y(n_1827)
);

NOR3xp33_ASAP7_75t_L g1828 ( 
.A(n_1803),
.B(n_1797),
.C(n_1780),
.Y(n_1828)
);

NOR2x1_ASAP7_75t_L g1829 ( 
.A(n_1812),
.B(n_1799),
.Y(n_1829)
);

INVx1_ASAP7_75t_SL g1830 ( 
.A(n_1813),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1807),
.B(n_1800),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1806),
.B(n_1791),
.Y(n_1832)
);

NAND3xp33_ASAP7_75t_L g1833 ( 
.A(n_1807),
.B(n_1715),
.C(n_1713),
.Y(n_1833)
);

AOI221xp5_ASAP7_75t_L g1834 ( 
.A1(n_1828),
.A2(n_1804),
.B1(n_1811),
.B2(n_1815),
.C(n_1817),
.Y(n_1834)
);

NAND4xp75_ASAP7_75t_L g1835 ( 
.A(n_1831),
.B(n_1817),
.C(n_1811),
.D(n_1802),
.Y(n_1835)
);

NAND3xp33_ASAP7_75t_L g1836 ( 
.A(n_1831),
.B(n_1821),
.C(n_1818),
.Y(n_1836)
);

NAND3xp33_ASAP7_75t_SL g1837 ( 
.A(n_1830),
.B(n_1809),
.C(n_1816),
.Y(n_1837)
);

NAND4xp75_ASAP7_75t_L g1838 ( 
.A(n_1829),
.B(n_1820),
.C(n_1810),
.D(n_1715),
.Y(n_1838)
);

OAI21xp33_ASAP7_75t_SL g1839 ( 
.A1(n_1830),
.A2(n_1820),
.B(n_1727),
.Y(n_1839)
);

NAND2x1p5_ASAP7_75t_L g1840 ( 
.A(n_1823),
.B(n_1810),
.Y(n_1840)
);

NOR4xp25_ASAP7_75t_L g1841 ( 
.A(n_1825),
.B(n_1727),
.C(n_1653),
.D(n_1730),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1822),
.Y(n_1842)
);

AOI21xp33_ASAP7_75t_L g1843 ( 
.A1(n_1832),
.A2(n_1733),
.B(n_1731),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1841),
.B(n_1827),
.Y(n_1844)
);

OAI221xp5_ASAP7_75t_L g1845 ( 
.A1(n_1834),
.A2(n_1833),
.B1(n_1826),
.B2(n_1824),
.C(n_1694),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1842),
.B(n_1840),
.Y(n_1846)
);

O2A1O1Ixp33_ASAP7_75t_L g1847 ( 
.A1(n_1837),
.A2(n_1733),
.B(n_1731),
.C(n_1730),
.Y(n_1847)
);

NAND4xp25_ASAP7_75t_SL g1848 ( 
.A(n_1839),
.B(n_1726),
.C(n_1724),
.D(n_1604),
.Y(n_1848)
);

O2A1O1Ixp33_ASAP7_75t_L g1849 ( 
.A1(n_1836),
.A2(n_1733),
.B(n_1726),
.C(n_1724),
.Y(n_1849)
);

AND4x1_ASAP7_75t_L g1850 ( 
.A(n_1846),
.B(n_1835),
.C(n_1838),
.D(n_1843),
.Y(n_1850)
);

AOI221xp5_ASAP7_75t_L g1851 ( 
.A1(n_1844),
.A2(n_1689),
.B1(n_1624),
.B2(n_1657),
.C(n_1656),
.Y(n_1851)
);

HB1xp67_ASAP7_75t_L g1852 ( 
.A(n_1848),
.Y(n_1852)
);

OAI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1845),
.A2(n_1643),
.B1(n_1646),
.B2(n_1593),
.Y(n_1853)
);

AOI211xp5_ASAP7_75t_L g1854 ( 
.A1(n_1847),
.A2(n_1611),
.B(n_1527),
.C(n_1605),
.Y(n_1854)
);

AO21x2_ASAP7_75t_L g1855 ( 
.A1(n_1849),
.A2(n_1676),
.B(n_1675),
.Y(n_1855)
);

NAND3xp33_ASAP7_75t_L g1856 ( 
.A(n_1844),
.B(n_1646),
.C(n_1601),
.Y(n_1856)
);

AO22x2_ASAP7_75t_L g1857 ( 
.A1(n_1856),
.A2(n_1676),
.B1(n_1675),
.B2(n_1667),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1852),
.Y(n_1858)
);

NOR2x1_ASAP7_75t_L g1859 ( 
.A(n_1853),
.B(n_1667),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1850),
.B(n_1673),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1855),
.Y(n_1861)
);

NAND4xp75_ASAP7_75t_L g1862 ( 
.A(n_1858),
.B(n_1851),
.C(n_1854),
.D(n_1460),
.Y(n_1862)
);

OAI322xp33_ASAP7_75t_L g1863 ( 
.A1(n_1860),
.A2(n_1623),
.A3(n_1621),
.B1(n_1619),
.B2(n_1657),
.C1(n_1656),
.C2(n_1675),
.Y(n_1863)
);

AOI32xp33_ASAP7_75t_L g1864 ( 
.A1(n_1861),
.A2(n_1683),
.A3(n_1661),
.B1(n_1670),
.B2(n_1669),
.Y(n_1864)
);

HB1xp67_ASAP7_75t_L g1865 ( 
.A(n_1862),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1865),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1866),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1866),
.Y(n_1868)
);

AOI21x1_ASAP7_75t_L g1869 ( 
.A1(n_1868),
.A2(n_1857),
.B(n_1859),
.Y(n_1869)
);

XNOR2x1_ASAP7_75t_L g1870 ( 
.A(n_1867),
.B(n_1864),
.Y(n_1870)
);

OAI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1870),
.A2(n_1863),
.B1(n_1667),
.B2(n_1676),
.Y(n_1871)
);

OAI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1869),
.A2(n_1683),
.B(n_1670),
.Y(n_1872)
);

XOR2xp5_ASAP7_75t_L g1873 ( 
.A(n_1871),
.B(n_1460),
.Y(n_1873)
);

OAI21xp5_ASAP7_75t_SL g1874 ( 
.A1(n_1873),
.A2(n_1872),
.B(n_1529),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1874),
.Y(n_1875)
);

OAI221xp5_ASAP7_75t_R g1876 ( 
.A1(n_1875),
.A2(n_1460),
.B1(n_1528),
.B2(n_1548),
.C(n_1627),
.Y(n_1876)
);

AOI211xp5_ASAP7_75t_L g1877 ( 
.A1(n_1876),
.A2(n_1529),
.B(n_1556),
.C(n_1514),
.Y(n_1877)
);


endmodule