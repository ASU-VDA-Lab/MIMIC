module fake_netlist_6_3068_n_1668 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1668);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1668;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_46),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_103),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_96),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_108),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_83),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_43),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_105),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_85),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_116),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_91),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_86),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_6),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_134),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_46),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_14),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_112),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_9),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_109),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_73),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_13),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_106),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_17),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_84),
.Y(n_183)
);

BUFx10_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_10),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_36),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_154),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_87),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_94),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_6),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_19),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_4),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_123),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_35),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_5),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_118),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_28),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_9),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_75),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_49),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_98),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_21),
.Y(n_203)
);

INVxp33_ASAP7_75t_R g204 ( 
.A(n_120),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_13),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_115),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_58),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_101),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_135),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_144),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_113),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_63),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_19),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_130),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_136),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_52),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_53),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_110),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_56),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_21),
.Y(n_220)
);

HB1xp67_ASAP7_75t_SL g221 ( 
.A(n_31),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_20),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_20),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_33),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_53),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_140),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_8),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_57),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_138),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_127),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_61),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_4),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_23),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_40),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_28),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_133),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_57),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_36),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_148),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_23),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_24),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_49),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_95),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_89),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_80),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_50),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_117),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_114),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_35),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_31),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_5),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_1),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_93),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_16),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_159),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_67),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_125),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_82),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_48),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_104),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_29),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_97),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_14),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_40),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_88),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_143),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_77),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_129),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_107),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_45),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_37),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_30),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_26),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_72),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_11),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_43),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_47),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_81),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_33),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_7),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_146),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_55),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_153),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_41),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_22),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_119),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_90),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_62),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_29),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_100),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_51),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_149),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_17),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_64),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_56),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_139),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_131),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_10),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_39),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_47),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_38),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_50),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_158),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_66),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_48),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_12),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_15),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_26),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_22),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_150),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_27),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_24),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_51),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_37),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_55),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_11),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_121),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_27),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_222),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_161),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_167),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_162),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_222),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_222),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_163),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_164),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_222),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_218),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_245),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_165),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_256),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_238),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_222),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_312),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_181),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_169),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_173),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_230),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_221),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_178),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_312),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_179),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_297),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_183),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_312),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_187),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_312),
.Y(n_347)
);

INVxp33_ASAP7_75t_SL g348 ( 
.A(n_201),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_189),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_197),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_312),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_200),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_202),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_242),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_206),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_241),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_205),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_207),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_208),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_211),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_242),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_214),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_174),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_174),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_175),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_226),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_229),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_168),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_241),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_175),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_231),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_244),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_255),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_180),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_180),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_185),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_168),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_185),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_258),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_195),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_165),
.B(n_0),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_195),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_166),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_171),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_199),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_199),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_170),
.B(n_0),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_260),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_216),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_266),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_170),
.B(n_1),
.Y(n_391)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_288),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_274),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_216),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_322),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_319),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_325),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_323),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_323),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_320),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_319),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_326),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_321),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_324),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_331),
.B(n_256),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_324),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_327),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_327),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_333),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_333),
.Y(n_410)
);

BUFx8_ASAP7_75t_L g411 ( 
.A(n_331),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_334),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_334),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_339),
.Y(n_414)
);

NAND2xp33_ASAP7_75t_L g415 ( 
.A(n_381),
.B(n_172),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_341),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_336),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_392),
.A2(n_160),
.B1(n_182),
.B2(n_196),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_341),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_345),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_345),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_347),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_347),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_351),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_351),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_330),
.B(n_288),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_337),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_340),
.B(n_342),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_368),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_350),
.B(n_210),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_353),
.B(n_210),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_363),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_355),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_368),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_377),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_335),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_339),
.B(n_184),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_363),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_369),
.A2(n_220),
.B1(n_235),
.B2(n_282),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_364),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_358),
.B(n_194),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_359),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_364),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_332),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_365),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_360),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_367),
.B(n_257),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_377),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_L g449 ( 
.A(n_354),
.B(n_243),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_384),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_365),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_371),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_370),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_373),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_370),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_374),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_374),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_384),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_388),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_375),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_375),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_331),
.Y(n_462)
);

AND2x6_ASAP7_75t_L g463 ( 
.A(n_331),
.B(n_257),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_331),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_390),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_348),
.A2(n_387),
.B1(n_391),
.B2(n_329),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_396),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_441),
.B(n_357),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_444),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_466),
.B(n_357),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_439),
.B(n_332),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_426),
.B(n_328),
.Y(n_472)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_405),
.B(n_171),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_405),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_405),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_430),
.B(n_383),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_405),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g478 ( 
.A1(n_426),
.A2(n_356),
.B1(n_213),
.B2(n_240),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_431),
.A2(n_213),
.B1(n_270),
.B2(n_224),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_432),
.B(n_354),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_411),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_414),
.Y(n_482)
);

OAI22xp33_ASAP7_75t_L g483 ( 
.A1(n_466),
.A2(n_251),
.B1(n_223),
.B2(n_219),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_462),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_432),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_437),
.A2(n_362),
.B1(n_393),
.B2(n_379),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_406),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_395),
.B(n_344),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_447),
.B(n_248),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_397),
.B(n_346),
.Y(n_490)
);

NAND2xp33_ASAP7_75t_L g491 ( 
.A(n_463),
.B(n_176),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_411),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_438),
.B(n_176),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_439),
.B(n_376),
.Y(n_494)
);

NAND2x1p5_ASAP7_75t_L g495 ( 
.A(n_464),
.B(n_188),
.Y(n_495)
);

INVx5_ASAP7_75t_L g496 ( 
.A(n_463),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_398),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_406),
.Y(n_498)
);

BUFx4f_ASAP7_75t_L g499 ( 
.A(n_463),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_406),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_464),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_398),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_413),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_402),
.B(n_349),
.Y(n_504)
);

INVx4_ASAP7_75t_SL g505 ( 
.A(n_463),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_413),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_411),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_396),
.Y(n_508)
);

NAND2x1p5_ASAP7_75t_L g509 ( 
.A(n_464),
.B(n_188),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_428),
.B(n_352),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_413),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_440),
.B(n_376),
.Y(n_512)
);

NOR3xp33_ASAP7_75t_L g513 ( 
.A(n_418),
.B(n_300),
.C(n_269),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_449),
.Y(n_514)
);

AND2x6_ASAP7_75t_L g515 ( 
.A(n_464),
.B(n_209),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_399),
.B(n_404),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_440),
.B(n_209),
.Y(n_517)
);

AND2x6_ASAP7_75t_L g518 ( 
.A(n_443),
.B(n_212),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_416),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_445),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_445),
.B(n_361),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_415),
.A2(n_224),
.B1(n_232),
.B2(n_308),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_451),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_465),
.B(n_417),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_451),
.B(n_212),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_400),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_427),
.A2(n_372),
.B1(n_366),
.B2(n_343),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_433),
.B(n_184),
.Y(n_528)
);

INVxp67_ASAP7_75t_SL g529 ( 
.A(n_462),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_442),
.B(n_338),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_463),
.A2(n_237),
.B1(n_232),
.B2(n_308),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_453),
.B(n_361),
.Y(n_532)
);

NOR3xp33_ASAP7_75t_L g533 ( 
.A(n_418),
.B(n_265),
.C(n_186),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_462),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_416),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_453),
.B(n_378),
.Y(n_536)
);

NAND2x1p5_ASAP7_75t_L g537 ( 
.A(n_462),
.B(n_215),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_399),
.B(n_278),
.Y(n_538)
);

AND2x6_ASAP7_75t_L g539 ( 
.A(n_455),
.B(n_215),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_449),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_446),
.B(n_204),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_403),
.Y(n_542)
);

BUFx10_ASAP7_75t_L g543 ( 
.A(n_452),
.Y(n_543)
);

AND2x6_ASAP7_75t_L g544 ( 
.A(n_455),
.B(n_236),
.Y(n_544)
);

AND2x2_ASAP7_75t_SL g545 ( 
.A(n_456),
.B(n_236),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_SL g546 ( 
.A(n_454),
.B(n_177),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_404),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_462),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_408),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_436),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_456),
.Y(n_551)
);

BUFx10_ASAP7_75t_L g552 ( 
.A(n_459),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_416),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_424),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_408),
.B(n_286),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_409),
.B(n_410),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_457),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_409),
.B(n_287),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_L g559 ( 
.A(n_463),
.B(n_239),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_424),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_424),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_463),
.A2(n_292),
.B1(n_294),
.B2(n_296),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_410),
.B(n_303),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_429),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_457),
.B(n_190),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_460),
.B(n_192),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_460),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_461),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_461),
.B(n_193),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_419),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_419),
.B(n_304),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_429),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_420),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_420),
.B(n_378),
.Y(n_574)
);

AND2x6_ASAP7_75t_L g575 ( 
.A(n_421),
.B(n_239),
.Y(n_575)
);

NOR2x1p5_ASAP7_75t_L g576 ( 
.A(n_421),
.B(n_198),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_423),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_422),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_422),
.B(n_380),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_435),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_458),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_458),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_425),
.B(n_310),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_425),
.B(n_407),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_435),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_407),
.B(n_203),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_435),
.B(n_380),
.Y(n_587)
);

NOR2x1p5_ASAP7_75t_L g588 ( 
.A(n_434),
.B(n_217),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_458),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_448),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_448),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_411),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_448),
.B(n_382),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_396),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_458),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_463),
.A2(n_275),
.B1(n_237),
.B2(n_240),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_450),
.B(n_382),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_450),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_458),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_458),
.Y(n_600)
);

OAI22xp33_ASAP7_75t_L g601 ( 
.A1(n_450),
.A2(n_234),
.B1(n_233),
.B2(n_228),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_396),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_407),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_407),
.Y(n_604)
);

OR2x6_ASAP7_75t_L g605 ( 
.A(n_434),
.B(n_246),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_396),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_396),
.Y(n_607)
);

INVx4_ASAP7_75t_SL g608 ( 
.A(n_401),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_412),
.B(n_225),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_412),
.Y(n_610)
);

INVx6_ASAP7_75t_L g611 ( 
.A(n_401),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_423),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_476),
.B(n_227),
.Y(n_613)
);

AOI22x1_ASAP7_75t_SL g614 ( 
.A1(n_485),
.A2(n_249),
.B1(n_252),
.B2(n_254),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_L g615 ( 
.A(n_473),
.B(n_247),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_489),
.B(n_250),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_545),
.B(n_247),
.Y(n_617)
);

NOR2xp67_ASAP7_75t_L g618 ( 
.A(n_527),
.B(n_412),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_477),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_477),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_474),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_543),
.Y(n_622)
);

NAND2x1_ASAP7_75t_L g623 ( 
.A(n_611),
.B(n_412),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_475),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_545),
.B(n_253),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_472),
.A2(n_290),
.B1(n_283),
.B2(n_317),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_468),
.B(n_264),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_494),
.A2(n_280),
.B1(n_279),
.B2(n_276),
.Y(n_628)
);

NAND2x1p5_ASAP7_75t_L g629 ( 
.A(n_499),
.B(n_253),
.Y(n_629)
);

NOR3xp33_ASAP7_75t_L g630 ( 
.A(n_470),
.B(n_291),
.C(n_271),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_471),
.B(n_469),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_499),
.B(n_262),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_536),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_586),
.B(n_423),
.Y(n_634)
);

NAND2x1_ASAP7_75t_L g635 ( 
.A(n_611),
.B(n_401),
.Y(n_635)
);

NOR2xp67_ASAP7_75t_SL g636 ( 
.A(n_481),
.B(n_262),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_499),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_472),
.B(n_184),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_514),
.B(n_540),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_543),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_510),
.B(n_205),
.Y(n_641)
);

OAI22xp33_ASAP7_75t_L g642 ( 
.A1(n_494),
.A2(n_290),
.B1(n_267),
.B2(n_268),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_609),
.B(n_423),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_483),
.B(n_272),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_520),
.B(n_401),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_536),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_518),
.A2(n_544),
.B1(n_539),
.B2(n_575),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_523),
.B(n_267),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_551),
.B(n_268),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_564),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_L g651 ( 
.A(n_473),
.B(n_281),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_518),
.A2(n_270),
.B1(n_298),
.B2(n_299),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_522),
.A2(n_281),
.B1(n_283),
.B2(n_317),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_557),
.B(n_385),
.Y(n_654)
);

A2O1A1Ixp33_ASAP7_75t_L g655 ( 
.A1(n_567),
.A2(n_275),
.B(n_302),
.C(n_298),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_473),
.Y(n_656)
);

AO221x1_ASAP7_75t_L g657 ( 
.A1(n_601),
.A2(n_279),
.B1(n_246),
.B2(n_259),
.C(n_261),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_568),
.B(n_385),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_497),
.B(n_386),
.Y(n_659)
);

NAND2xp33_ASAP7_75t_L g660 ( 
.A(n_473),
.B(n_518),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_528),
.B(n_538),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_480),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_497),
.B(n_386),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_543),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_565),
.B(n_184),
.Y(n_665)
);

A2O1A1Ixp33_ASAP7_75t_L g666 ( 
.A1(n_566),
.A2(n_299),
.B(n_306),
.C(n_259),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_480),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_502),
.B(n_389),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_552),
.B(n_205),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_SL g670 ( 
.A1(n_541),
.A2(n_191),
.B1(n_205),
.B2(n_261),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_518),
.A2(n_302),
.B1(n_263),
.B2(n_276),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_569),
.B(n_191),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_572),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_576),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_502),
.B(n_547),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_572),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_521),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_580),
.Y(n_678)
);

O2A1O1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_512),
.A2(n_263),
.B(n_280),
.C(n_306),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_481),
.B(n_191),
.Y(n_680)
);

NAND3xp33_ASAP7_75t_L g681 ( 
.A(n_478),
.B(n_305),
.C(n_273),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_580),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_521),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_547),
.B(n_389),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_585),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_471),
.B(n_482),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_532),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_549),
.B(n_394),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_555),
.B(n_277),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_558),
.B(n_284),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_549),
.B(n_394),
.Y(n_691)
);

NOR2xp67_ASAP7_75t_L g692 ( 
.A(n_486),
.B(n_92),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_570),
.B(n_318),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_532),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_585),
.Y(n_695)
);

BUFx6f_ASAP7_75t_SL g696 ( 
.A(n_552),
.Y(n_696)
);

NOR3xp33_ASAP7_75t_L g697 ( 
.A(n_546),
.B(n_316),
.C(n_315),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_570),
.B(n_314),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_512),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_574),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_573),
.B(n_313),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_590),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_588),
.Y(n_703)
);

OAI221xp5_ASAP7_75t_L g704 ( 
.A1(n_479),
.A2(n_311),
.B1(n_309),
.B2(n_307),
.C(n_301),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_573),
.B(n_295),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_SL g706 ( 
.A(n_552),
.B(n_530),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_578),
.B(n_293),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_590),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_546),
.A2(n_191),
.B1(n_289),
.B2(n_285),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_496),
.B(n_68),
.Y(n_710)
);

AOI221xp5_ASAP7_75t_L g711 ( 
.A1(n_513),
.A2(n_2),
.B1(n_3),
.B2(n_7),
.C(n_8),
.Y(n_711)
);

NOR2xp67_ASAP7_75t_L g712 ( 
.A(n_524),
.B(n_70),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_488),
.B(n_2),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_578),
.B(n_71),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_591),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_SL g716 ( 
.A(n_526),
.B(n_3),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_584),
.B(n_74),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_563),
.B(n_69),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_571),
.B(n_12),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_L g720 ( 
.A(n_473),
.B(n_76),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_490),
.B(n_15),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_496),
.B(n_78),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_526),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_591),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_473),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_493),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_583),
.B(n_79),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_598),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_610),
.B(n_65),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_610),
.B(n_99),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_518),
.A2(n_60),
.B1(n_157),
.B2(n_156),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_501),
.B(n_59),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_598),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_516),
.B(n_155),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_496),
.B(n_152),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_587),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_SL g737 ( 
.A1(n_542),
.A2(n_16),
.B1(n_18),
.B2(n_25),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_556),
.B(n_587),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_493),
.B(n_18),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_593),
.B(n_151),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_504),
.B(n_25),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_542),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_529),
.A2(n_145),
.B(n_142),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_593),
.B(n_141),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_518),
.A2(n_137),
.B1(n_132),
.B2(n_128),
.Y(n_745)
);

NAND3xp33_ASAP7_75t_SL g746 ( 
.A(n_533),
.B(n_30),
.C(n_32),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_539),
.A2(n_32),
.B1(n_34),
.B2(n_38),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_550),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_597),
.B(n_124),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_539),
.A2(n_122),
.B1(n_102),
.B2(n_41),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_574),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_579),
.B(n_493),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_492),
.B(n_54),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_579),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_495),
.A2(n_34),
.B1(n_39),
.B2(n_42),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_597),
.B(n_54),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_496),
.B(n_42),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_605),
.Y(n_758)
);

BUFx6f_ASAP7_75t_SL g759 ( 
.A(n_517),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_487),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_517),
.B(n_44),
.Y(n_761)
);

OAI22xp33_ASAP7_75t_L g762 ( 
.A1(n_605),
.A2(n_44),
.B1(n_45),
.B2(n_52),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_517),
.B(n_525),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_525),
.B(n_603),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_539),
.A2(n_544),
.B1(n_575),
.B2(n_525),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_603),
.B(n_604),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_604),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_492),
.B(n_592),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_605),
.B(n_600),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_595),
.B(n_599),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_487),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_496),
.B(n_509),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_498),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_599),
.B(n_539),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_616),
.B(n_539),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_764),
.A2(n_607),
.B(n_606),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_641),
.B(n_495),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_613),
.B(n_495),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_763),
.A2(n_589),
.B(n_491),
.Y(n_779)
);

CKINVDCx8_ASAP7_75t_R g780 ( 
.A(n_723),
.Y(n_780)
);

O2A1O1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_617),
.A2(n_625),
.B(n_642),
.C(n_756),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_616),
.B(n_544),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_613),
.B(n_507),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_706),
.B(n_592),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_763),
.A2(n_559),
.B(n_491),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_661),
.A2(n_544),
.B1(n_575),
.B2(n_515),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_742),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_736),
.A2(n_765),
.B1(n_726),
.B2(n_661),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_634),
.A2(n_559),
.B(n_612),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_631),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_633),
.B(n_505),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_736),
.B(n_544),
.Y(n_792)
);

A2O1A1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_719),
.A2(n_562),
.B(n_507),
.C(n_596),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_643),
.A2(n_484),
.B(n_534),
.Y(n_794)
);

NOR2xp67_ASAP7_75t_L g795 ( 
.A(n_622),
.B(n_640),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_689),
.A2(n_575),
.B1(n_515),
.B2(n_509),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_689),
.B(n_575),
.Y(n_797)
);

OAI21xp5_ASAP7_75t_L g798 ( 
.A1(n_766),
.A2(n_509),
.B(n_553),
.Y(n_798)
);

AO21x1_ASAP7_75t_L g799 ( 
.A1(n_617),
.A2(n_537),
.B(n_612),
.Y(n_799)
);

A2O1A1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_719),
.A2(n_531),
.B(n_594),
.C(n_467),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_621),
.Y(n_801)
);

A2O1A1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_644),
.A2(n_467),
.B(n_594),
.C(n_508),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_690),
.B(n_575),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_SL g804 ( 
.A(n_696),
.B(n_515),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_660),
.A2(n_548),
.B(n_612),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_686),
.B(n_537),
.Y(n_806)
);

INVx4_ASAP7_75t_L g807 ( 
.A(n_620),
.Y(n_807)
);

OAI321xp33_ASAP7_75t_L g808 ( 
.A1(n_762),
.A2(n_711),
.A3(n_644),
.B1(n_737),
.B2(n_747),
.C(n_746),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_772),
.A2(n_548),
.B(n_577),
.Y(n_809)
);

A2O1A1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_627),
.A2(n_467),
.B(n_594),
.C(n_508),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_772),
.A2(n_577),
.B(n_582),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_765),
.A2(n_537),
.B1(n_508),
.B2(n_611),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_624),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_774),
.A2(n_577),
.B(n_582),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_690),
.B(n_515),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_650),
.Y(n_816)
);

BUFx12f_ASAP7_75t_L g817 ( 
.A(n_674),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_675),
.B(n_515),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_627),
.A2(n_498),
.B(n_500),
.C(n_503),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_650),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_646),
.B(n_515),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_696),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_748),
.B(n_582),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_700),
.B(n_500),
.Y(n_824)
);

BUFx12f_ASAP7_75t_L g825 ( 
.A(n_703),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_639),
.B(n_582),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_751),
.B(n_503),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_754),
.B(n_662),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_713),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_740),
.A2(n_581),
.B(n_602),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_667),
.B(n_554),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_677),
.B(n_554),
.Y(n_832)
);

OAI321xp33_ASAP7_75t_L g833 ( 
.A1(n_747),
.A2(n_755),
.A3(n_625),
.B1(n_709),
.B2(n_628),
.C(n_626),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_744),
.A2(n_749),
.B(n_619),
.Y(n_834)
);

NOR2x1p5_ASAP7_75t_SL g835 ( 
.A(n_760),
.B(n_553),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_699),
.B(n_560),
.Y(n_836)
);

INVx1_ASAP7_75t_SL g837 ( 
.A(n_721),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_619),
.A2(n_581),
.B(n_602),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_620),
.B(n_505),
.Y(n_839)
);

NAND3xp33_ASAP7_75t_L g840 ( 
.A(n_670),
.B(n_535),
.C(n_506),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_683),
.B(n_535),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_687),
.B(n_505),
.Y(n_842)
);

INVx5_ASAP7_75t_L g843 ( 
.A(n_656),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_694),
.B(n_693),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_717),
.A2(n_602),
.B(n_506),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_698),
.B(n_511),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_739),
.A2(n_511),
.B(n_519),
.C(n_560),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_669),
.B(n_519),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_701),
.B(n_561),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_632),
.A2(n_561),
.B(n_505),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_664),
.B(n_608),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_705),
.B(n_707),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_659),
.B(n_663),
.Y(n_853)
);

OAI21xp33_ASAP7_75t_L g854 ( 
.A1(n_628),
.A2(n_608),
.B(n_716),
.Y(n_854)
);

O2A1O1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_666),
.A2(n_653),
.B(n_757),
.C(n_648),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_770),
.A2(n_608),
.B(n_769),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_668),
.B(n_608),
.Y(n_857)
);

NOR2x1p5_ASAP7_75t_SL g858 ( 
.A(n_760),
.B(n_773),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_647),
.A2(n_620),
.B1(n_629),
.B2(n_769),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_645),
.A2(n_734),
.B(n_770),
.Y(n_860)
);

NAND2x1p5_ASAP7_75t_L g861 ( 
.A(n_725),
.B(n_620),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_638),
.B(n_741),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_623),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_718),
.A2(n_727),
.B(n_615),
.Y(n_864)
);

AOI22x1_ASAP7_75t_L g865 ( 
.A1(n_629),
.A2(n_767),
.B1(n_773),
.B2(n_702),
.Y(n_865)
);

BUFx2_ASAP7_75t_L g866 ( 
.A(n_758),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_758),
.B(n_618),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_651),
.A2(n_720),
.B(n_714),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_758),
.B(n_692),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_732),
.A2(n_771),
.B(n_729),
.Y(n_870)
);

NAND3xp33_ASAP7_75t_SL g871 ( 
.A(n_697),
.B(n_630),
.C(n_704),
.Y(n_871)
);

OAI21x1_ASAP7_75t_L g872 ( 
.A1(n_673),
.A2(n_695),
.B(n_715),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_R g873 ( 
.A(n_759),
.B(n_758),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_673),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_665),
.A2(n_672),
.B1(n_759),
.B2(n_761),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_657),
.A2(n_739),
.B1(n_761),
.B2(n_652),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_681),
.B(n_658),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_684),
.B(n_691),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_652),
.A2(n_671),
.B1(n_725),
.B2(n_712),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_730),
.A2(n_708),
.B(n_728),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_688),
.B(n_649),
.Y(n_881)
);

OAI22x1_ASAP7_75t_L g882 ( 
.A1(n_753),
.A2(n_680),
.B1(n_768),
.B2(n_750),
.Y(n_882)
);

A2O1A1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_679),
.A2(n_654),
.B(n_671),
.C(n_728),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_725),
.B(n_708),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_676),
.A2(n_685),
.B(n_724),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_678),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_678),
.A2(n_715),
.B(n_733),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_682),
.B(n_724),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_SL g889 ( 
.A(n_636),
.B(n_655),
.Y(n_889)
);

NAND2xp33_ASAP7_75t_L g890 ( 
.A(n_682),
.B(n_685),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_695),
.B(n_635),
.Y(n_891)
);

OAI21xp5_ASAP7_75t_L g892 ( 
.A1(n_710),
.A2(n_722),
.B(n_735),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_710),
.A2(n_722),
.B(n_735),
.Y(n_893)
);

INVx5_ASAP7_75t_L g894 ( 
.A(n_731),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_743),
.A2(n_745),
.B(n_614),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_738),
.B(n_616),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_613),
.B(n_510),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_738),
.B(n_616),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_706),
.B(n_661),
.Y(n_899)
);

BUFx4f_ASAP7_75t_L g900 ( 
.A(n_758),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_738),
.A2(n_764),
.B(n_763),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_764),
.A2(n_738),
.B(n_766),
.Y(n_902)
);

AO22x1_ASAP7_75t_L g903 ( 
.A1(n_644),
.A2(n_533),
.B1(n_513),
.B2(n_627),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_613),
.B(n_510),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_736),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_613),
.B(n_510),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_641),
.B(n_472),
.Y(n_907)
);

A2O1A1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_763),
.A2(n_616),
.B(n_613),
.C(n_661),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_738),
.B(n_616),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_738),
.A2(n_764),
.B(n_763),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_738),
.B(n_616),
.Y(n_911)
);

NOR3xp33_ASAP7_75t_L g912 ( 
.A(n_644),
.B(n_339),
.C(n_541),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_738),
.A2(n_764),
.B(n_763),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_622),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_706),
.B(n_661),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_620),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_738),
.B(n_616),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_738),
.B(n_616),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_641),
.B(n_472),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_738),
.B(n_616),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_736),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_764),
.A2(n_738),
.B(n_766),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_764),
.A2(n_738),
.B(n_766),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_706),
.B(n_661),
.Y(n_924)
);

NAND2xp33_ASAP7_75t_L g925 ( 
.A(n_637),
.B(n_656),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_738),
.A2(n_764),
.B(n_763),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_R g927 ( 
.A(n_622),
.B(n_400),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_764),
.A2(n_738),
.B(n_766),
.Y(n_928)
);

OAI21x1_ASAP7_75t_L g929 ( 
.A1(n_774),
.A2(n_766),
.B(n_764),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_736),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_738),
.B(n_616),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_613),
.B(n_510),
.Y(n_932)
);

INVx4_ASAP7_75t_L g933 ( 
.A(n_620),
.Y(n_933)
);

AOI21xp33_ASAP7_75t_L g934 ( 
.A1(n_613),
.A2(n_644),
.B(n_616),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_738),
.A2(n_764),
.B(n_763),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_661),
.A2(n_763),
.B1(n_752),
.B2(n_690),
.Y(n_936)
);

BUFx10_ASAP7_75t_L g937 ( 
.A(n_696),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_738),
.B(n_616),
.Y(n_938)
);

NOR2xp67_ASAP7_75t_L g939 ( 
.A(n_622),
.B(n_640),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_613),
.B(n_510),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_763),
.A2(n_738),
.B1(n_736),
.B2(n_765),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_738),
.B(n_616),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_738),
.A2(n_764),
.B(n_763),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_738),
.A2(n_764),
.B(n_763),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_622),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_934),
.A2(n_904),
.B1(n_906),
.B2(n_897),
.Y(n_946)
);

NOR2xp67_ASAP7_75t_L g947 ( 
.A(n_914),
.B(n_795),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_905),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_834),
.A2(n_868),
.B(n_902),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_868),
.A2(n_923),
.B(n_922),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_896),
.B(n_898),
.Y(n_951)
);

AO31x2_ASAP7_75t_L g952 ( 
.A1(n_802),
.A2(n_799),
.A3(n_810),
.B(n_847),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_928),
.A2(n_910),
.B(n_901),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_927),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_901),
.A2(n_913),
.B(n_910),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_913),
.A2(n_935),
.B(n_926),
.Y(n_956)
);

AOI21xp33_ASAP7_75t_L g957 ( 
.A1(n_932),
.A2(n_940),
.B(n_781),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_909),
.B(n_911),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_916),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_790),
.B(n_907),
.Y(n_960)
);

OAI21x1_ASAP7_75t_L g961 ( 
.A1(n_880),
.A2(n_845),
.B(n_929),
.Y(n_961)
);

NOR2x1p5_ASAP7_75t_L g962 ( 
.A(n_817),
.B(n_825),
.Y(n_962)
);

NAND2x1p5_ASAP7_75t_L g963 ( 
.A(n_843),
.B(n_900),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_874),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_943),
.A2(n_944),
.B(n_798),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_921),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_780),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_944),
.A2(n_918),
.B(n_917),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_899),
.A2(n_915),
.B1(n_924),
.B2(n_919),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_945),
.Y(n_970)
);

AOI21xp33_ASAP7_75t_L g971 ( 
.A1(n_833),
.A2(n_931),
.B(n_920),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_938),
.B(n_942),
.Y(n_972)
);

OAI21x1_ASAP7_75t_L g973 ( 
.A1(n_814),
.A2(n_887),
.B(n_885),
.Y(n_973)
);

NOR2xp67_ASAP7_75t_L g974 ( 
.A(n_939),
.B(n_871),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_916),
.Y(n_975)
);

INVxp67_ASAP7_75t_L g976 ( 
.A(n_787),
.Y(n_976)
);

AOI21xp33_ASAP7_75t_L g977 ( 
.A1(n_808),
.A2(n_908),
.B(n_862),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_801),
.Y(n_978)
);

NAND2x1p5_ASAP7_75t_L g979 ( 
.A(n_843),
.B(n_900),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_797),
.A2(n_803),
.B(n_864),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_864),
.A2(n_805),
.B(n_925),
.Y(n_981)
);

AOI221xp5_ASAP7_75t_L g982 ( 
.A1(n_903),
.A2(n_912),
.B1(n_876),
.B2(n_844),
.C(n_882),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_936),
.B(n_852),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_813),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_829),
.B(n_837),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_853),
.B(n_878),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_855),
.A2(n_893),
.B(n_783),
.C(n_892),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_941),
.A2(n_893),
.B(n_785),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_815),
.A2(n_794),
.B(n_789),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_789),
.A2(n_775),
.B(n_782),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_776),
.A2(n_811),
.B(n_865),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_930),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_828),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_894),
.A2(n_854),
.B1(n_788),
.B2(n_879),
.Y(n_994)
);

OAI22x1_ASAP7_75t_L g995 ( 
.A1(n_875),
.A2(n_784),
.B1(n_894),
.B2(n_828),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_860),
.A2(n_818),
.B(n_785),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_806),
.B(n_848),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_894),
.A2(n_859),
.B1(n_786),
.B2(n_796),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_860),
.A2(n_881),
.B(n_809),
.Y(n_999)
);

NAND3xp33_ASAP7_75t_L g1000 ( 
.A(n_877),
.B(n_826),
.C(n_777),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_778),
.B(n_846),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_779),
.A2(n_800),
.B(n_792),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_836),
.B(n_866),
.Y(n_1003)
);

INVx1_ASAP7_75t_SL g1004 ( 
.A(n_873),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_849),
.B(n_824),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_SL g1006 ( 
.A1(n_895),
.A2(n_821),
.B(n_856),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_823),
.B(n_867),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_870),
.A2(n_812),
.B(n_838),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_827),
.B(n_832),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_779),
.A2(n_890),
.B(n_857),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_819),
.A2(n_883),
.B(n_793),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_869),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_884),
.A2(n_888),
.B(n_843),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_869),
.B(n_851),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_831),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_840),
.A2(n_850),
.B(n_841),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_874),
.B(n_886),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_843),
.A2(n_894),
.B(n_891),
.Y(n_1018)
);

AND2x2_ASAP7_75t_SL g1019 ( 
.A(n_804),
.B(n_889),
.Y(n_1019)
);

NAND2x1_ASAP7_75t_L g1020 ( 
.A(n_807),
.B(n_933),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_839),
.A2(n_842),
.B(n_791),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_791),
.A2(n_842),
.B(n_863),
.Y(n_1022)
);

AND2x2_ASAP7_75t_SL g1023 ( 
.A(n_807),
.B(n_933),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_816),
.B(n_820),
.Y(n_1024)
);

NOR2xp67_ASAP7_75t_SL g1025 ( 
.A(n_822),
.B(n_863),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_861),
.A2(n_937),
.B1(n_858),
.B2(n_835),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_861),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_934),
.A2(n_908),
.B(n_901),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_934),
.A2(n_908),
.B(n_901),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_901),
.A2(n_913),
.B(n_910),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_901),
.A2(n_913),
.B(n_910),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_901),
.A2(n_913),
.B(n_910),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_896),
.B(n_898),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_874),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_896),
.B(n_898),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_905),
.Y(n_1036)
);

INVx5_ASAP7_75t_L g1037 ( 
.A(n_843),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_916),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_896),
.B(n_898),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_916),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_896),
.B(n_898),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_872),
.A2(n_880),
.B(n_830),
.Y(n_1042)
);

AOI21x1_ASAP7_75t_L g1043 ( 
.A1(n_901),
.A2(n_913),
.B(n_910),
.Y(n_1043)
);

BUFx12f_ASAP7_75t_L g1044 ( 
.A(n_937),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_896),
.B(n_898),
.Y(n_1045)
);

AO31x2_ASAP7_75t_L g1046 ( 
.A1(n_802),
.A2(n_799),
.A3(n_810),
.B(n_847),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_934),
.A2(n_908),
.B(n_901),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_897),
.B(n_940),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_828),
.B(n_866),
.Y(n_1049)
);

NAND2xp33_ASAP7_75t_L g1050 ( 
.A(n_908),
.B(n_637),
.Y(n_1050)
);

AOI21xp33_ASAP7_75t_L g1051 ( 
.A1(n_897),
.A2(n_906),
.B(n_904),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_872),
.A2(n_880),
.B(n_830),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_897),
.B(n_940),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_916),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_872),
.A2(n_880),
.B(n_830),
.Y(n_1055)
);

AOI21x1_ASAP7_75t_L g1056 ( 
.A1(n_901),
.A2(n_913),
.B(n_910),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_872),
.A2(n_880),
.B(n_830),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_934),
.B(n_940),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_872),
.A2(n_880),
.B(n_830),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_934),
.A2(n_908),
.B(n_901),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_897),
.B(n_940),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_791),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_896),
.B(n_898),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_872),
.A2(n_880),
.B(n_830),
.Y(n_1064)
);

AOI211x1_ASAP7_75t_L g1065 ( 
.A1(n_934),
.A2(n_903),
.B(n_642),
.C(n_844),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_927),
.Y(n_1066)
);

OAI22x1_ASAP7_75t_L g1067 ( 
.A1(n_897),
.A2(n_906),
.B1(n_932),
.B2(n_904),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_872),
.A2(n_880),
.B(n_830),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_825),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_934),
.A2(n_908),
.B(n_901),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_896),
.B(n_898),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_897),
.B(n_940),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_896),
.B(n_898),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_791),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_907),
.B(n_919),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_901),
.A2(n_913),
.B(n_910),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_1049),
.B(n_1014),
.Y(n_1077)
);

INVx4_ASAP7_75t_L g1078 ( 
.A(n_1037),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_1048),
.A2(n_1053),
.B1(n_1061),
.B2(n_1072),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1051),
.B(n_986),
.Y(n_1080)
);

NOR2xp67_ASAP7_75t_L g1081 ( 
.A(n_954),
.B(n_976),
.Y(n_1081)
);

OR2x6_ASAP7_75t_L g1082 ( 
.A(n_963),
.B(n_979),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_1049),
.B(n_1012),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_946),
.B(n_957),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_986),
.A2(n_972),
.B1(n_1041),
.B2(n_958),
.Y(n_1085)
);

BUFx4f_ASAP7_75t_L g1086 ( 
.A(n_1044),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_1037),
.Y(n_1087)
);

O2A1O1Ixp5_ASAP7_75t_SL g1088 ( 
.A1(n_957),
.A2(n_1058),
.B(n_977),
.C(n_1051),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_978),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_967),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_993),
.B(n_1062),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_1062),
.B(n_1074),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_984),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_1037),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_951),
.B(n_958),
.Y(n_1095)
);

OR2x6_ASAP7_75t_L g1096 ( 
.A(n_963),
.B(n_979),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_1033),
.A2(n_1035),
.B1(n_1045),
.B2(n_1073),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1033),
.B(n_1035),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_1074),
.B(n_1003),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_960),
.Y(n_1100)
);

AOI222xp33_ASAP7_75t_L g1101 ( 
.A1(n_1067),
.A2(n_982),
.B1(n_1075),
.B2(n_983),
.C1(n_1073),
.C2(n_1071),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1039),
.B(n_1045),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1063),
.A2(n_1071),
.B1(n_983),
.B2(n_987),
.Y(n_1103)
);

INVx4_ASAP7_75t_L g1104 ( 
.A(n_1037),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_968),
.A2(n_965),
.B(n_956),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_1066),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_970),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_955),
.A2(n_1076),
.B(n_1030),
.Y(n_1108)
);

OAI21xp33_ASAP7_75t_SL g1109 ( 
.A1(n_1019),
.A2(n_977),
.B(n_1063),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_997),
.B(n_1015),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_985),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_969),
.B(n_971),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_948),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_959),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1001),
.B(n_1005),
.Y(n_1115)
);

AOI222xp33_ASAP7_75t_L g1116 ( 
.A1(n_982),
.A2(n_994),
.B1(n_1070),
.B2(n_1028),
.C1(n_1029),
.C2(n_1060),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_1004),
.B(n_966),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_971),
.B(n_1001),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_1017),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_995),
.B(n_974),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1005),
.B(n_1009),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1009),
.B(n_1065),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_1007),
.B(n_1000),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_1069),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_947),
.A2(n_994),
.B1(n_998),
.B2(n_1050),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_959),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1036),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_992),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1047),
.B(n_988),
.Y(n_1129)
);

BUFx2_ASAP7_75t_SL g1130 ( 
.A(n_962),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_959),
.Y(n_1131)
);

AND2x2_ASAP7_75t_SL g1132 ( 
.A(n_1023),
.B(n_998),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1030),
.A2(n_1076),
.B(n_1031),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1021),
.A2(n_1011),
.B1(n_1022),
.B2(n_981),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1031),
.A2(n_1032),
.B(n_999),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1024),
.B(n_1032),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_975),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_964),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1026),
.A2(n_1018),
.B1(n_1017),
.B2(n_1008),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1034),
.B(n_1025),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1027),
.B(n_1038),
.Y(n_1141)
);

O2A1O1Ixp5_ASAP7_75t_L g1142 ( 
.A1(n_980),
.A2(n_989),
.B(n_990),
.C(n_1056),
.Y(n_1142)
);

BUFx8_ASAP7_75t_SL g1143 ( 
.A(n_975),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_1038),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_SL g1145 ( 
.A1(n_1020),
.A2(n_1038),
.B1(n_1054),
.B2(n_1040),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_1040),
.Y(n_1146)
);

AO21x2_ASAP7_75t_L g1147 ( 
.A1(n_996),
.A2(n_1006),
.B(n_1043),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_1054),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1010),
.A2(n_1002),
.B(n_1016),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1013),
.B(n_952),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_1046),
.Y(n_1151)
);

OR2x6_ASAP7_75t_L g1152 ( 
.A(n_973),
.B(n_991),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_1046),
.Y(n_1153)
);

INVx3_ASAP7_75t_SL g1154 ( 
.A(n_961),
.Y(n_1154)
);

INVxp67_ASAP7_75t_L g1155 ( 
.A(n_1042),
.Y(n_1155)
);

INVx2_ASAP7_75t_SL g1156 ( 
.A(n_1052),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1055),
.A2(n_1057),
.B(n_1059),
.C(n_1064),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1068),
.B(n_1048),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1048),
.B(n_1053),
.Y(n_1159)
);

O2A1O1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1051),
.A2(n_934),
.B(n_1053),
.C(n_1048),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_978),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_1037),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1048),
.B(n_1053),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_978),
.Y(n_1164)
);

INVxp67_ASAP7_75t_L g1165 ( 
.A(n_960),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_978),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1048),
.B(n_1053),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_978),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_978),
.Y(n_1169)
);

HB1xp67_ASAP7_75t_L g1170 ( 
.A(n_1003),
.Y(n_1170)
);

NAND3xp33_ASAP7_75t_SL g1171 ( 
.A(n_946),
.B(n_904),
.C(n_897),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1048),
.A2(n_1053),
.B1(n_1072),
.B2(n_1061),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1048),
.B(n_1053),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_1037),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_1049),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1048),
.A2(n_1053),
.B1(n_1072),
.B2(n_1061),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1048),
.B(n_1053),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1049),
.B(n_1014),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1048),
.B(n_1053),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_954),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_953),
.A2(n_950),
.B(n_949),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_978),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1048),
.B(n_1053),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_1037),
.Y(n_1184)
);

OR2x6_ASAP7_75t_L g1185 ( 
.A(n_963),
.B(n_979),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1048),
.B(n_1053),
.Y(n_1186)
);

INVx4_ASAP7_75t_L g1187 ( 
.A(n_1037),
.Y(n_1187)
);

AO32x2_ASAP7_75t_L g1188 ( 
.A1(n_994),
.A2(n_998),
.A3(n_788),
.B1(n_941),
.B2(n_755),
.Y(n_1188)
);

OR2x2_ASAP7_75t_L g1189 ( 
.A(n_960),
.B(n_790),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_946),
.B(n_934),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_1066),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1048),
.B(n_1053),
.Y(n_1192)
);

OA21x2_ASAP7_75t_L g1193 ( 
.A1(n_988),
.A2(n_1029),
.B(n_1028),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1049),
.B(n_1014),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1048),
.B(n_1053),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1048),
.B(n_1053),
.Y(n_1196)
);

HB1xp67_ASAP7_75t_L g1197 ( 
.A(n_1003),
.Y(n_1197)
);

OAI21xp33_ASAP7_75t_L g1198 ( 
.A1(n_1048),
.A2(n_1061),
.B(n_1053),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1048),
.B(n_1053),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_954),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_976),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1048),
.B(n_1053),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1049),
.B(n_1014),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1171),
.A2(n_1190),
.B1(n_1176),
.B2(n_1172),
.Y(n_1204)
);

AO21x2_ASAP7_75t_L g1205 ( 
.A1(n_1135),
.A2(n_1133),
.B(n_1157),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_1087),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_1180),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1171),
.A2(n_1190),
.B1(n_1173),
.B2(n_1198),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_1084),
.B(n_1129),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1173),
.A2(n_1079),
.B1(n_1084),
.B2(n_1101),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1163),
.B(n_1179),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1079),
.A2(n_1192),
.B1(n_1177),
.B2(n_1186),
.Y(n_1212)
);

CKINVDCx11_ASAP7_75t_R g1213 ( 
.A(n_1191),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1200),
.Y(n_1214)
);

BUFx4f_ASAP7_75t_SL g1215 ( 
.A(n_1126),
.Y(n_1215)
);

CKINVDCx11_ASAP7_75t_R g1216 ( 
.A(n_1107),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1166),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1170),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1182),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1093),
.Y(n_1220)
);

OR2x6_ASAP7_75t_L g1221 ( 
.A(n_1149),
.B(n_1134),
.Y(n_1221)
);

OR2x2_ASAP7_75t_L g1222 ( 
.A(n_1103),
.B(n_1193),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1170),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1197),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1161),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1193),
.B(n_1115),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1143),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_SL g1228 ( 
.A1(n_1160),
.A2(n_1167),
.B(n_1159),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1164),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1168),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1080),
.B(n_1095),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1183),
.B(n_1195),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1136),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1098),
.B(n_1102),
.Y(n_1234)
);

OAI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1110),
.A2(n_1125),
.B1(n_1121),
.B2(n_1085),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_1106),
.Y(n_1236)
);

BUFx4f_ASAP7_75t_SL g1237 ( 
.A(n_1124),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1169),
.Y(n_1238)
);

CKINVDCx11_ASAP7_75t_R g1239 ( 
.A(n_1090),
.Y(n_1239)
);

CKINVDCx6p67_ASAP7_75t_R g1240 ( 
.A(n_1130),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1197),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1196),
.A2(n_1199),
.B1(n_1202),
.B2(n_1097),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1132),
.A2(n_1123),
.B1(n_1112),
.B2(n_1116),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1087),
.Y(n_1244)
);

NAND2x1p5_ASAP7_75t_L g1245 ( 
.A(n_1132),
.B(n_1153),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1113),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1127),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1109),
.B(n_1118),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1128),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1160),
.B(n_1189),
.Y(n_1250)
);

OAI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1117),
.A2(n_1123),
.B1(n_1100),
.B2(n_1111),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1120),
.A2(n_1118),
.B1(n_1193),
.B2(n_1140),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1119),
.Y(n_1253)
);

AO21x1_ASAP7_75t_L g1254 ( 
.A1(n_1149),
.A2(n_1122),
.B(n_1139),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1138),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1165),
.A2(n_1099),
.B1(n_1201),
.B2(n_1083),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1119),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1147),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1088),
.B(n_1188),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1147),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1141),
.Y(n_1261)
);

INVx6_ASAP7_75t_L g1262 ( 
.A(n_1087),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_1143),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1165),
.A2(n_1099),
.B1(n_1083),
.B2(n_1151),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1151),
.A2(n_1077),
.B1(n_1203),
.B2(n_1178),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1077),
.B(n_1178),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1194),
.A2(n_1203),
.B1(n_1175),
.B2(n_1091),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1194),
.A2(n_1175),
.B1(n_1091),
.B2(n_1158),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_1081),
.Y(n_1269)
);

AO21x2_ASAP7_75t_L g1270 ( 
.A1(n_1157),
.A2(n_1108),
.B(n_1105),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1082),
.B(n_1185),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1082),
.A2(n_1096),
.B1(n_1185),
.B2(n_1150),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1144),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1188),
.B(n_1092),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1145),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1146),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1148),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_1131),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_1086),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1184),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1137),
.Y(n_1281)
);

NOR2x1_ASAP7_75t_L g1282 ( 
.A(n_1078),
.B(n_1187),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1142),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1188),
.B(n_1096),
.Y(n_1284)
);

BUFx12f_ASAP7_75t_L g1285 ( 
.A(n_1114),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1181),
.B(n_1114),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1155),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1152),
.A2(n_1156),
.B1(n_1094),
.B2(n_1104),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1152),
.Y(n_1289)
);

AO21x1_ASAP7_75t_SL g1290 ( 
.A1(n_1154),
.A2(n_1152),
.B(n_1094),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1078),
.A2(n_1187),
.B1(n_1162),
.B2(n_1174),
.Y(n_1291)
);

NAND2x1p5_ASAP7_75t_L g1292 ( 
.A(n_1104),
.B(n_1162),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1154),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1171),
.A2(n_904),
.B1(n_906),
.B2(n_897),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1089),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1087),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_SL g1297 ( 
.A1(n_1172),
.A2(n_906),
.B1(n_904),
.B2(n_897),
.Y(n_1297)
);

AOI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1173),
.A2(n_904),
.B1(n_906),
.B2(n_897),
.Y(n_1298)
);

NAND2x1p5_ASAP7_75t_L g1299 ( 
.A(n_1125),
.B(n_1132),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1079),
.A2(n_1048),
.B1(n_1061),
.B2(n_1053),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1171),
.A2(n_904),
.B1(n_906),
.B2(n_897),
.Y(n_1301)
);

INVxp33_ASAP7_75t_L g1302 ( 
.A(n_1189),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1089),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1287),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1218),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1226),
.B(n_1222),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_1213),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_SL g1308 ( 
.A1(n_1235),
.A2(n_1299),
.B(n_1233),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1234),
.B(n_1231),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1254),
.A2(n_1258),
.A3(n_1260),
.B(n_1283),
.Y(n_1310)
);

CKINVDCx11_ASAP7_75t_R g1311 ( 
.A(n_1213),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1226),
.B(n_1222),
.Y(n_1312)
);

AOI222xp33_ASAP7_75t_L g1313 ( 
.A1(n_1300),
.A2(n_1243),
.B1(n_1210),
.B2(n_1301),
.C1(n_1294),
.C2(n_1212),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1234),
.B(n_1231),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1253),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1297),
.A2(n_1298),
.B(n_1204),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1223),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1274),
.B(n_1248),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1274),
.B(n_1248),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1209),
.B(n_1284),
.Y(n_1320)
);

OR2x6_ASAP7_75t_L g1321 ( 
.A(n_1221),
.B(n_1299),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1289),
.B(n_1271),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1223),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1253),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1224),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1224),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1286),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1241),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1215),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_SL g1330 ( 
.A1(n_1208),
.A2(n_1228),
.B(n_1250),
.Y(n_1330)
);

INVx5_ASAP7_75t_SL g1331 ( 
.A(n_1221),
.Y(n_1331)
);

INVx5_ASAP7_75t_SL g1332 ( 
.A(n_1221),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1245),
.B(n_1259),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1241),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1289),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1271),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1245),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1271),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1221),
.B(n_1257),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1261),
.Y(n_1340)
);

OA21x2_ASAP7_75t_L g1341 ( 
.A1(n_1288),
.A2(n_1246),
.B(n_1247),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1242),
.B(n_1252),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1293),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1290),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1247),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1290),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1220),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1272),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1270),
.B(n_1251),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1225),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1229),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1292),
.A2(n_1291),
.B(n_1249),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1230),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1238),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1273),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1205),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1211),
.B(n_1232),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1303),
.B(n_1217),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1219),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1330),
.A2(n_1264),
.B1(n_1265),
.B2(n_1275),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1318),
.B(n_1295),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1306),
.B(n_1302),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1319),
.B(n_1255),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1327),
.B(n_1268),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1333),
.B(n_1280),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1344),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1306),
.B(n_1276),
.Y(n_1367)
);

AOI221xp5_ASAP7_75t_L g1368 ( 
.A1(n_1316),
.A2(n_1256),
.B1(n_1269),
.B2(n_1267),
.C(n_1278),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1341),
.Y(n_1369)
);

NAND2x1_ASAP7_75t_L g1370 ( 
.A(n_1308),
.B(n_1282),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1312),
.B(n_1277),
.Y(n_1371)
);

INVx1_ASAP7_75t_SL g1372 ( 
.A(n_1315),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1341),
.Y(n_1373)
);

INVxp67_ASAP7_75t_L g1374 ( 
.A(n_1315),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1322),
.B(n_1206),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1320),
.B(n_1296),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1357),
.A2(n_1263),
.B1(n_1279),
.B2(n_1227),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1341),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1341),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1310),
.B(n_1296),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1304),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1310),
.B(n_1296),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1310),
.B(n_1244),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1313),
.A2(n_1239),
.B1(n_1216),
.B2(n_1266),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1310),
.B(n_1244),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1324),
.Y(n_1386)
);

AND2x4_ASAP7_75t_SL g1387 ( 
.A(n_1346),
.B(n_1240),
.Y(n_1387)
);

NAND2x1_ASAP7_75t_L g1388 ( 
.A(n_1308),
.B(n_1262),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1362),
.B(n_1305),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1362),
.B(n_1323),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1384),
.A2(n_1348),
.B1(n_1321),
.B2(n_1342),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_SL g1392 ( 
.A1(n_1384),
.A2(n_1342),
.B(n_1348),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1362),
.B(n_1325),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1377),
.B(n_1329),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1377),
.B(n_1309),
.Y(n_1395)
);

NAND3xp33_ASAP7_75t_L g1396 ( 
.A(n_1368),
.B(n_1349),
.C(n_1355),
.Y(n_1396)
);

NAND3xp33_ASAP7_75t_L g1397 ( 
.A(n_1368),
.B(n_1340),
.C(n_1343),
.Y(n_1397)
);

OAI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1370),
.A2(n_1321),
.B1(n_1314),
.B2(n_1339),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1371),
.B(n_1326),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1376),
.B(n_1331),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1371),
.B(n_1334),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1371),
.B(n_1328),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1376),
.B(n_1331),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1376),
.B(n_1331),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_SL g1405 ( 
.A(n_1360),
.B(n_1364),
.Y(n_1405)
);

OAI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1360),
.A2(n_1336),
.B1(n_1338),
.B2(n_1339),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1367),
.B(n_1317),
.Y(n_1407)
);

NAND3xp33_ASAP7_75t_L g1408 ( 
.A(n_1364),
.B(n_1343),
.C(n_1317),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1367),
.B(n_1345),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1381),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1367),
.B(n_1311),
.Y(n_1411)
);

NAND3xp33_ASAP7_75t_L g1412 ( 
.A(n_1370),
.B(n_1335),
.C(n_1356),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1372),
.B(n_1347),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1361),
.B(n_1363),
.Y(n_1414)
);

AND2x2_ASAP7_75t_SL g1415 ( 
.A(n_1369),
.B(n_1346),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1388),
.A2(n_1352),
.B(n_1307),
.Y(n_1416)
);

AOI221xp5_ASAP7_75t_L g1417 ( 
.A1(n_1374),
.A2(n_1335),
.B1(n_1350),
.B2(n_1351),
.C(n_1353),
.Y(n_1417)
);

NAND3xp33_ASAP7_75t_L g1418 ( 
.A(n_1369),
.B(n_1354),
.C(n_1353),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1363),
.B(n_1374),
.Y(n_1419)
);

OAI21xp5_ASAP7_75t_SL g1420 ( 
.A1(n_1387),
.A2(n_1346),
.B(n_1337),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1388),
.A2(n_1337),
.B1(n_1332),
.B2(n_1331),
.Y(n_1421)
);

AOI221xp5_ASAP7_75t_L g1422 ( 
.A1(n_1373),
.A2(n_1379),
.B1(n_1378),
.B2(n_1351),
.C(n_1354),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1363),
.B(n_1350),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1381),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1375),
.B(n_1216),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1410),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1415),
.Y(n_1427)
);

NOR2x1_ASAP7_75t_L g1428 ( 
.A(n_1418),
.B(n_1366),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1410),
.Y(n_1429)
);

INVxp67_ASAP7_75t_SL g1430 ( 
.A(n_1418),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1424),
.Y(n_1431)
);

AOI221xp5_ASAP7_75t_L g1432 ( 
.A1(n_1396),
.A2(n_1379),
.B1(n_1378),
.B2(n_1373),
.C(n_1358),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1415),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1424),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1415),
.B(n_1380),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1422),
.B(n_1382),
.Y(n_1436)
);

NAND4xp25_ASAP7_75t_L g1437 ( 
.A(n_1396),
.B(n_1227),
.C(n_1359),
.D(n_1358),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1413),
.B(n_1383),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1423),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1409),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1407),
.Y(n_1441)
);

INVx4_ASAP7_75t_L g1442 ( 
.A(n_1400),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1403),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1403),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1419),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1414),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1404),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1389),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1416),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1390),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1421),
.B(n_1385),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1434),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1435),
.B(n_1421),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1431),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1426),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1448),
.B(n_1450),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1434),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1434),
.Y(n_1458)
);

INVxp67_ASAP7_75t_SL g1459 ( 
.A(n_1428),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1435),
.B(n_1411),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1448),
.B(n_1417),
.Y(n_1461)
);

OAI21xp33_ASAP7_75t_L g1462 ( 
.A1(n_1436),
.A2(n_1405),
.B(n_1392),
.Y(n_1462)
);

OAI21xp5_ASAP7_75t_SL g1463 ( 
.A1(n_1449),
.A2(n_1391),
.B(n_1397),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1427),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1435),
.B(n_1365),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1448),
.B(n_1450),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1450),
.B(n_1393),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1436),
.B(n_1402),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1436),
.B(n_1399),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1441),
.B(n_1401),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1438),
.B(n_1386),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1438),
.B(n_1386),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1426),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1428),
.B(n_1366),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1431),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1431),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1431),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1431),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1438),
.B(n_1408),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_SL g1480 ( 
.A(n_1449),
.B(n_1398),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1435),
.B(n_1365),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1431),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_1426),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1426),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1429),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1429),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1441),
.B(n_1408),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1429),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1441),
.B(n_1395),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1440),
.B(n_1430),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1452),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1453),
.B(n_1464),
.Y(n_1492)
);

NAND2x1p5_ASAP7_75t_L g1493 ( 
.A(n_1474),
.B(n_1428),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1452),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1479),
.B(n_1430),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1453),
.B(n_1427),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1483),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1457),
.Y(n_1498)
);

INVxp67_ASAP7_75t_SL g1499 ( 
.A(n_1459),
.Y(n_1499)
);

CKINVDCx20_ASAP7_75t_R g1500 ( 
.A(n_1460),
.Y(n_1500)
);

NAND2xp33_ASAP7_75t_SL g1501 ( 
.A(n_1460),
.B(n_1449),
.Y(n_1501)
);

NOR2x1p5_ASAP7_75t_L g1502 ( 
.A(n_1459),
.B(n_1437),
.Y(n_1502)
);

INVxp67_ASAP7_75t_SL g1503 ( 
.A(n_1487),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1457),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1458),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1458),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1464),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1465),
.B(n_1427),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1455),
.Y(n_1509)
);

AND3x2_ASAP7_75t_L g1510 ( 
.A(n_1474),
.B(n_1433),
.C(n_1394),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1479),
.B(n_1439),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1483),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1455),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1490),
.B(n_1439),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1474),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1483),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1488),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1486),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1462),
.B(n_1440),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1462),
.B(n_1440),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1488),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1465),
.B(n_1433),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1486),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1490),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1486),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1489),
.B(n_1445),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1489),
.B(n_1445),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1461),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1461),
.B(n_1445),
.Y(n_1529)
);

INVx2_ASAP7_75t_SL g1530 ( 
.A(n_1474),
.Y(n_1530)
);

INVxp33_ASAP7_75t_L g1531 ( 
.A(n_1463),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1469),
.B(n_1446),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1481),
.B(n_1433),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1528),
.B(n_1463),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1531),
.B(n_1469),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1500),
.B(n_1501),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1503),
.B(n_1487),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1491),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1491),
.Y(n_1539)
);

AOI221xp5_ASAP7_75t_L g1540 ( 
.A1(n_1519),
.A2(n_1480),
.B1(n_1432),
.B2(n_1437),
.C(n_1468),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1494),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1520),
.B(n_1468),
.Y(n_1542)
);

INVx2_ASAP7_75t_SL g1543 ( 
.A(n_1515),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1502),
.A2(n_1442),
.B1(n_1397),
.B2(n_1432),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1496),
.B(n_1481),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1494),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1496),
.B(n_1442),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1495),
.B(n_1456),
.Y(n_1548)
);

CKINVDCx16_ASAP7_75t_R g1549 ( 
.A(n_1492),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1492),
.B(n_1442),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1529),
.B(n_1467),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1526),
.B(n_1442),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1508),
.B(n_1442),
.Y(n_1553)
);

INVx1_ASAP7_75t_SL g1554 ( 
.A(n_1510),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1515),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1508),
.B(n_1442),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1522),
.B(n_1451),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1527),
.B(n_1425),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1495),
.B(n_1207),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1512),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1522),
.B(n_1451),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1533),
.B(n_1451),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1498),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1498),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1532),
.B(n_1456),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1504),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_1507),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1524),
.B(n_1467),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1511),
.B(n_1466),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1541),
.Y(n_1570)
);

AOI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1536),
.A2(n_1499),
.B(n_1493),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1534),
.A2(n_1502),
.B1(n_1530),
.B2(n_1432),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1541),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1549),
.B(n_1533),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1559),
.B(n_1207),
.Y(n_1575)
);

INVxp67_ASAP7_75t_L g1576 ( 
.A(n_1535),
.Y(n_1576)
);

NAND4xp25_ASAP7_75t_L g1577 ( 
.A(n_1554),
.B(n_1437),
.C(n_1513),
.D(n_1509),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1546),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1544),
.A2(n_1493),
.B1(n_1420),
.B2(n_1530),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1567),
.B(n_1466),
.Y(n_1580)
);

OAI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1540),
.A2(n_1493),
.B(n_1514),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1546),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1543),
.B(n_1504),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1545),
.B(n_1443),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1552),
.A2(n_1451),
.B1(n_1406),
.B2(n_1398),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1537),
.B(n_1511),
.Y(n_1586)
);

OR2x6_ASAP7_75t_L g1587 ( 
.A(n_1543),
.B(n_1285),
.Y(n_1587)
);

OAI322xp33_ASAP7_75t_L g1588 ( 
.A1(n_1542),
.A2(n_1514),
.A3(n_1513),
.B1(n_1521),
.B2(n_1517),
.C1(n_1509),
.C2(n_1505),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1563),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1558),
.B(n_1470),
.Y(n_1590)
);

OAI321xp33_ASAP7_75t_L g1591 ( 
.A1(n_1555),
.A2(n_1521),
.A3(n_1517),
.B1(n_1512),
.B2(n_1525),
.C(n_1523),
.Y(n_1591)
);

INVxp67_ASAP7_75t_L g1592 ( 
.A(n_1555),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1545),
.B(n_1470),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1551),
.B(n_1471),
.Y(n_1594)
);

O2A1O1Ixp33_ASAP7_75t_L g1595 ( 
.A1(n_1568),
.A2(n_1506),
.B(n_1505),
.C(n_1512),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1592),
.B(n_1557),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1574),
.B(n_1557),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1587),
.B(n_1547),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1586),
.B(n_1548),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1587),
.B(n_1547),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1576),
.B(n_1548),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1587),
.B(n_1550),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1583),
.B(n_1550),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1570),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1573),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1578),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1582),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1590),
.B(n_1557),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1575),
.B(n_1556),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1572),
.A2(n_1556),
.B1(n_1562),
.B2(n_1561),
.Y(n_1610)
);

NAND2x1p5_ASAP7_75t_L g1611 ( 
.A(n_1583),
.B(n_1571),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1589),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1580),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1581),
.B(n_1561),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1604),
.Y(n_1615)
);

NAND4xp75_ASAP7_75t_L g1616 ( 
.A(n_1614),
.B(n_1591),
.C(n_1588),
.D(n_1553),
.Y(n_1616)
);

NOR3x1_ASAP7_75t_L g1617 ( 
.A(n_1596),
.B(n_1577),
.C(n_1579),
.Y(n_1617)
);

AOI221xp5_ASAP7_75t_L g1618 ( 
.A1(n_1610),
.A2(n_1591),
.B1(n_1595),
.B2(n_1577),
.C(n_1585),
.Y(n_1618)
);

AOI221xp5_ASAP7_75t_L g1619 ( 
.A1(n_1601),
.A2(n_1593),
.B1(n_1566),
.B2(n_1563),
.C(n_1564),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1601),
.B(n_1562),
.Y(n_1620)
);

NOR3xp33_ASAP7_75t_SL g1621 ( 
.A(n_1609),
.B(n_1214),
.C(n_1564),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1603),
.B(n_1594),
.Y(n_1622)
);

NOR3x1_ASAP7_75t_L g1623 ( 
.A(n_1597),
.B(n_1613),
.C(n_1608),
.Y(n_1623)
);

O2A1O1Ixp33_ASAP7_75t_L g1624 ( 
.A1(n_1611),
.A2(n_1538),
.B(n_1539),
.C(n_1566),
.Y(n_1624)
);

NAND3xp33_ASAP7_75t_SL g1625 ( 
.A(n_1611),
.B(n_1263),
.C(n_1279),
.Y(n_1625)
);

NOR3xp33_ASAP7_75t_L g1626 ( 
.A(n_1625),
.B(n_1609),
.C(n_1606),
.Y(n_1626)
);

AO22x2_ASAP7_75t_L g1627 ( 
.A1(n_1616),
.A2(n_1612),
.B1(n_1605),
.B2(n_1607),
.Y(n_1627)
);

NOR3xp33_ASAP7_75t_L g1628 ( 
.A(n_1618),
.B(n_1602),
.C(n_1599),
.Y(n_1628)
);

AOI21xp33_ASAP7_75t_L g1629 ( 
.A1(n_1624),
.A2(n_1600),
.B(n_1598),
.Y(n_1629)
);

AND4x1_ASAP7_75t_L g1630 ( 
.A(n_1623),
.B(n_1617),
.C(n_1621),
.D(n_1622),
.Y(n_1630)
);

AOI211xp5_ASAP7_75t_L g1631 ( 
.A1(n_1619),
.A2(n_1600),
.B(n_1598),
.C(n_1603),
.Y(n_1631)
);

NOR3xp33_ASAP7_75t_L g1632 ( 
.A(n_1620),
.B(n_1239),
.C(n_1214),
.Y(n_1632)
);

NOR3xp33_ASAP7_75t_L g1633 ( 
.A(n_1615),
.B(n_1560),
.C(n_1584),
.Y(n_1633)
);

OA22x2_ASAP7_75t_SL g1634 ( 
.A1(n_1616),
.A2(n_1560),
.B1(n_1516),
.B2(n_1497),
.Y(n_1634)
);

NOR3x1_ASAP7_75t_L g1635 ( 
.A(n_1625),
.B(n_1565),
.C(n_1569),
.Y(n_1635)
);

NOR3x1_ASAP7_75t_L g1636 ( 
.A(n_1625),
.B(n_1565),
.C(n_1569),
.Y(n_1636)
);

OAI211xp5_ASAP7_75t_SL g1637 ( 
.A1(n_1629),
.A2(n_1523),
.B(n_1525),
.C(n_1518),
.Y(n_1637)
);

AOI221xp5_ASAP7_75t_L g1638 ( 
.A1(n_1627),
.A2(n_1556),
.B1(n_1553),
.B2(n_1518),
.C(n_1516),
.Y(n_1638)
);

AOI221xp5_ASAP7_75t_L g1639 ( 
.A1(n_1628),
.A2(n_1518),
.B1(n_1497),
.B2(n_1506),
.C(n_1412),
.Y(n_1639)
);

NAND3xp33_ASAP7_75t_L g1640 ( 
.A(n_1630),
.B(n_1281),
.C(n_1236),
.Y(n_1640)
);

OAI211xp5_ASAP7_75t_SL g1641 ( 
.A1(n_1631),
.A2(n_1443),
.B(n_1472),
.C(n_1471),
.Y(n_1641)
);

OR3x1_ASAP7_75t_L g1642 ( 
.A(n_1634),
.B(n_1636),
.C(n_1635),
.Y(n_1642)
);

OR2x6_ASAP7_75t_L g1643 ( 
.A(n_1640),
.B(n_1237),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1642),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1637),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1641),
.B(n_1633),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_SL g1647 ( 
.A(n_1638),
.B(n_1626),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1639),
.Y(n_1648)
);

NAND4xp75_ASAP7_75t_L g1649 ( 
.A(n_1644),
.B(n_1632),
.C(n_1240),
.D(n_1236),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1646),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1643),
.B(n_1443),
.Y(n_1651)
);

CKINVDCx16_ASAP7_75t_R g1652 ( 
.A(n_1643),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_1647),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1650),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1652),
.B(n_1645),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1653),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1656),
.Y(n_1657)
);

AOI311xp33_ASAP7_75t_L g1658 ( 
.A1(n_1657),
.A2(n_1655),
.A3(n_1648),
.B(n_1653),
.C(n_1654),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1658),
.A2(n_1651),
.B(n_1649),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1658),
.B(n_1454),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1659),
.A2(n_1285),
.B1(n_1475),
.B2(n_1476),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1660),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_SL g1663 ( 
.A(n_1661),
.B(n_1454),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1662),
.B(n_1472),
.Y(n_1664)
);

OAI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1664),
.A2(n_1447),
.B(n_1444),
.Y(n_1665)
);

AOI322xp5_ASAP7_75t_L g1666 ( 
.A1(n_1665),
.A2(n_1663),
.A3(n_1478),
.B1(n_1477),
.B2(n_1475),
.C1(n_1482),
.C2(n_1476),
.Y(n_1666)
);

AOI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1666),
.A2(n_1454),
.B1(n_1475),
.B2(n_1476),
.C(n_1482),
.Y(n_1667)
);

AOI211xp5_ASAP7_75t_L g1668 ( 
.A1(n_1667),
.A2(n_1485),
.B(n_1484),
.C(n_1473),
.Y(n_1668)
);


endmodule