module fake_jpeg_12374_n_188 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_188);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_15),
.B(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_5),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_31),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_22),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_26),
.C(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_25),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_9),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_6),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_10),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_11),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_57),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_32),
.B1(n_30),
.B2(n_33),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_53),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_48),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_28),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_65),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_32),
.B1(n_18),
.B2(n_29),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_27),
.B1(n_30),
.B2(n_24),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_21),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_26),
.B1(n_29),
.B2(n_27),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_66),
.A2(n_48),
.B1(n_2),
.B2(n_3),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_18),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_74),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_37),
.B(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_37),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_28),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_92),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_29),
.B1(n_37),
.B2(n_48),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_70),
.B1(n_52),
.B2(n_54),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_94),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_24),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_83),
.B(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_14),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_1),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_95),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_88),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_13),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_89),
.B(n_93),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_73),
.B1(n_55),
.B2(n_68),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_12),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_1),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_58),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_101),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_2),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_97),
.B(n_99),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_54),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_4),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_4),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_114),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_70),
.B(n_72),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_106),
.A2(n_117),
.B(n_79),
.Y(n_134)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_81),
.B(n_12),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_111),
.B(n_78),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_116),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_86),
.A2(n_5),
.B1(n_55),
.B2(n_92),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_120),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_L g120 ( 
.A1(n_76),
.A2(n_87),
.B(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_130),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_95),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_102),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_83),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_126),
.C(n_103),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_99),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_117),
.A2(n_78),
.B1(n_77),
.B2(n_98),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_129),
.A2(n_103),
.B1(n_114),
.B2(n_106),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_115),
.B(n_96),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_138),
.B1(n_119),
.B2(n_110),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_121),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_137),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_105),
.B(n_101),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_103),
.A2(n_77),
.B1(n_98),
.B2(n_100),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_145),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_143),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g143 ( 
.A1(n_136),
.A2(n_112),
.A3(n_114),
.B1(n_111),
.B2(n_98),
.C1(n_77),
.C2(n_104),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_132),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_108),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_150),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_132),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_148),
.Y(n_157)
);

AND2x4_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_151),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_88),
.C(n_109),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_133),
.C(n_138),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_148),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_129),
.C(n_133),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_159),
.C(n_163),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_133),
.C(n_131),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_118),
.C(n_127),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_144),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_152),
.B(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_168),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_139),
.C(n_146),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_164),
.C(n_158),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_145),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_171),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_164),
.Y(n_174)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_165),
.A2(n_162),
.B1(n_157),
.B2(n_119),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_167),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_174),
.B(n_175),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_172),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_173),
.B(n_174),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_180),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_176),
.B(n_175),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_177),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_183),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_178),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_185),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_184),
.Y(n_187)
);

BUFx24_ASAP7_75t_SL g188 ( 
.A(n_187),
.Y(n_188)
);


endmodule