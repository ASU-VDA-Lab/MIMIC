module real_jpeg_15090_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_331, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_331;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_3),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_3),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_56),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_56),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_4),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_4),
.A2(n_39),
.B1(n_58),
.B2(n_59),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_4),
.A2(n_39),
.B1(n_53),
.B2(n_54),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_254)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_6),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_6),
.A2(n_35),
.B1(n_58),
.B2(n_59),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_6),
.A2(n_35),
.B1(n_53),
.B2(n_54),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_7),
.A2(n_40),
.B1(n_41),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_7),
.A2(n_49),
.B1(n_58),
.B2(n_59),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_49),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_7),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_8),
.A2(n_53),
.B1(n_54),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_8),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_68),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_68),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_68),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_9),
.A2(n_58),
.B1(n_59),
.B2(n_79),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_9),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_9),
.A2(n_53),
.B1(n_54),
.B2(n_79),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_9),
.A2(n_40),
.B1(n_41),
.B2(n_79),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_79),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_10),
.A2(n_53),
.B1(n_54),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_10),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_121),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_121),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_121),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_12),
.A2(n_40),
.B1(n_41),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_12),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_161),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_12),
.A2(n_58),
.B1(n_59),
.B2(n_161),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_12),
.A2(n_53),
.B1(n_54),
.B2(n_161),
.Y(n_264)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_13),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_149),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_14),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_14),
.B(n_30),
.C(n_44),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_14),
.B(n_77),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_14),
.A2(n_112),
.B(n_165),
.Y(n_181)
);

O2A1O1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_14),
.A2(n_58),
.B(n_76),
.C(n_192),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_149),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_14),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_14),
.B(n_53),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_15),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_57)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_15),
.A2(n_53),
.B1(n_54),
.B2(n_61),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g250 ( 
.A(n_15),
.B(n_59),
.Y(n_250)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_322),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_309),
.B(n_321),
.Y(n_18)
);

AO21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_137),
.B(n_306),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_124),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_99),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_22),
.B(n_99),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_69),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_23),
.B(n_70),
.C(n_85),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.B(n_51),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_24),
.A2(n_25),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_36),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_26),
.A2(n_27),
.B1(n_51),
.B2(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_26),
.A2(n_27),
.B1(n_36),
.B2(n_37),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_32),
.B(n_33),
.Y(n_27)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_28),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_28),
.A2(n_32),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_28),
.B(n_166),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_28),
.A2(n_32),
.B1(n_111),
.B2(n_254),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_30),
.B1(n_44),
.B2(n_45),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_29),
.B(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_32),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_32),
.B(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_34),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B1(n_47),
.B2(n_50),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_38),
.A2(n_42),
.B1(n_50),
.B2(n_116),
.Y(n_115)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

AO22x1_ASAP7_75t_SL g77 ( 
.A1(n_40),
.A2(n_41),
.B1(n_75),
.B2(n_76),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_40),
.B(n_153),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_41),
.A2(n_75),
.B(n_149),
.Y(n_192)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_42),
.A2(n_50),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_42),
.B(n_151),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_42),
.A2(n_50),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_42),
.A2(n_50),
.B1(n_116),
.B2(n_243),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_46),
.A2(n_48),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_46),
.A2(n_160),
.B(n_162),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_46),
.B(n_149),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_46),
.A2(n_162),
.B(n_242),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_50),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_57),
.B(n_62),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_57),
.B1(n_64),
.B2(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_54),
.A2(n_64),
.B(n_149),
.C(n_236),
.Y(n_235)
);

AOI32xp33_ASAP7_75t_L g249 ( 
.A1(n_54),
.A2(n_58),
.A3(n_61),
.B1(n_237),
.B2(n_250),
.Y(n_249)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_57),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_57),
.B(n_67),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_57),
.A2(n_64),
.B1(n_88),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_57),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_57),
.A2(n_62),
.B(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_57),
.A2(n_64),
.B1(n_120),
.B2(n_264),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_59),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_63),
.A2(n_217),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_63),
.A2(n_217),
.B1(n_316),
.B2(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_64),
.A2(n_120),
.B(n_122),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_85),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_71),
.B(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_82),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_72),
.A2(n_78),
.B1(n_80),
.B2(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_72),
.A2(n_80),
.B1(n_93),
.B2(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_72),
.A2(n_197),
.B(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_72),
.A2(n_80),
.B1(n_212),
.B2(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_72),
.A2(n_198),
.B(n_240),
.Y(n_262)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_77),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_73),
.B(n_199),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_73),
.A2(n_77),
.B(n_313),
.Y(n_312)
);

NOR2x1_ASAP7_75t_R g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_77),
.B(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_80),
.A2(n_212),
.B(n_213),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_80),
.A2(n_118),
.B(n_213),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_83),
.A2(n_148),
.B(n_150),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_83),
.A2(n_150),
.B(n_225),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_98),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_86),
.A2(n_87),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_SL g135 ( 
.A(n_87),
.B(n_90),
.C(n_95),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_87),
.B(n_128),
.C(n_135),
.Y(n_320)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_94),
.A2(n_95),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_95),
.B(n_129),
.C(n_133),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_105),
.C(n_106),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_100),
.A2(n_101),
.B1(n_105),
.B2(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_105),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_106),
.B(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_117),
.C(n_119),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_107),
.A2(n_108),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_114),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_109),
.A2(n_114),
.B1(n_115),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_109),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_112),
.A2(n_164),
.B(n_165),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_112),
.A2(n_113),
.B1(n_194),
.B2(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_112),
.A2(n_113),
.B1(n_220),
.B2(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_113),
.A2(n_171),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_113),
.B(n_149),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_113),
.A2(n_179),
.B(n_194),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_117),
.B(n_119),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_123),
.B(n_235),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_L g306 ( 
.A1(n_124),
.A2(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_136),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_125),
.B(n_136),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_135),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_130),
.Y(n_315)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_134),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_300),
.B(n_305),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_288),
.B(n_299),
.Y(n_138)
);

OAI321xp33_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_256),
.A3(n_281),
.B1(n_286),
.B2(n_287),
.C(n_331),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_229),
.B(n_255),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_206),
.B(n_228),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_187),
.B(n_205),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_167),
.B(n_186),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_154),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_145),
.B(n_154),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_152),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_147),
.B1(n_152),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_152),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_163),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_159),
.C(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_164),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_175),
.B(n_185),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_169),
.B(n_173),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_180),
.B(n_184),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_177),
.B(n_178),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_188),
.B(n_189),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_195),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_200),
.C(n_204),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_193),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_200),
.B1(n_203),
.B2(n_204),
.Y(n_195)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_200),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_202),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_207),
.B(n_208),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_221),
.B2(n_222),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_224),
.C(n_226),
.Y(n_230)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_215),
.C(n_219),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_226),
.B2(n_227),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_223),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_230),
.B(n_231),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_245),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_232),
.B(n_246),
.C(n_247),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_238),
.B2(n_244),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_233),
.B(n_239),
.C(n_241),
.Y(n_270)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_238),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_251),
.B2(n_252),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_252),
.Y(n_266)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_271),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_271),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_267),
.C(n_270),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_258),
.A2(n_259),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_266),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_265),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_265),
.C(n_266),
.Y(n_280)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_263),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_267),
.B(n_270),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_269),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_280),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_275),
.C(n_280),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_279),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_278),
.C(n_279),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_282),
.B(n_283),
.Y(n_286)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_298),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_298),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_293),
.C(n_294),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_302),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_320),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_320),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_319),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_314),
.B1(n_317),
.B2(n_318),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_312),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_314),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_317),
.C(n_319),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_327),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_326),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_324),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_326),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);


endmodule