module fake_jpeg_25473_n_275 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_275);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_275;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_6),
.B(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_38),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_20),
.B1(n_25),
.B2(n_15),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_25),
.B1(n_20),
.B2(n_19),
.Y(n_56)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_20),
.B1(n_15),
.B2(n_25),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_26),
.B1(n_18),
.B2(n_29),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_16),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_47),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_21),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_50),
.B(n_45),
.C(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_23),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_21),
.Y(n_50)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_53),
.B(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_22),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_64),
.B1(n_80),
.B2(n_50),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_54),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_58),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_47),
.Y(n_58)
);

INVxp67_ASAP7_75t_SL g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_70),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_22),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_60),
.B(n_73),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_29),
.B1(n_24),
.B2(n_19),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_61),
.A2(n_65),
.B1(n_48),
.B2(n_51),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_50),
.B1(n_44),
.B2(n_18),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_63),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_39),
.A2(n_29),
.B1(n_28),
.B2(n_26),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_50),
.B(n_41),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_51),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_40),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_72),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_28),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_76),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_39),
.A2(n_30),
.B1(n_27),
.B2(n_3),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_78),
.B1(n_48),
.B2(n_43),
.Y(n_85)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_38),
.C(n_23),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_48),
.C(n_52),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_43),
.A2(n_30),
.B1(n_27),
.B2(n_3),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_42),
.A2(n_23),
.B1(n_28),
.B2(n_1),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_83),
.B(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_85),
.A2(n_92),
.B1(n_97),
.B2(n_79),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_72),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_86),
.B(n_87),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_51),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_94),
.Y(n_124)
);

AO21x2_ASAP7_75t_L g97 ( 
.A1(n_59),
.A2(n_48),
.B(n_49),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_105),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_63),
.B(n_71),
.Y(n_111)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_77),
.C(n_74),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_76),
.A2(n_52),
.B1(n_2),
.B2(n_1),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_104),
.A2(n_62),
.B1(n_81),
.B2(n_58),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_10),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_68),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_106),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_55),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_116),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_111),
.A2(n_88),
.B(n_90),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_112),
.A2(n_82),
.B1(n_52),
.B2(n_84),
.Y(n_162)
);

BUFx24_ASAP7_75t_SL g113 ( 
.A(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_119),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_55),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_103),
.C(n_88),
.Y(n_153)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_118),
.B(n_121),
.Y(n_143)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_89),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_89),
.B(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_123),
.Y(n_142)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_63),
.C(n_5),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_128),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_91),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_127),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_106),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_95),
.B(n_73),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_133),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_66),
.Y(n_131)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

AND2x6_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_88),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_136),
.B(n_140),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_129),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_108),
.Y(n_141)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_101),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_155),
.Y(n_163)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_147),
.Y(n_169)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_97),
.B(n_90),
.C(n_83),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_149),
.A2(n_151),
.B(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_160),
.Y(n_167)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_112),
.C(n_124),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_107),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_82),
.B(n_92),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_110),
.B(n_96),
.Y(n_157)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

MAJx2_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_116),
.C(n_122),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_7),
.Y(n_185)
);

AOI22x1_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_104),
.B1(n_80),
.B2(n_56),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_182)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_114),
.B(n_102),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_161),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_114),
.B1(n_119),
.B2(n_81),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_139),
.A2(n_133),
.B1(n_123),
.B2(n_125),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_149),
.B1(n_154),
.B2(n_145),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_SL g192 ( 
.A(n_166),
.B(n_174),
.C(n_176),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_128),
.Y(n_170)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_127),
.Y(n_171)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_132),
.C(n_115),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_179),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_99),
.B1(n_81),
.B2(n_66),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_99),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_155),
.Y(n_206)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_138),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_180),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_187),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_159),
.A2(n_14),
.B1(n_7),
.B2(n_8),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_159),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_185),
.B(n_137),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_144),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_186),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_143),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_160),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_193),
.B1(n_200),
.B2(n_208),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_145),
.B1(n_150),
.B2(n_156),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_199),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_195),
.B(n_197),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_185),
.B(n_135),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_169),
.A2(n_147),
.B1(n_152),
.B2(n_162),
.Y(n_200)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_167),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_209),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_167),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_189),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_166),
.C(n_175),
.Y(n_215)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_172),
.A2(n_136),
.B1(n_158),
.B2(n_151),
.Y(n_208)
);

INVxp67_ASAP7_75t_SL g209 ( 
.A(n_168),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_163),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_211),
.C(n_215),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_163),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_171),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_217),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_170),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_218),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_179),
.B1(n_188),
.B2(n_182),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_221),
.A2(n_225),
.B1(n_193),
.B2(n_190),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_188),
.B(n_181),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_223),
.Y(n_236)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_184),
.B1(n_173),
.B2(n_178),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_228),
.A2(n_232),
.B1(n_238),
.B2(n_224),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_196),
.B1(n_206),
.B2(n_199),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_229),
.A2(n_213),
.B1(n_212),
.B2(n_12),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_214),
.B(n_204),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_230),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_203),
.B(n_165),
.Y(n_231)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_221),
.A2(n_206),
.B1(n_187),
.B2(n_177),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_194),
.C(n_177),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_211),
.C(n_216),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_225),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_235),
.Y(n_239)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_210),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_246),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_241),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_243),
.C(n_248),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_218),
.C(n_217),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_245),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_236),
.A2(n_229),
.B(n_227),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_237),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_12),
.C(n_13),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_239),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_253),
.B(n_254),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_228),
.C(n_232),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_247),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_255),
.B(n_249),
.Y(n_259)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_244),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_238),
.C(n_245),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_253),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_254),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_248),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_263),
.C(n_264),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_240),
.C(n_241),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_266),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_267),
.B(n_258),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_268),
.A2(n_258),
.B(n_251),
.Y(n_269)
);

AOI31xp33_ASAP7_75t_L g272 ( 
.A1(n_269),
.A2(n_270),
.A3(n_265),
.B(n_235),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_272),
.A2(n_271),
.B(n_227),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_233),
.C(n_13),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_233),
.Y(n_275)
);


endmodule