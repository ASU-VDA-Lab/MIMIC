module real_jpeg_6655_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_286;
wire n_221;
wire n_176;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_148;
wire n_19;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_213;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_1),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_1),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_2),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_2),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_2),
.A2(n_39),
.B1(n_67),
.B2(n_69),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_2),
.A2(n_39),
.B1(n_97),
.B2(n_99),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_2),
.A2(n_39),
.B1(n_141),
.B2(n_143),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_2),
.B(n_69),
.C(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_2),
.B(n_200),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_2),
.A2(n_207),
.B(n_209),
.C(n_210),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_2),
.B(n_221),
.C(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_2),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_2),
.B(n_162),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_2),
.B(n_18),
.Y(n_247)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_4),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_4),
.Y(n_234)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_5),
.Y(n_188)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_7),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_7),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_7),
.A2(n_58),
.B1(n_82),
.B2(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_8),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_9),
.A2(n_84),
.B1(n_92),
.B2(n_94),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_9),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_9),
.A2(n_94),
.B1(n_133),
.B2(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_10),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_10),
.Y(n_111)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_10),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_172),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_171),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_151),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_14),
.B(n_151),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_122),
.C(n_136),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_15),
.B(n_122),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_70),
.B1(n_120),
.B2(n_121),
.Y(n_15)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_16),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_16),
.B(n_137),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_16),
.A2(n_120),
.B1(n_181),
.B2(n_270),
.Y(n_269)
);

XNOR2x1_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_41),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_17),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_17),
.B(n_148),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_17),
.A2(n_123),
.B1(n_124),
.B2(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_17),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_17),
.A2(n_169),
.B1(n_203),
.B2(n_214),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_17),
.B(n_95),
.Y(n_277)
);

OA21x2_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_28),
.B(n_37),
.Y(n_17)
);

NOR2x1_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_29),
.Y(n_28)
);

AO22x1_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_21),
.B1(n_25),
.B2(n_26),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_24),
.Y(n_212)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_29)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_39),
.A2(n_55),
.B(n_58),
.Y(n_209)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_41),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_41),
.B(n_157),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_41),
.A2(n_150),
.B(n_169),
.C(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_41),
.A2(n_95),
.B1(n_148),
.B2(n_178),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_41),
.A2(n_148),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

AO21x2_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_54),
.B(n_66),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_54),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_43)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_44),
.Y(n_208)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_54),
.Y(n_200)
);

OA22x2_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_57),
.B1(n_60),
.B2(n_63),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_70),
.A2(n_147),
.B(n_149),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_95),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_71),
.A2(n_95),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_71),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_78),
.B1(n_87),
.B2(n_91),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_76),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_72),
.A2(n_78),
.B1(n_139),
.B2(n_145),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_74),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_91),
.B(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_95),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_95),
.B(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_95),
.A2(n_178),
.B1(n_199),
.B2(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_95),
.A2(n_178),
.B1(n_218),
.B2(n_219),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_95),
.A2(n_178),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

O2A1O1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_95),
.A2(n_148),
.B(n_205),
.C(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_95),
.B(n_148),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_95),
.A2(n_138),
.B1(n_178),
.B2(n_274),
.Y(n_273)
);

AND2x4_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g223 ( 
.A(n_98),
.Y(n_223)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_112),
.Y(n_102)
);

NAND2x1_ASAP7_75t_SL g112 ( 
.A(n_103),
.B(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_112),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_106),
.B1(n_108),
.B2(n_111),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_104),
.B(n_231),
.Y(n_230)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_117),
.B2(n_119),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_116),
.Y(n_222)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_135),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_127),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_126),
.B(n_140),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_130),
.A2(n_158),
.B1(n_159),
.B2(n_162),
.Y(n_157)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_136),
.B(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_147),
.B(n_149),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_138),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_156),
.B(n_163),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_148),
.B(n_189),
.C(n_246),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AND3x1_ASAP7_75t_L g276 ( 
.A(n_150),
.B(n_253),
.C(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_170),
.Y(n_151)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_164),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_192),
.B(n_286),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_190),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_175),
.B(n_190),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.C(n_180),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_176),
.B(n_177),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_199),
.C(n_201),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_178),
.B(n_243),
.C(n_250),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_180),
.B(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_181),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_189),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_182),
.A2(n_183),
.B1(n_189),
.B2(n_201),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_189),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_189),
.A2(n_201),
.B1(n_206),
.B2(n_213),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_189),
.B(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_189),
.A2(n_201),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_189),
.B(n_206),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_265),
.B(n_283),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_255),
.B(n_264),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_241),
.B(n_254),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_215),
.B(n_240),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_202),
.Y(n_240)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_201),
.B(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_201),
.B(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_214),
.Y(n_202)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_203),
.Y(n_214)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_227),
.B(n_239),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_224),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_224),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_237),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_235),
.Y(n_228)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_251),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_251),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_248),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_257),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_261),
.C(n_262),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NOR2x1_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_278),
.Y(n_265)
);

NOR2x1_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_268),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_275),
.B2(n_276),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_275),
.C(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_278),
.A2(n_284),
.B(n_285),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_281),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);


endmodule