module real_aes_17730_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_867;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_617;
wire n_402;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_855;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AND2x4_ASAP7_75t_L g121 ( .A(n_0), .B(n_122), .Y(n_121) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_1), .A2(n_34), .B1(n_149), .B2(n_241), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_2), .A2(n_10), .B1(n_546), .B2(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g122 ( .A(n_3), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_4), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_5), .A2(n_11), .B1(n_547), .B2(n_583), .Y(n_582) );
XNOR2xp5_ASAP7_75t_L g832 ( .A(n_6), .B(n_833), .Y(n_832) );
BUFx2_ASAP7_75t_L g113 ( .A(n_7), .Y(n_113) );
OR2x2_ASAP7_75t_L g842 ( .A(n_7), .B(n_30), .Y(n_842) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_8), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_9), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_12), .B(n_164), .Y(n_163) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_13), .A2(n_101), .B1(n_194), .B2(n_546), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_14), .A2(n_31), .B1(n_564), .B2(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_15), .B(n_164), .Y(n_561) );
OAI21x1_ASAP7_75t_L g144 ( .A1(n_16), .A2(n_47), .B(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_17), .B(n_245), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_18), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_19), .A2(n_38), .B1(n_201), .B2(n_216), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_20), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_21), .A2(n_44), .B1(n_216), .B2(n_546), .Y(n_602) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_22), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_23), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_24), .B(n_224), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_25), .Y(n_553) );
XNOR2x1_ASAP7_75t_L g833 ( .A(n_26), .B(n_39), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_27), .B(n_142), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_28), .Y(n_873) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_29), .Y(n_193) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_30), .Y(n_111) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_32), .A2(n_84), .B1(n_149), .B2(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_33), .A2(n_37), .B1(n_149), .B2(n_549), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_35), .A2(n_50), .B1(n_546), .B2(n_601), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_36), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_40), .B(n_164), .Y(n_212) );
INVx2_ASAP7_75t_L g837 ( .A(n_41), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_42), .B(n_197), .Y(n_239) );
INVx1_ASAP7_75t_L g116 ( .A(n_43), .Y(n_116) );
BUFx3_ASAP7_75t_L g840 ( .A(n_43), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_45), .B(n_183), .Y(n_247) );
XOR2x2_ASAP7_75t_L g131 ( .A(n_46), .B(n_132), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g855 ( .A1(n_46), .A2(n_856), .B1(n_857), .B2(n_860), .Y(n_855) );
INVx1_ASAP7_75t_L g860 ( .A(n_46), .Y(n_860) );
AND2x2_ASAP7_75t_L g275 ( .A(n_48), .B(n_183), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_49), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_51), .B(n_224), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_52), .B(n_201), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_53), .A2(n_70), .B1(n_201), .B2(n_601), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_54), .A2(n_73), .B1(n_149), .B2(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_55), .B(n_305), .Y(n_304) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_56), .A2(n_153), .B(n_162), .C(n_268), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_57), .A2(n_98), .B1(n_546), .B2(n_547), .Y(n_545) );
INVx1_ASAP7_75t_L g145 ( .A(n_58), .Y(n_145) );
AND2x4_ASAP7_75t_L g167 ( .A(n_59), .B(n_168), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_60), .A2(n_61), .B1(n_216), .B2(n_228), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g857 ( .A1(n_62), .A2(n_81), .B1(n_858), .B2(n_859), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_62), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_63), .B(n_142), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_64), .B(n_183), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_65), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_66), .B(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g168 ( .A(n_67), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_68), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_69), .B(n_142), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_71), .B(n_149), .Y(n_300) );
NAND3xp33_ASAP7_75t_L g240 ( .A(n_72), .B(n_197), .C(n_241), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g870 ( .A(n_74), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_75), .B(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g155 ( .A(n_76), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_77), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_78), .B(n_164), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_79), .B(n_158), .Y(n_157) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_80), .A2(n_97), .B1(n_162), .B2(n_216), .Y(n_533) );
INVx1_ASAP7_75t_L g859 ( .A(n_81), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_82), .Y(n_604) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_83), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_85), .A2(n_91), .B1(n_223), .B2(n_224), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_86), .B(n_164), .Y(n_196) );
NAND2xp33_ASAP7_75t_SL g181 ( .A(n_87), .B(n_152), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_88), .B(n_195), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g881 ( .A(n_89), .Y(n_881) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_90), .B(n_142), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_92), .Y(n_586) );
INVx1_ASAP7_75t_L g120 ( .A(n_93), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g866 ( .A(n_93), .B(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g845 ( .A(n_94), .Y(n_845) );
NAND2xp33_ASAP7_75t_L g565 ( .A(n_95), .B(n_164), .Y(n_565) );
NAND2xp33_ASAP7_75t_L g151 ( .A(n_96), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_99), .B(n_183), .Y(n_307) );
NAND3xp33_ASAP7_75t_L g177 ( .A(n_100), .B(n_152), .C(n_176), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_102), .B(n_149), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_103), .B(n_224), .Y(n_303) );
AOI21xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_123), .B(n_880), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx6p67_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx12_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx5_ASAP7_75t_L g882 ( .A(n_108), .Y(n_882) );
OR2x6_ASAP7_75t_L g108 ( .A(n_109), .B(n_114), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NOR2x1p5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_117), .Y(n_114) );
AND3x2_ASAP7_75t_L g852 ( .A(n_115), .B(n_119), .C(n_841), .Y(n_852) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g867 ( .A(n_116), .Y(n_867) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g130 ( .A(n_120), .Y(n_130) );
AO21x2_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_834), .B(n_843), .Y(n_123) );
XOR2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_831), .Y(n_124) );
AOI21x1_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_131), .B(n_520), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g520 ( .A(n_127), .B(n_521), .Y(n_520) );
INVx8_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx12f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g878 ( .A(n_130), .B(n_879), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_132), .A2(n_854), .B1(n_855), .B2(n_861), .Y(n_853) );
INVx2_ASAP7_75t_L g861 ( .A(n_132), .Y(n_861) );
OR2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_452), .Y(n_132) );
NAND4xp25_ASAP7_75t_L g133 ( .A(n_134), .B(n_327), .C(n_367), .D(n_416), .Y(n_133) );
NOR2xp67_ASAP7_75t_L g134 ( .A(n_135), .B(n_276), .Y(n_134) );
OAI22xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_186), .B1(n_248), .B2(n_257), .Y(n_135) );
INVx1_ASAP7_75t_L g448 ( .A(n_136), .Y(n_448) );
INVx1_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_137), .B(n_295), .Y(n_364) );
AND2x2_ASAP7_75t_L g395 ( .A(n_137), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_169), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_138), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g319 ( .A(n_138), .Y(n_319) );
AND2x2_ASAP7_75t_L g494 ( .A(n_138), .B(n_362), .Y(n_494) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx2_ASAP7_75t_L g259 ( .A(n_139), .Y(n_259) );
AND2x2_ASAP7_75t_L g347 ( .A(n_139), .B(n_309), .Y(n_347) );
AND2x2_ASAP7_75t_L g391 ( .A(n_139), .B(n_296), .Y(n_391) );
OR2x2_ASAP7_75t_L g409 ( .A(n_139), .B(n_410), .Y(n_409) );
INVx4_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g313 ( .A(n_140), .B(n_296), .Y(n_313) );
BUFx2_ASAP7_75t_L g370 ( .A(n_140), .Y(n_370) );
OR2x2_ASAP7_75t_L g378 ( .A(n_140), .B(n_336), .Y(n_378) );
INVx1_ASAP7_75t_L g433 ( .A(n_140), .Y(n_433) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_146), .Y(n_140) );
INVx2_ASAP7_75t_L g573 ( .A(n_142), .Y(n_573) );
INVx4_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_SL g165 ( .A(n_143), .B(n_166), .Y(n_165) );
INVx1_ASAP7_75t_SL g172 ( .A(n_143), .Y(n_172) );
INVx2_ASAP7_75t_L g208 ( .A(n_143), .Y(n_208) );
BUFx3_ASAP7_75t_L g529 ( .A(n_143), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_143), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_SL g557 ( .A(n_143), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_143), .B(n_575), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_143), .B(n_596), .Y(n_595) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g185 ( .A(n_144), .Y(n_185) );
OAI21x1_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_156), .B(n_165), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_151), .B(n_153), .Y(n_147) );
OAI22xp33_ASAP7_75t_L g272 ( .A1(n_149), .A2(n_216), .B1(n_273), .B2(n_274), .Y(n_272) );
INVx1_ASAP7_75t_L g547 ( .A(n_149), .Y(n_547) );
INVx4_ASAP7_75t_L g549 ( .A(n_149), .Y(n_549) );
INVx1_ASAP7_75t_L g601 ( .A(n_149), .Y(n_601) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_150), .Y(n_152) );
INVx1_ASAP7_75t_L g162 ( .A(n_150), .Y(n_162) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_150), .Y(n_164) );
INVx1_ASAP7_75t_L g180 ( .A(n_150), .Y(n_180) );
INVx1_ASAP7_75t_L g195 ( .A(n_150), .Y(n_195) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_150), .Y(n_216) );
INVx1_ASAP7_75t_L g225 ( .A(n_150), .Y(n_225) );
INVx1_ASAP7_75t_L g228 ( .A(n_150), .Y(n_228) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_150), .Y(n_241) );
INVx2_ASAP7_75t_L g270 ( .A(n_150), .Y(n_270) );
INVx2_ASAP7_75t_L g201 ( .A(n_152), .Y(n_201) );
INVx1_ASAP7_75t_L g564 ( .A(n_152), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_153), .A2(n_179), .B(n_181), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_153), .A2(n_211), .B(n_212), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_153), .A2(n_300), .B(n_301), .Y(n_299) );
BUFx4f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g160 ( .A(n_155), .Y(n_160) );
INVx1_ASAP7_75t_L g176 ( .A(n_155), .Y(n_176) );
BUFx8_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .B1(n_161), .B2(n_163), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_158), .A2(n_199), .B(n_200), .Y(n_198) );
INVx2_ASAP7_75t_SL g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx3_ASAP7_75t_L g230 ( .A(n_160), .Y(n_230) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OAI21xp5_ASAP7_75t_L g174 ( .A1(n_164), .A2(n_175), .B(n_177), .Y(n_174) );
INVx1_ASAP7_75t_L g245 ( .A(n_164), .Y(n_245) );
INVx3_ASAP7_75t_L g546 ( .A(n_164), .Y(n_546) );
OAI21x1_ASAP7_75t_L g173 ( .A1(n_166), .A2(n_174), .B(n_178), .Y(n_173) );
OAI21x1_ASAP7_75t_L g191 ( .A1(n_166), .A2(n_192), .B(n_198), .Y(n_191) );
OAI21x1_ASAP7_75t_L g209 ( .A1(n_166), .A2(n_210), .B(n_213), .Y(n_209) );
OAI21x1_ASAP7_75t_L g237 ( .A1(n_166), .A2(n_238), .B(n_242), .Y(n_237) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_166), .A2(n_299), .B(n_302), .Y(n_298) );
BUFx10_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx10_ASAP7_75t_L g232 ( .A(n_167), .Y(n_232) );
INVx1_ASAP7_75t_L g536 ( .A(n_167), .Y(n_536) );
AND2x2_ASAP7_75t_L g260 ( .A(n_169), .B(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g372 ( .A(n_169), .B(n_349), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_169), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g410 ( .A(n_170), .Y(n_410) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_170), .Y(n_415) );
AND2x2_ASAP7_75t_L g432 ( .A(n_170), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g322 ( .A(n_171), .B(n_262), .Y(n_322) );
INVx1_ASAP7_75t_L g336 ( .A(n_171), .Y(n_336) );
OAI21x1_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_182), .Y(n_171) );
INVx1_ASAP7_75t_L g246 ( .A(n_176), .Y(n_246) );
INVx1_ASAP7_75t_L g534 ( .A(n_176), .Y(n_534) );
INVx1_ASAP7_75t_SL g550 ( .A(n_176), .Y(n_550) );
INVx1_ASAP7_75t_L g592 ( .A(n_180), .Y(n_592) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g190 ( .A(n_184), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_184), .B(n_604), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_184), .B(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g231 ( .A(n_185), .Y(n_231) );
INVx2_ASAP7_75t_L g235 ( .A(n_185), .Y(n_235) );
NAND2x1_ASAP7_75t_L g186 ( .A(n_187), .B(n_203), .Y(n_186) );
AND2x4_ASAP7_75t_L g497 ( .A(n_187), .B(n_425), .Y(n_497) );
INVxp67_ASAP7_75t_SL g187 ( .A(n_188), .Y(n_187) );
INVxp67_ASAP7_75t_SL g256 ( .A(n_188), .Y(n_256) );
BUFx3_ASAP7_75t_L g291 ( .A(n_188), .Y(n_291) );
INVx1_ASAP7_75t_L g357 ( .A(n_188), .Y(n_357) );
AND2x2_ASAP7_75t_L g360 ( .A(n_188), .B(n_206), .Y(n_360) );
AND2x2_ASAP7_75t_L g385 ( .A(n_188), .B(n_236), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_188), .Y(n_388) );
AND2x2_ASAP7_75t_L g420 ( .A(n_188), .B(n_285), .Y(n_420) );
INVx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
OAI21x1_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_202), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g286 ( .A1(n_190), .A2(n_191), .B(n_202), .Y(n_286) );
OAI21x1_ASAP7_75t_L g297 ( .A1(n_190), .A2(n_298), .B(n_307), .Y(n_297) );
OAI21xp33_ASAP7_75t_SL g325 ( .A1(n_190), .A2(n_298), .B(n_307), .Y(n_325) );
O2A1O1Ixp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_196), .C(n_197), .Y(n_192) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_197), .A2(n_214), .B(n_215), .Y(n_213) );
INVx6_ASAP7_75t_L g226 ( .A(n_197), .Y(n_226) );
O2A1O1Ixp5_ASAP7_75t_L g559 ( .A1(n_197), .A2(n_549), .B(n_560), .C(n_561), .Y(n_559) );
AND2x4_ASAP7_75t_L g203 ( .A(n_204), .B(n_218), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g329 ( .A(n_205), .B(n_315), .Y(n_329) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g355 ( .A(n_207), .B(n_342), .Y(n_355) );
AND2x2_ASAP7_75t_L g384 ( .A(n_207), .B(n_220), .Y(n_384) );
OR2x2_ASAP7_75t_L g480 ( .A(n_207), .B(n_220), .Y(n_480) );
OAI21x1_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_217), .Y(n_207) );
OA21x2_ASAP7_75t_L g236 ( .A1(n_208), .A2(n_237), .B(n_247), .Y(n_236) );
OAI21x1_ASAP7_75t_L g254 ( .A1(n_208), .A2(n_209), .B(n_217), .Y(n_254) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_208), .A2(n_237), .B(n_247), .Y(n_285) );
INVx2_ASAP7_75t_L g223 ( .A(n_216), .Y(n_223) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_216), .A2(n_239), .B(n_240), .Y(n_238) );
AND2x2_ASAP7_75t_L g359 ( .A(n_218), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g508 ( .A(n_218), .Y(n_508) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_219), .Y(n_250) );
OR2x2_ASAP7_75t_L g442 ( .A(n_219), .B(n_252), .Y(n_442) );
INVx1_ASAP7_75t_L g464 ( .A(n_219), .Y(n_464) );
OR2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_236), .Y(n_219) );
AND2x2_ASAP7_75t_L g280 ( .A(n_220), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g315 ( .A(n_220), .B(n_285), .Y(n_315) );
INVx1_ASAP7_75t_L g342 ( .A(n_220), .Y(n_342) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_220), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_220), .B(n_236), .Y(n_429) );
AO31x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_231), .A3(n_232), .B(n_233), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_226), .B1(n_227), .B2(n_229), .Y(n_221) );
INVx1_ASAP7_75t_L g583 ( .A(n_224), .Y(n_583) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_226), .A2(n_531), .B1(n_533), .B2(n_534), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_226), .A2(n_545), .B1(n_548), .B2(n_550), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_226), .A2(n_563), .B(n_565), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_226), .A2(n_229), .B1(n_571), .B2(n_572), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_226), .A2(n_550), .B1(n_582), .B2(n_584), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_226), .A2(n_229), .B1(n_591), .B2(n_593), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_226), .A2(n_229), .B1(n_600), .B2(n_602), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_226), .A2(n_229), .B1(n_616), .B2(n_617), .Y(n_615) );
INVx1_ASAP7_75t_L g594 ( .A(n_228), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_229), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g306 ( .A(n_230), .Y(n_306) );
INVx2_ASAP7_75t_L g264 ( .A(n_231), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_231), .B(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_SL g585 ( .A(n_231), .B(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g265 ( .A(n_232), .Y(n_265) );
AO31x2_ASAP7_75t_L g569 ( .A1(n_232), .A2(n_570), .A3(n_573), .B(n_574), .Y(n_569) );
AO31x2_ASAP7_75t_L g580 ( .A1(n_232), .A2(n_543), .A3(n_581), .B(n_585), .Y(n_580) );
AO31x2_ASAP7_75t_L g589 ( .A1(n_232), .A2(n_529), .A3(n_590), .B(n_595), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
BUFx2_ASAP7_75t_L g543 ( .A(n_235), .Y(n_543) );
AND2x2_ASAP7_75t_L g366 ( .A(n_236), .B(n_286), .Y(n_366) );
INVx2_ASAP7_75t_L g305 ( .A(n_241), .Y(n_305) );
AOI21x1_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_246), .Y(n_242) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NOR3x1_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .C(n_255), .Y(n_249) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_252), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g314 ( .A(n_252), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g365 ( .A(n_252), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g405 ( .A(n_252), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_252), .B(n_428), .Y(n_460) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NOR2xp67_ASAP7_75t_L g401 ( .A(n_253), .B(n_341), .Y(n_401) );
AND2x2_ASAP7_75t_L g425 ( .A(n_253), .B(n_285), .Y(n_425) );
BUFx3_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g281 ( .A(n_254), .Y(n_281) );
BUFx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g436 ( .A(n_256), .B(n_315), .Y(n_436) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_259), .B(n_322), .Y(n_501) );
AND2x4_ASAP7_75t_L g493 ( .A(n_260), .B(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_260), .B(n_313), .Y(n_507) );
INVx2_ASAP7_75t_L g309 ( .A(n_261), .Y(n_309) );
INVx1_ASAP7_75t_L g312 ( .A(n_261), .Y(n_312) );
INVx2_ASAP7_75t_L g397 ( .A(n_261), .Y(n_397) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g381 ( .A(n_262), .Y(n_381) );
AOI21x1_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_266), .B(n_275), .Y(n_262) );
NOR2xp67_ASAP7_75t_SL g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx2_ASAP7_75t_L g598 ( .A(n_264), .Y(n_598) );
INVx1_ASAP7_75t_L g551 ( .A(n_265), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_271), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx2_ASAP7_75t_SL g532 ( .A(n_270), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_316), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_292), .B1(n_310), .B2(n_314), .Y(n_277) );
OAI21xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_282), .B(n_287), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g344 ( .A(n_280), .B(n_291), .Y(n_344) );
AND2x2_ASAP7_75t_L g504 ( .A(n_280), .B(n_385), .Y(n_504) );
BUFx2_ASAP7_75t_L g375 ( .A(n_281), .Y(n_375) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g374 ( .A(n_284), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g289 ( .A(n_285), .Y(n_289) );
INVx1_ASAP7_75t_L g341 ( .A(n_285), .Y(n_341) );
INVx1_ASAP7_75t_L g466 ( .A(n_286), .Y(n_466) );
AOI31xp33_ASAP7_75t_L g484 ( .A1(n_287), .A2(n_485), .A3(n_486), .B(n_487), .Y(n_484) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_288), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_289), .B(n_384), .Y(n_483) );
INVx2_ASAP7_75t_L g511 ( .A(n_289), .Y(n_511) );
INVxp67_ASAP7_75t_SL g326 ( .A(n_290), .Y(n_326) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g339 ( .A(n_291), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_291), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g469 ( .A(n_291), .B(n_429), .Y(n_469) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_308), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g380 ( .A(n_296), .B(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g349 ( .A(n_297), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B(n_306), .Y(n_302) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_312), .Y(n_333) );
INVx1_ASAP7_75t_L g373 ( .A(n_312), .Y(n_373) );
INVx1_ASAP7_75t_L g353 ( .A(n_313), .Y(n_353) );
AND2x2_ASAP7_75t_L g414 ( .A(n_313), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g470 ( .A(n_313), .B(n_397), .Y(n_470) );
OAI21xp5_ASAP7_75t_L g386 ( .A1(n_314), .A2(n_387), .B(n_389), .Y(n_386) );
OR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_326), .Y(n_316) );
NAND3x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .C(n_323), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g488 ( .A(n_319), .B(n_408), .Y(n_488) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NOR2x1_ASAP7_75t_SL g441 ( .A(n_321), .B(n_353), .Y(n_441) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g361 ( .A(n_322), .B(n_362), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_323), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_323), .B(n_432), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_323), .B(n_432), .Y(n_505) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g408 ( .A(n_325), .B(n_381), .Y(n_408) );
AND2x2_ASAP7_75t_L g328 ( .A(n_326), .B(n_329), .Y(n_328) );
AOI221x1_ASAP7_75t_SL g327 ( .A1(n_328), .A2(n_330), .B1(n_337), .B2(n_346), .C(n_350), .Y(n_327) );
AOI32xp33_ASAP7_75t_L g509 ( .A1(n_329), .A2(n_510), .A3(n_515), .B1(n_516), .B2(n_518), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_331), .B(n_334), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_334), .B(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g348 ( .A(n_336), .B(n_349), .Y(n_348) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_336), .Y(n_352) );
OR2x2_ASAP7_75t_L g465 ( .A(n_336), .B(n_466), .Y(n_465) );
NAND3xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_343), .C(n_345), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_L g387 ( .A(n_340), .B(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g404 ( .A(n_340), .B(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_343), .A2(n_440), .B1(n_442), .B2(n_443), .Y(n_439) );
INVx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g517 ( .A(n_347), .Y(n_517) );
INVx2_ASAP7_75t_L g362 ( .A(n_349), .Y(n_362) );
OAI21xp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_354), .B(n_358), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g486 ( .A(n_355), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_356), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_361), .B1(n_363), .B2(n_365), .Y(n_358) );
AND2x4_ASAP7_75t_L g455 ( .A(n_361), .B(n_370), .Y(n_455) );
INVx1_ASAP7_75t_L g514 ( .A(n_362), .Y(n_514) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g393 ( .A(n_366), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_366), .B(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_366), .B(n_394), .Y(n_485) );
AOI211x1_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_374), .B(n_376), .C(n_402), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OR3x2_ASAP7_75t_L g477 ( .A(n_370), .B(n_372), .C(n_373), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_371), .A2(n_393), .B1(n_395), .B2(n_398), .Y(n_392) );
NOR2x1p5_ASAP7_75t_SL g371 ( .A(n_372), .B(n_373), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_372), .A2(n_511), .B1(n_512), .B2(n_513), .Y(n_510) );
INVx2_ASAP7_75t_L g394 ( .A(n_375), .Y(n_394) );
OAI211xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_382), .B(n_386), .C(n_392), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_384), .B(n_388), .Y(n_399) );
INVx1_ASAP7_75t_L g426 ( .A(n_384), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_384), .B(n_491), .Y(n_499) );
OAI32xp33_ASAP7_75t_L g474 ( .A1(n_385), .A2(n_430), .A3(n_475), .B1(n_477), .B2(n_478), .Y(n_474) );
INVx1_ASAP7_75t_L g491 ( .A(n_385), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_385), .B(n_405), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_388), .B(n_422), .Y(n_457) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g435 ( .A(n_394), .B(n_420), .Y(n_435) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g444 ( .A(n_397), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g412 ( .A(n_400), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_406), .B1(n_411), .B2(n_413), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_409), .Y(n_406) );
INVx1_ASAP7_75t_L g450 ( .A(n_407), .Y(n_450) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g431 ( .A(n_408), .B(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_408), .B(n_415), .Y(n_519) );
INVx1_ASAP7_75t_SL g445 ( .A(n_409), .Y(n_445) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NOR3xp33_ASAP7_75t_L g416 ( .A(n_417), .B(n_439), .C(n_446), .Y(n_416) );
OAI21xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_430), .B(n_434), .Y(n_417) );
NOR2xp33_ASAP7_75t_SL g418 ( .A(n_419), .B(n_423), .Y(n_418) );
INVxp67_ASAP7_75t_L g451 ( .A(n_419), .Y(n_451) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g476 ( .A(n_421), .Y(n_476) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NAND3xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_426), .C(n_427), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g438 ( .A(n_432), .Y(n_438) );
OAI21xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_436), .B(n_437), .Y(n_434) );
INVx1_ASAP7_75t_L g447 ( .A(n_435), .Y(n_447) );
OAI221xp5_ASAP7_75t_L g490 ( .A1(n_440), .A2(n_491), .B1(n_492), .B2(n_495), .C(n_496), .Y(n_490) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OAI32xp33_ASAP7_75t_L g446 ( .A1(n_443), .A2(n_447), .A3(n_448), .B1(n_449), .B2(n_451), .Y(n_446) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI221xp5_ASAP7_75t_L g458 ( .A1(n_449), .A2(n_459), .B1(n_460), .B2(n_461), .C(n_467), .Y(n_458) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND3xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_471), .C(n_489), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_456), .B(n_458), .Y(n_453) );
AOI211x1_ASAP7_75t_L g471 ( .A1(n_454), .A2(n_472), .B(n_474), .C(n_481), .Y(n_471) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVxp67_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NOR2x1_ASAP7_75t_SL g462 ( .A(n_463), .B(n_465), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g473 ( .A(n_464), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_470), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AO21x1_ASAP7_75t_L g481 ( .A1(n_470), .A2(n_482), .B(n_484), .Y(n_481) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVxp67_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g515 ( .A(n_486), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_502), .Y(n_489) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OAI21xp33_ASAP7_75t_SL g496 ( .A1(n_497), .A2(n_498), .B(n_500), .Y(n_496) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_509), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_505), .B(n_506), .Y(n_503) );
NOR2xp67_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g512 ( .A(n_511), .Y(n_512) );
INVxp67_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NAND4xp75_ASAP7_75t_L g521 ( .A(n_522), .B(n_671), .C(n_747), .D(n_799), .Y(n_521) );
AND3x1_ASAP7_75t_L g522 ( .A(n_523), .B(n_644), .C(n_657), .Y(n_522) );
AOI221x1_ASAP7_75t_SL g523 ( .A1(n_524), .A2(n_576), .B1(n_605), .B2(n_609), .C(n_621), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g644 ( .A1(n_524), .A2(n_645), .B(n_647), .C(n_648), .Y(n_644) );
AND2x4_ASAP7_75t_L g524 ( .A(n_525), .B(n_539), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g608 ( .A(n_528), .Y(n_608) );
BUFx2_ASAP7_75t_L g626 ( .A(n_528), .Y(n_626) );
OR2x2_ASAP7_75t_L g668 ( .A(n_528), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g675 ( .A(n_528), .B(n_542), .Y(n_675) );
AND2x4_ASAP7_75t_L g710 ( .A(n_528), .B(n_541), .Y(n_710) );
OR2x2_ASAP7_75t_L g753 ( .A(n_528), .B(n_569), .Y(n_753) );
AO31x2_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .A3(n_535), .B(n_537), .Y(n_528) );
AO31x2_ASAP7_75t_L g597 ( .A1(n_535), .A2(n_598), .A3(n_599), .B(n_603), .Y(n_597) );
INVx2_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_SL g566 ( .A(n_536), .Y(n_566) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_554), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_541), .B(n_624), .Y(n_623) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_541), .Y(n_640) );
INVx2_ASAP7_75t_L g667 ( .A(n_541), .Y(n_667) );
INVx3_ASAP7_75t_L g680 ( .A(n_541), .Y(n_680) );
AND2x2_ASAP7_75t_L g798 ( .A(n_541), .B(n_627), .Y(n_798) );
INVx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g607 ( .A(n_542), .B(n_608), .Y(n_607) );
BUFx2_ASAP7_75t_L g663 ( .A(n_542), .Y(n_663) );
AO31x2_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .A3(n_551), .B(n_552), .Y(n_542) );
AO31x2_ASAP7_75t_L g614 ( .A1(n_551), .A2(n_598), .A3(n_615), .B(n_618), .Y(n_614) );
INVxp67_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g683 ( .A(n_555), .Y(n_683) );
INVx1_ASAP7_75t_L g810 ( .A(n_555), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_568), .Y(n_555) );
AND2x2_ASAP7_75t_L g606 ( .A(n_556), .B(n_569), .Y(n_606) );
INVx1_ASAP7_75t_L g669 ( .A(n_556), .Y(n_669) );
OAI21x1_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_558), .B(n_567), .Y(n_556) );
OAI21x1_ASAP7_75t_L g628 ( .A1(n_557), .A2(n_558), .B(n_567), .Y(n_628) );
OAI21x1_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_562), .B(n_566), .Y(n_558) );
INVx2_ASAP7_75t_L g624 ( .A(n_568), .Y(n_624) );
AND2x2_ASAP7_75t_L g676 ( .A(n_568), .B(n_627), .Y(n_676) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g638 ( .A(n_569), .Y(n_638) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_569), .Y(n_698) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_578), .A2(n_670), .B1(n_674), .B2(n_677), .Y(n_673) );
AND2x4_ASAP7_75t_L g578 ( .A(n_579), .B(n_587), .Y(n_578) );
INVx1_ASAP7_75t_L g691 ( .A(n_579), .Y(n_691) );
BUFx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g611 ( .A(n_580), .B(n_589), .Y(n_611) );
AND2x2_ASAP7_75t_L g642 ( .A(n_580), .B(n_597), .Y(n_642) );
INVx4_ASAP7_75t_SL g653 ( .A(n_580), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_580), .B(n_687), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_580), .B(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g724 ( .A(n_588), .B(n_702), .Y(n_724) );
OR2x2_ASAP7_75t_L g757 ( .A(n_588), .B(n_739), .Y(n_757) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_597), .Y(n_588) );
INVx2_ASAP7_75t_L g631 ( .A(n_589), .Y(n_631) );
INVx1_ASAP7_75t_L g636 ( .A(n_589), .Y(n_636) );
AND2x2_ASAP7_75t_L g643 ( .A(n_589), .B(n_613), .Y(n_643) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_589), .Y(n_659) );
INVx1_ASAP7_75t_L g687 ( .A(n_589), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_589), .B(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g620 ( .A(n_597), .Y(n_620) );
AND2x4_ASAP7_75t_L g630 ( .A(n_597), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g656 ( .A(n_597), .Y(n_656) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_597), .Y(n_733) );
INVx1_ASAP7_75t_L g826 ( .A(n_597), .Y(n_826) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_606), .B(n_679), .Y(n_746) );
AND2x2_ASAP7_75t_L g759 ( .A(n_606), .B(n_675), .Y(n_759) );
AND2x2_ASAP7_75t_L g829 ( .A(n_606), .B(n_680), .Y(n_829) );
AND2x4_ASAP7_75t_L g664 ( .A(n_608), .B(n_627), .Y(n_664) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
AND2x2_ASAP7_75t_L g731 ( .A(n_611), .B(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g745 ( .A(n_611), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_611), .B(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g647 ( .A(n_612), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_612), .B(n_685), .Y(n_684) );
AOI211xp5_ASAP7_75t_L g741 ( .A1(n_612), .A2(n_742), .B(n_745), .C(n_746), .Y(n_741) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_620), .Y(n_612) );
AND2x2_ASAP7_75t_L g712 ( .A(n_613), .B(n_653), .Y(n_712) );
INVx3_ASAP7_75t_L g739 ( .A(n_613), .Y(n_739) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g634 ( .A(n_614), .Y(n_634) );
AND2x4_ASAP7_75t_L g660 ( .A(n_614), .B(n_620), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_620), .B(n_653), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_629), .B1(n_637), .B2(n_641), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
INVx1_ASAP7_75t_L g778 ( .A(n_623), .Y(n_778) );
AND2x4_ASAP7_75t_L g689 ( .A(n_624), .B(n_669), .Y(n_689) );
INVx1_ASAP7_75t_L g709 ( .A(n_624), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_626), .A2(n_682), .B1(n_692), .B2(n_694), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_626), .B(n_683), .Y(n_740) );
NAND2x1_ASAP7_75t_L g797 ( .A(n_626), .B(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g812 ( .A(n_626), .Y(n_812) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
BUFx2_ASAP7_75t_L g751 ( .A(n_628), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
AND2x2_ASAP7_75t_L g670 ( .A(n_630), .B(n_652), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_630), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g711 ( .A(n_630), .B(n_712), .Y(n_711) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_630), .Y(n_785) );
NAND2x1p5_ASAP7_75t_L g792 ( .A(n_630), .B(n_693), .Y(n_792) );
AND2x4_ASAP7_75t_L g815 ( .A(n_630), .B(n_743), .Y(n_815) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
INVx3_ASAP7_75t_L g693 ( .A(n_633), .Y(n_693) );
AND2x2_ASAP7_75t_L g705 ( .A(n_633), .B(n_698), .Y(n_705) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g655 ( .A(n_634), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g703 ( .A(n_634), .Y(n_703) );
INVx1_ASAP7_75t_L g646 ( .A(n_635), .Y(n_646) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g803 ( .A(n_636), .B(n_653), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
AND2x2_ASAP7_75t_L g729 ( .A(n_638), .B(n_710), .Y(n_729) );
INVx2_ASAP7_75t_L g770 ( .A(n_638), .Y(n_770) );
AND2x4_ASAP7_75t_L g771 ( .A(n_638), .B(n_664), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_639), .B(n_689), .Y(n_819) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_642), .B(n_702), .Y(n_701) );
AND2x4_ASAP7_75t_L g714 ( .A(n_642), .B(n_659), .Y(n_714) );
INVx1_ASAP7_75t_L g806 ( .A(n_642), .Y(n_806) );
AND2x2_ASAP7_75t_L g805 ( .A(n_643), .B(n_732), .Y(n_805) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OAI22xp33_ASAP7_75t_L g776 ( .A1(n_647), .A2(n_777), .B1(n_779), .B2(n_781), .Y(n_776) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x4_ASAP7_75t_L g650 ( .A(n_651), .B(n_654), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x4_ASAP7_75t_L g685 ( .A(n_653), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g721 ( .A(n_653), .Y(n_721) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_653), .Y(n_727) );
INVx2_ASAP7_75t_L g744 ( .A(n_653), .Y(n_744) );
OR2x2_ASAP7_75t_L g765 ( .A(n_653), .B(n_728), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_653), .B(n_723), .Y(n_775) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OR2x2_ASAP7_75t_L g742 ( .A(n_655), .B(n_743), .Y(n_742) );
HB1xp67_ASAP7_75t_L g796 ( .A(n_655), .Y(n_796) );
INVx1_ASAP7_75t_L g723 ( .A(n_656), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_661), .B(n_665), .Y(n_657) );
AND2x4_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_660), .B(n_691), .Y(n_690) );
INVx3_ASAP7_75t_L g728 ( .A(n_660), .Y(n_728) );
AND2x2_ASAP7_75t_L g802 ( .A(n_660), .B(n_803), .Y(n_802) );
AOI211x1_ASAP7_75t_SL g730 ( .A1(n_661), .A2(n_731), .B(n_734), .C(n_741), .Y(n_730) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x4_ASAP7_75t_L g787 ( .A(n_663), .B(n_664), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_664), .B(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g780 ( .A(n_664), .Y(n_780) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_670), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g695 ( .A(n_667), .Y(n_695) );
NOR2x1p5_ASAP7_75t_L g752 ( .A(n_667), .B(n_753), .Y(n_752) );
NOR2x1_ASAP7_75t_L g696 ( .A(n_668), .B(n_697), .Y(n_696) );
NOR2xp67_ASAP7_75t_SL g769 ( .A(n_668), .B(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g830 ( .A(n_670), .B(n_738), .Y(n_830) );
NOR2x1_ASAP7_75t_L g671 ( .A(n_672), .B(n_715), .Y(n_671) );
NAND3xp33_ASAP7_75t_SL g672 ( .A(n_673), .B(n_681), .C(n_699), .Y(n_672) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_675), .Y(n_706) );
AND2x2_ASAP7_75t_L g713 ( .A(n_675), .B(n_709), .Y(n_713) );
AND2x4_ASAP7_75t_SL g827 ( .A(n_675), .B(n_689), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_676), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_678), .A2(n_720), .B1(n_792), .B2(n_793), .Y(n_791) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AND2x4_ASAP7_75t_L g809 ( .A(n_680), .B(n_810), .Y(n_809) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .B1(n_688), .B2(n_690), .Y(n_682) );
NAND2x1_ASAP7_75t_L g758 ( .A(n_685), .B(n_738), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g768 ( .A(n_685), .B(n_732), .Y(n_768) );
INVx1_ASAP7_75t_L g795 ( .A(n_685), .Y(n_795) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OAI21xp5_ASAP7_75t_L g813 ( .A1(n_688), .A2(n_814), .B(n_817), .Y(n_813) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OAI21xp5_ASAP7_75t_L g700 ( .A1(n_689), .A2(n_701), .B(n_704), .Y(n_700) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g774 ( .A(n_693), .Y(n_774) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVx1_ASAP7_75t_L g718 ( .A(n_696), .Y(n_718) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI222xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_706), .B1(n_707), .B2(n_711), .C1(n_713), .C2(n_714), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g734 ( .A1(n_701), .A2(n_735), .B(n_740), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_702), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g816 ( .A(n_702), .Y(n_816) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
HB1xp67_ASAP7_75t_L g822 ( .A(n_703), .Y(n_822) );
AND2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_710), .Y(n_707) );
AND2x2_ASAP7_75t_L g786 ( .A(n_708), .B(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OR2x2_ASAP7_75t_L g779 ( .A(n_709), .B(n_780), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_730), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_719), .B1(n_725), .B2(n_729), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NAND2xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_724), .Y(n_719) );
OR2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx1_ASAP7_75t_L g736 ( .A(n_722), .Y(n_736) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx4_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OR2x2_ASAP7_75t_L g764 ( .A(n_739), .B(n_756), .Y(n_764) );
OR2x2_ASAP7_75t_L g824 ( .A(n_739), .B(n_825), .Y(n_824) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
NAND5xp2_ASAP7_75t_L g800 ( .A(n_745), .B(n_792), .C(n_801), .D(n_804), .E(n_806), .Y(n_800) );
NOR2x1_ASAP7_75t_L g747 ( .A(n_748), .B(n_783), .Y(n_747) );
NAND2xp67_ASAP7_75t_SL g748 ( .A(n_749), .B(n_766), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_754), .B1(n_759), .B2(n_760), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
NAND3xp33_ASAP7_75t_SL g754 ( .A(n_755), .B(n_757), .C(n_758), .Y(n_754) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g789 ( .A(n_758), .Y(n_789) );
NAND3xp33_ASAP7_75t_SL g760 ( .A(n_761), .B(n_764), .C(n_765), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g782 ( .A(n_763), .Y(n_782) );
O2A1O1Ixp33_ASAP7_75t_SL g794 ( .A1(n_764), .A2(n_795), .B(n_796), .C(n_797), .Y(n_794) );
AOI221xp5_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_769), .B1(n_771), .B2(n_772), .C(n_776), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_773), .B(n_821), .Y(n_820) );
OR2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
INVx1_ASAP7_75t_L g790 ( .A(n_777), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_788), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
INVx1_ASAP7_75t_L g793 ( .A(n_787), .Y(n_793) );
AOI211xp5_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_790), .B(n_791), .C(n_794), .Y(n_788) );
AOI211x1_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_807), .B(n_813), .C(n_828), .Y(n_799) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
NAND2x1p5_ASAP7_75t_L g808 ( .A(n_809), .B(n_811), .Y(n_808) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
NAND2x1_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_820), .B1(n_823), .B2(n_827), .Y(n_817) );
INVxp67_ASAP7_75t_SL g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
AND2x2_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
BUFx12f_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
AND2x6_ASAP7_75t_SL g835 ( .A(n_836), .B(n_838), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx3_ASAP7_75t_L g849 ( .A(n_837), .Y(n_849) );
NOR2xp33_ASAP7_75t_L g876 ( .A(n_837), .B(n_877), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_841), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
NOR2x1_ASAP7_75t_L g879 ( .A(n_840), .B(n_842), .Y(n_879) );
AND2x6_ASAP7_75t_SL g865 ( .A(n_841), .B(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
OAI21xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_850), .B(n_862), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .Y(n_844) );
OAI31xp33_ASAP7_75t_SL g863 ( .A1(n_845), .A2(n_853), .A3(n_864), .B(n_868), .Y(n_863) );
AOI21xp33_ASAP7_75t_SL g862 ( .A1(n_846), .A2(n_863), .B(n_872), .Y(n_862) );
INVx2_ASAP7_75t_SL g846 ( .A(n_847), .Y(n_846) );
BUFx3_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
BUFx8_ASAP7_75t_SL g848 ( .A(n_849), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_851), .B(n_853), .Y(n_850) );
INVx4_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
BUFx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx5_ASAP7_75t_L g871 ( .A(n_865), .Y(n_871) );
OAI21xp5_ASAP7_75t_L g872 ( .A1(n_868), .A2(n_873), .B(n_874), .Y(n_872) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_870), .B(n_871), .Y(n_869) );
INVx5_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
BUFx10_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
NOR2xp33_ASAP7_75t_L g880 ( .A(n_881), .B(n_882), .Y(n_880) );
endmodule