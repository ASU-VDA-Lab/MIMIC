module fake_jpeg_26731_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_4),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_22),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_0),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_26),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_27),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_25),
.A2(n_17),
.B1(n_15),
.B2(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_31),
.B(n_32),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_2),
.B(n_13),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_39),
.B(n_3),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_26),
.B(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_34),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_49),
.Y(n_53)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_43),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_22),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_21),
.B1(n_17),
.B2(n_12),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_21),
.B1(n_12),
.B2(n_19),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_27),
.C(n_28),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_29),
.C(n_35),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_32),
.B(n_31),
.C(n_35),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_56),
.B1(n_44),
.B2(n_43),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_46),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_52),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_55),
.C(n_48),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_29),
.C(n_10),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_49),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_60),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_61),
.Y(n_65)
);

FAx1_ASAP7_75t_SL g60 ( 
.A(n_55),
.B(n_41),
.CI(n_42),
.CON(n_60),
.SN(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_19),
.B1(n_14),
.B2(n_30),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_30),
.C(n_10),
.Y(n_62)
);

A2O1A1O1Ixp25_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_53),
.B(n_11),
.C(n_50),
.D(n_10),
.Y(n_63)
);

AOI322xp5_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_57),
.A3(n_62),
.B1(n_58),
.B2(n_13),
.C1(n_14),
.C2(n_8),
.Y(n_67)
);

FAx1_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_53),
.CI(n_11),
.CON(n_66),
.SN(n_66)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_66),
.B(n_5),
.Y(n_68)
);

AOI31xp67_ASAP7_75t_SL g69 ( 
.A1(n_67),
.A2(n_66),
.A3(n_64),
.B(n_8),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_7),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_70),
.C(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_65),
.Y(n_72)
);


endmodule