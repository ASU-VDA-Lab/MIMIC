module real_jpeg_8020_n_21 (n_17, n_8, n_0, n_82, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_81, n_1, n_20, n_19, n_16, n_15, n_13, n_21);

input n_17;
input n_8;
input n_0;
input n_82;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_81;
input n_1;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_21;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_49;
wire n_68;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_26;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_61;
wire n_70;
wire n_41;
wire n_74;
wire n_32;
wire n_30;
wire n_57;
wire n_43;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_0),
.A2(n_11),
.B(n_28),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_0),
.B(n_30),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_1),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_3),
.A2(n_14),
.B(n_32),
.Y(n_51)
);

NAND3xp33_ASAP7_75t_SL g52 ( 
.A(n_3),
.B(n_14),
.C(n_32),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_4),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_6),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_8),
.A2(n_18),
.B(n_32),
.Y(n_63)
);

NAND3xp33_ASAP7_75t_L g64 ( 
.A(n_8),
.B(n_18),
.C(n_32),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_9),
.A2(n_20),
.B(n_32),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_SL g58 ( 
.A(n_9),
.B(n_20),
.C(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_25),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_10),
.A2(n_45),
.B(n_46),
.Y(n_44)
);

NOR3xp33_ASAP7_75t_L g50 ( 
.A(n_10),
.B(n_45),
.C(n_46),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_10),
.A2(n_54),
.B(n_55),
.Y(n_53)
);

NOR3xp33_ASAP7_75t_L g56 ( 
.A(n_10),
.B(n_54),
.C(n_55),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_10),
.A2(n_60),
.B(n_61),
.Y(n_59)
);

NOR3xp33_ASAP7_75t_L g62 ( 
.A(n_10),
.B(n_60),
.C(n_61),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_10),
.A2(n_66),
.B(n_67),
.Y(n_65)
);

NOR3xp33_ASAP7_75t_L g68 ( 
.A(n_10),
.B(n_66),
.C(n_67),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_11),
.B(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_11),
.A2(n_12),
.B(n_28),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_11),
.B(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_11),
.B(n_17),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_12),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_13),
.B(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_16),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_17),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_19),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_33),
.B2(n_34),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_31),
.B(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_31),
.A2(n_78),
.B(n_79),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_82),
.Y(n_49)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI311xp33_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_71),
.A3(n_72),
.B1(n_73),
.C1(n_74),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NOR3xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_69),
.C(n_70),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_65),
.B(n_68),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_63),
.B(n_64),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_59),
.B(n_62),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_57),
.B(n_58),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_53),
.B(n_56),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_51),
.B(n_52),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B(n_50),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_81),
.Y(n_45)
);


endmodule