module fake_jpeg_28309_n_297 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_297);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_0),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_6),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_14),
.B1(n_17),
.B2(n_16),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_47),
.B1(n_14),
.B2(n_29),
.Y(n_57)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_42),
.Y(n_54)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_14),
.B1(n_17),
.B2(n_20),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_24),
.C(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_35),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_13),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_29),
.B1(n_28),
.B2(n_14),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_50),
.B1(n_45),
.B2(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_53),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_64),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_68),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_58),
.B1(n_71),
.B2(n_26),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_26),
.B1(n_16),
.B2(n_13),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVxp67_ASAP7_75t_SL g91 ( 
.A(n_59),
.Y(n_91)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_60),
.Y(n_77)
);

AO22x1_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_30),
.B1(n_35),
.B2(n_32),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_90)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_22),
.B(n_24),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_SL g87 ( 
.A(n_63),
.B(n_24),
.C(n_23),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_49),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_67),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_69),
.B(n_18),
.Y(n_80)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_66),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_26),
.B1(n_13),
.B2(n_18),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_50),
.B1(n_45),
.B2(n_42),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_74),
.A2(n_78),
.B1(n_87),
.B2(n_88),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_76),
.A2(n_86),
.B1(n_82),
.B2(n_85),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_50),
.B1(n_45),
.B2(n_39),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_39),
.B1(n_43),
.B2(n_41),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_57),
.B1(n_58),
.B2(n_68),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_92),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_94),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_64),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_67),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_111),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_92),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_100),
.B(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_104),
.Y(n_128)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_56),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_31),
.C(n_80),
.Y(n_129)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_107),
.B(n_108),
.Y(n_139)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_53),
.Y(n_109)
);

BUFx24_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_76),
.B1(n_61),
.B2(n_62),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_117),
.B1(n_84),
.B2(n_81),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_115),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_88),
.A2(n_61),
.B1(n_71),
.B2(n_59),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_116),
.A2(n_73),
.B1(n_65),
.B2(n_60),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_83),
.A2(n_61),
.B1(n_59),
.B2(n_62),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_134),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_83),
.B(n_87),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_130),
.B(n_132),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_133),
.B1(n_95),
.B2(n_116),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_125),
.A2(n_136),
.B1(n_144),
.B2(n_23),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_61),
.B1(n_73),
.B2(n_70),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_126),
.A2(n_44),
.B1(n_23),
.B2(n_24),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_106),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_100),
.B(n_98),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_77),
.B(n_75),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_131),
.A2(n_138),
.B(n_141),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_31),
.B(n_75),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_60),
.B1(n_65),
.B2(n_77),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_115),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_143),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_105),
.A2(n_25),
.B(n_24),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_108),
.A2(n_72),
.B1(n_66),
.B2(n_25),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_104),
.A2(n_72),
.B1(n_43),
.B2(n_41),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_148),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_173),
.B1(n_174),
.B2(n_168),
.Y(n_186)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_149),
.B(n_19),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_96),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_151),
.B(n_154),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_110),
.B(n_25),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_118),
.B(n_115),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_152),
.Y(n_178)
);

INVxp33_ASAP7_75t_SL g153 ( 
.A(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_110),
.B(n_25),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_124),
.C(n_134),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_164),
.C(n_167),
.Y(n_179)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_160),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_141),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_139),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_168),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_43),
.Y(n_163)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_32),
.C(n_43),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_129),
.B(n_132),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_15),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_126),
.B(n_36),
.C(n_110),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_122),
.B(n_131),
.C(n_125),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_136),
.C(n_137),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_120),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_170),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_140),
.B(n_119),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_171),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_120),
.Y(n_172)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

AO21x2_ASAP7_75t_SL g173 ( 
.A1(n_138),
.A2(n_44),
.B(n_24),
.Y(n_173)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_189),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_143),
.C(n_135),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_158),
.C(n_159),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_186),
.A2(n_190),
.B1(n_200),
.B2(n_173),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_188),
.B(n_196),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_145),
.B(n_15),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_146),
.A2(n_23),
.B1(n_19),
.B2(n_22),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_145),
.B(n_15),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_199),
.Y(n_214)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_155),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_8),
.C(n_1),
.Y(n_195)
);

NOR3xp33_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_165),
.C(n_172),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_149),
.B(n_15),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_198),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_148),
.A2(n_23),
.B1(n_19),
.B2(n_22),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_169),
.B1(n_173),
.B2(n_174),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_204),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_183),
.B(n_150),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_208),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_211),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_192),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_210),
.Y(n_238)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_197),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_198),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_216),
.Y(n_235)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_196),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_173),
.B1(n_160),
.B2(n_156),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_217),
.A2(n_218),
.B(n_220),
.Y(n_233)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_186),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_150),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

BUFx12_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_154),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_179),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_226),
.C(n_231),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_179),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_220),
.A2(n_156),
.B(n_157),
.C(n_176),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_157),
.B(n_219),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_228),
.B(n_230),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_180),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_188),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_205),
.C(n_214),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_239),
.C(n_151),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_199),
.C(n_187),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_202),
.B1(n_219),
.B2(n_216),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_240),
.A2(n_231),
.B1(n_224),
.B2(n_228),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_238),
.B(n_163),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_245),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_223),
.B1(n_233),
.B2(n_235),
.Y(n_243)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_243),
.Y(n_259)
);

OAI321xp33_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_230),
.A3(n_237),
.B1(n_226),
.B2(n_175),
.C(n_4),
.Y(n_256)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_229),
.Y(n_245)
);

NAND4xp25_ASAP7_75t_SL g246 ( 
.A(n_236),
.B(n_221),
.C(n_200),
.D(n_190),
.Y(n_246)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_225),
.B(n_164),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_247),
.B(n_248),
.Y(n_254)
);

OAI21xp33_ASAP7_75t_L g248 ( 
.A1(n_227),
.A2(n_176),
.B(n_189),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_251),
.Y(n_260)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_239),
.A2(n_214),
.B1(n_167),
.B2(n_191),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_252),
.B(n_253),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_253),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_256),
.A2(n_264),
.B(n_7),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_23),
.C(n_19),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_265),
.C(n_22),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_240),
.B(n_22),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_246),
.Y(n_266)
);

OAI321xp33_ASAP7_75t_L g264 ( 
.A1(n_248),
.A2(n_23),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_22),
.C(n_0),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_269),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_267),
.B(n_270),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_252),
.B(n_250),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_268),
.A2(n_272),
.B(n_273),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_0),
.C(n_2),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_271),
.B(n_5),
.Y(n_283)
);

AOI21xp33_ASAP7_75t_L g272 ( 
.A1(n_258),
.A2(n_2),
.B(n_3),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_3),
.B(n_4),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_3),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_275),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_4),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_5),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_5),
.Y(n_284)
);

NAND4xp25_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_265),
.C(n_261),
.D(n_7),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_9),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_270),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_283),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_284),
.A2(n_9),
.B(n_10),
.Y(n_289)
);

AOI21x1_ASAP7_75t_L g285 ( 
.A1(n_281),
.A2(n_6),
.B(n_7),
.Y(n_285)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_285),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_279),
.A2(n_8),
.B(n_9),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_288),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_282),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_SL g294 ( 
.A1(n_290),
.A2(n_11),
.B(n_12),
.C(n_292),
.Y(n_294)
);

NOR4xp25_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_278),
.C(n_287),
.D(n_280),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_293),
.A2(n_294),
.B(n_11),
.Y(n_295)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_11),
.C(n_12),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_12),
.Y(n_297)
);


endmodule