module real_jpeg_18529_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_546;
wire n_285;
wire n_172;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B(n_545),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_0),
.B(n_546),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_1),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_1),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_1),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_1),
.B(n_29),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_1),
.B(n_169),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_1),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_1),
.B(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_1),
.A2(n_3),
.B1(n_288),
.B2(n_290),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_1),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_2),
.Y(n_105)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_2),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_3),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_3),
.B(n_241),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_3),
.B(n_356),
.Y(n_355)
);

AOI31xp33_ASAP7_75t_SL g388 ( 
.A1(n_3),
.A2(n_287),
.A3(n_389),
.B(n_391),
.Y(n_388)
);

NAND2x1_ASAP7_75t_SL g430 ( 
.A(n_3),
.B(n_431),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_3),
.B(n_73),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_3),
.B(n_455),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_3),
.B(n_503),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_4),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_4),
.Y(n_212)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_4),
.Y(n_244)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_4),
.Y(n_409)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_5),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_5),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_5),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_6),
.Y(n_107)
);

NAND2x1_ASAP7_75t_SL g109 ( 
.A(n_6),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_6),
.B(n_250),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g268 ( 
.A(n_6),
.B(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_SL g306 ( 
.A(n_6),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_6),
.B(n_73),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_6),
.B(n_396),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_6),
.B(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_7),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_7),
.B(n_62),
.Y(n_61)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_7),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_7),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_7),
.B(n_214),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_7),
.B(n_300),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_7),
.B(n_316),
.Y(n_315)
);

AND2x2_ASAP7_75t_SL g353 ( 
.A(n_7),
.B(n_258),
.Y(n_353)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_8),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_8),
.Y(n_201)
);

BUFx4f_ASAP7_75t_L g398 ( 
.A(n_8),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_8),
.Y(n_457)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_9),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_10),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_10),
.B(n_406),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_10),
.B(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_10),
.B(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_10),
.B(n_494),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_10),
.B(n_508),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_10),
.B(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_11),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_11),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_11),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g136 ( 
.A(n_11),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_11),
.B(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_12),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_12),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_13),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_13),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_13),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_13),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_13),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_13),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_13),
.B(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_14),
.Y(n_118)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_14),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_14),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_15),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_15),
.B(n_133),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_15),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_15),
.B(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_15),
.B(n_361),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_15),
.B(n_459),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_15),
.B(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_15),
.B(n_311),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_16),
.B(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_16),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_16),
.B(n_90),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_16),
.B(n_246),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_16),
.B(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_16),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_16),
.B(n_400),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_17),
.Y(n_98)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

BUFx8_ASAP7_75t_L g110 ( 
.A(n_18),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_18),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_177),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_175),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_149),
.Y(n_22)
);

NOR2xp67_ASAP7_75t_SL g176 ( 
.A(n_23),
.B(n_149),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_114),
.C(n_125),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_24),
.B(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_80),
.C(n_100),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_26),
.B(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_43),
.C(n_60),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_27),
.B(n_43),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_28),
.B(n_33),
.C(n_38),
.Y(n_124)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_31),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_38),
.Y(n_32)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_42),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_50),
.C(n_55),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_44),
.B(n_55),
.Y(n_193)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_48),
.Y(n_432)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

XNOR2x1_ASAP7_75t_L g192 ( 
.A(n_50),
.B(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_54),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_59),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_60),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_68),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_61),
.B(n_70),
.C(n_74),
.Y(n_123)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_65),
.Y(n_269)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_67),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_74),
.B2(n_75),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_69),
.A2(n_70),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_SL g128 ( 
.A(n_70),
.B(n_117),
.C(n_120),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_74),
.A2(n_75),
.B1(n_103),
.B2(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

MAJx2_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_103),
.C(n_106),
.Y(n_102)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_78),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_80),
.B(n_100),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_81),
.B(n_88),
.C(n_99),
.Y(n_140)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_86),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_94),
.B2(n_99),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_93),
.Y(n_252)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_96),
.Y(n_322)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_97),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_98),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_109),
.C(n_111),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_101),
.A2(n_102),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_103),
.B(n_195),
.C(n_198),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_103),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_103),
.A2(n_198),
.B1(n_206),
.B2(n_238),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_105),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_106),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_106),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_106),
.A2(n_203),
.B1(n_299),
.B2(n_348),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_109),
.B(n_111),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_109),
.B(n_257),
.C(n_261),
.Y(n_256)
);

XNOR2x2_ASAP7_75t_SL g284 ( 
.A(n_109),
.B(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_111),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_111),
.A2(n_219),
.B1(n_220),
.B2(n_273),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_114),
.A2(n_125),
.B1(n_126),
.B2(n_182),
.Y(n_181)
);

INVxp33_ASAP7_75t_SL g182 ( 
.A(n_114),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_123),
.C(n_124),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_115),
.B(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_117),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_119),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_119),
.B(n_130),
.C(n_136),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_123),
.B(n_124),
.Y(n_188)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_139),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_129),
.C(n_139),
.Y(n_174)
);

XOR2x1_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_135),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_136),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_138),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_142),
.C(n_143),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_174),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_166),
.B2(n_167),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_161),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx2_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_168),
.Y(n_172)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_170),
.Y(n_309)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_225),
.B(n_541),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_179),
.A2(n_543),
.B(n_544),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_180),
.B(n_183),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_189),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_184),
.A2(n_185),
.B1(n_187),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_187),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_189),
.B(n_275),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_207),
.C(n_221),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_230),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.C(n_202),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_192),
.B(n_194),
.Y(n_331)
);

XNOR2x1_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_198),
.Y(n_238)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_201),
.Y(n_263)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_201),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_202),
.Y(n_330)
);

MAJx2_ASAP7_75t_L g293 ( 
.A(n_203),
.B(n_294),
.C(n_299),
.Y(n_293)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_222),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_219),
.C(n_220),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_208),
.B(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_213),
.C(n_218),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_209),
.B(n_218),
.Y(n_254)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_219),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_223),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_277),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_274),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_228),
.B(n_274),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.C(n_234),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_229),
.B(n_231),
.Y(n_371)
);

XNOR2x1_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_234),
.B(n_371),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_255),
.C(n_270),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_235),
.B(n_328),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.C(n_253),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_236),
.B(n_239),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_245),
.C(n_248),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_240),
.A2(n_248),
.B1(n_249),
.B2(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_240),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_245),
.B(n_367),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_247),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_248),
.B(n_426),
.C(n_430),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_248),
.A2(n_249),
.B1(n_426),
.B2(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2x1_ASAP7_75t_L g340 ( 
.A(n_253),
.B(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_255),
.B(n_271),
.Y(n_328)
);

MAJx2_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_264),
.C(n_267),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g324 ( 
.A(n_256),
.B(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_261),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_260),
.Y(n_402)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_264),
.B(n_268),
.Y(n_325)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_265),
.Y(n_509)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_267),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_267),
.A2(n_268),
.B1(n_404),
.B2(n_405),
.Y(n_525)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

AO21x2_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_375),
.B(n_538),
.Y(n_277)
);

NOR2xp67_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_369),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_334),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_280),
.B(n_334),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_326),
.Y(n_280)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_281),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_303),
.C(n_323),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_283),
.B(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.C(n_293),
.Y(n_283)
);

XNOR2x1_ASAP7_75t_L g410 ( 
.A(n_284),
.B(n_411),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_286),
.A2(n_287),
.B1(n_293),
.B2(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_289),
.B(n_392),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_293),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_294),
.B(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_298),
.Y(n_450)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_299),
.Y(n_348)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_304),
.A2(n_323),
.B1(n_324),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_304),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_314),
.C(n_321),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_305),
.B(n_364),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.C(n_310),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_306),
.B(n_310),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_306),
.B(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_306),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_308),
.B(n_387),
.Y(n_386)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_314),
.A2(n_315),
.B1(n_321),
.B2(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx6_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_321),
.Y(n_365)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_329),
.B1(n_332),
.B2(n_333),
.Y(n_326)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_327),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_329),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_329),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_332),
.B(n_373),
.C(n_374),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_340),
.C(n_342),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_336),
.A2(n_337),
.B1(n_340),
.B2(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_340),
.Y(n_380)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_343),
.B(n_379),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_363),
.C(n_366),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_344),
.B(n_384),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_349),
.C(n_354),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

XNOR2x1_ASAP7_75t_SL g435 ( 
.A(n_346),
.B(n_436),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_349),
.B(n_354),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_353),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_350),
.B(n_353),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_352),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_359),
.C(n_360),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_355),
.A2(n_359),
.B1(n_422),
.B2(n_423),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_355),
.Y(n_422)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_359),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_359),
.B(n_490),
.C(n_492),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_359),
.A2(n_423),
.B1(n_492),
.B2(n_493),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_360),
.B(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_362),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_363),
.B(n_366),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_369),
.A2(n_539),
.B(n_540),
.Y(n_538)
);

AND2x2_ASAP7_75t_SL g369 ( 
.A(n_370),
.B(n_372),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g540 ( 
.A(n_370),
.B(n_372),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_437),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_381),
.C(n_413),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_378),
.B(n_382),
.Y(n_439)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_385),
.C(n_410),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_383),
.B(n_415),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_385),
.B(n_410),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_388),
.C(n_393),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_386),
.B(n_388),
.Y(n_418)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_393),
.B(n_418),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_403),
.C(n_404),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g524 ( 
.A(n_394),
.B(n_525),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_399),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_395),
.B(n_399),
.Y(n_476)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_395),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_395),
.A2(n_501),
.B1(n_502),
.B2(n_511),
.Y(n_510)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_402),
.Y(n_460)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

NOR2x1_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_416),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_414),
.B(n_416),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_419),
.C(n_435),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_417),
.B(n_536),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_419),
.B(n_435),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_424),
.C(n_433),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_420),
.B(n_530),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_425),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_425),
.B(n_434),
.Y(n_530)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_426),
.Y(n_483)
);

INVx8_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

XOR2x2_ASAP7_75t_L g481 ( 
.A(n_430),
.B(n_482),
.Y(n_481)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

NAND3xp33_ASAP7_75t_SL g437 ( 
.A(n_438),
.B(n_439),
.C(n_440),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_441),
.A2(n_533),
.B(n_537),
.Y(n_440)
);

AOI21x1_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_519),
.B(n_532),
.Y(n_441)
);

OAI21x1_ASAP7_75t_SL g442 ( 
.A1(n_443),
.A2(n_484),
.B(n_518),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_472),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_444),
.B(n_472),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_452),
.C(n_461),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_445),
.B(n_487),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_451),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_447),
.B(n_451),
.C(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_452),
.A2(n_453),
.B1(n_461),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_458),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g491 ( 
.A(n_454),
.B(n_458),
.Y(n_491)
);

INVx5_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_457),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_461),
.Y(n_488)
);

AO22x1_ASAP7_75t_SL g461 ( 
.A1(n_462),
.A2(n_467),
.B1(n_470),
.B2(n_471),
.Y(n_461)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_462),
.Y(n_470)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_467),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_467),
.B(n_470),
.Y(n_474)
);

INVx6_ASAP7_75t_L g504 ( 
.A(n_468),
.Y(n_504)
);

INVx5_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_471),
.B(n_513),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_478),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_473),
.B(n_479),
.C(n_481),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_475),
.Y(n_473)
);

MAJx2_ASAP7_75t_L g527 ( 
.A(n_474),
.B(n_476),
.C(n_477),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_481),
.Y(n_478)
);

AOI21x1_ASAP7_75t_L g484 ( 
.A1(n_485),
.A2(n_495),
.B(n_517),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_486),
.B(n_489),
.Y(n_485)
);

NOR2x1_ASAP7_75t_L g517 ( 
.A(n_486),
.B(n_489),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_490),
.A2(n_491),
.B1(n_498),
.B2(n_499),
.Y(n_497)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_496),
.A2(n_505),
.B(n_516),
.Y(n_495)
);

NOR2xp67_ASAP7_75t_SL g496 ( 
.A(n_497),
.B(n_500),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_497),
.B(n_500),
.Y(n_516)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_501),
.B(n_502),
.Y(n_500)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_502),
.Y(n_511)
);

INVx5_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_506),
.A2(n_512),
.B(n_515),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_510),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_507),
.B(n_510),
.Y(n_515)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_520),
.B(n_531),
.Y(n_519)
);

NOR2x1p5_ASAP7_75t_L g532 ( 
.A(n_520),
.B(n_531),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_521),
.A2(n_522),
.B1(n_528),
.B2(n_529),
.Y(n_520)
);

INVxp67_ASAP7_75t_SL g521 ( 
.A(n_522),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_523),
.A2(n_524),
.B1(n_526),
.B2(n_527),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_523),
.B(n_527),
.C(n_528),
.Y(n_534)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

NOR2xp67_ASAP7_75t_SL g533 ( 
.A(n_534),
.B(n_535),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_534),
.B(n_535),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);


endmodule