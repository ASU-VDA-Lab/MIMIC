module fake_jpeg_18195_n_284 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_284);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_SL g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

NAND2xp33_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_43),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_22),
.B(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_37),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_30),
.B1(n_19),
.B2(n_24),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_33),
.B1(n_34),
.B2(n_30),
.Y(n_67)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_37),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_59),
.B(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_61),
.Y(n_108)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_63),
.B(n_65),
.Y(n_116)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_67),
.A2(n_68),
.B1(n_75),
.B2(n_84),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_33),
.B1(n_40),
.B2(n_42),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_19),
.B1(n_30),
.B2(n_13),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_69),
.A2(n_91),
.B1(n_92),
.B2(n_27),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_42),
.B1(n_24),
.B2(n_19),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_71),
.A2(n_94),
.B1(n_75),
.B2(n_26),
.Y(n_128)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx8_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_13),
.B(n_37),
.C(n_17),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_80),
.Y(n_127)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_82),
.Y(n_102)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_54),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_87),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_13),
.B1(n_31),
.B2(n_22),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_51),
.B(n_31),
.Y(n_85)
);

BUFx24_ASAP7_75t_SL g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_86),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_20),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_52),
.B(n_18),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_89),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_53),
.B(n_18),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_28),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_96),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_45),
.A2(n_17),
.B1(n_14),
.B2(n_26),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_50),
.A2(n_44),
.B1(n_41),
.B2(n_15),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_100),
.B1(n_15),
.B2(n_41),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_20),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_36),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_23),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_23),
.Y(n_130)
);

INVxp33_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_76),
.B1(n_77),
.B2(n_64),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_68),
.A2(n_59),
.B(n_99),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_120),
.A2(n_23),
.B(n_25),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_66),
.Y(n_147)
);

AOI22x1_ASAP7_75t_L g123 ( 
.A1(n_59),
.A2(n_44),
.B1(n_36),
.B2(n_35),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_128),
.B1(n_131),
.B2(n_90),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_71),
.A2(n_15),
.B1(n_27),
.B2(n_32),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_97),
.B1(n_72),
.B2(n_21),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_130),
.B(n_23),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_60),
.A2(n_62),
.B1(n_98),
.B2(n_93),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_100),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_137),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_99),
.C(n_90),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_155),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_138),
.A2(n_140),
.B1(n_126),
.B2(n_123),
.Y(n_177)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_128),
.A2(n_71),
.B1(n_70),
.B2(n_74),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_106),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_144),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_71),
.B(n_86),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_143),
.A2(n_151),
.B(n_154),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_106),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_104),
.A2(n_70),
.B(n_23),
.C(n_82),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_35),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_149),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_32),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_79),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_152),
.Y(n_171)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_105),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_112),
.A2(n_25),
.B(n_23),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_109),
.B1(n_127),
.B2(n_108),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_157),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_131),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_148),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_139),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_161),
.B(n_168),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_115),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_167),
.B(n_185),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_141),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_172),
.A2(n_158),
.B1(n_134),
.B2(n_154),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_126),
.B1(n_123),
.B2(n_104),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_173),
.A2(n_177),
.B1(n_184),
.B2(n_144),
.Y(n_192)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_142),
.Y(n_200)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g178 ( 
.A1(n_143),
.A2(n_132),
.B1(n_107),
.B2(n_125),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_178),
.A2(n_179),
.B(n_16),
.Y(n_205)
);

AND2x6_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_113),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_116),
.Y(n_181)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_140),
.A2(n_102),
.B1(n_121),
.B2(n_124),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_72),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_187),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_201),
.B1(n_173),
.B2(n_169),
.Y(n_212)
);

INVxp33_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_191),
.Y(n_211)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_192),
.A2(n_204),
.B1(n_172),
.B2(n_180),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_170),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_197),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_200),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_170),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_146),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_198),
.B(n_118),
.Y(n_227)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_199),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_159),
.A2(n_153),
.B1(n_152),
.B2(n_117),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_182),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_202),
.B(n_206),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_159),
.A2(n_105),
.B(n_6),
.C(n_11),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_205),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_177),
.A2(n_145),
.B1(n_118),
.B2(n_9),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_169),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_166),
.C(n_185),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_213),
.C(n_198),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_212),
.A2(n_218),
.B1(n_220),
.B2(n_192),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_166),
.C(n_180),
.Y(n_213)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_226),
.Y(n_236)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_217),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_175),
.B1(n_178),
.B2(n_161),
.Y(n_218)
);

AND2x6_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_179),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_219),
.A2(n_224),
.B(n_221),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_201),
.A2(n_178),
.B1(n_168),
.B2(n_164),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_178),
.B1(n_164),
.B2(n_183),
.Y(n_222)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_160),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_213),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_231),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_233),
.Y(n_254)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_189),
.B1(n_191),
.B2(n_160),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_234),
.B(n_237),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_208),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_240),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_225),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_207),
.C(n_193),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_242),
.C(n_244),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_226),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_239),
.B(n_243),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_203),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_186),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_187),
.B(n_207),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_194),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_241),
.A2(n_221),
.B1(n_216),
.B2(n_215),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_249),
.B1(n_256),
.B2(n_8),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_229),
.A2(n_220),
.B1(n_215),
.B2(n_217),
.Y(n_249)
);

XNOR2x1_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_223),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_251),
.A2(n_252),
.B1(n_8),
.B2(n_12),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_145),
.C(n_176),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_230),
.C(n_235),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_240),
.B1(n_242),
.B2(n_244),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_259),
.C(n_265),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_253),
.A2(n_231),
.B(n_163),
.Y(n_258)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_254),
.C(n_1),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_21),
.C(n_16),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_260),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_262),
.Y(n_269)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_263),
.A2(n_252),
.B1(n_251),
.B2(n_245),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_8),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_245),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_21),
.C(n_25),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_268),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_254),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_21),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_265),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_257),
.C(n_258),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_274),
.A2(n_275),
.B(n_276),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_266),
.C(n_271),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_278),
.B(n_279),
.Y(n_280)
);

O2A1O1Ixp33_ASAP7_75t_SL g279 ( 
.A1(n_274),
.A2(n_272),
.B(n_266),
.C(n_9),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_281),
.A2(n_277),
.B1(n_6),
.B2(n_5),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_282),
.A2(n_5),
.B(n_6),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_11),
.Y(n_284)
);


endmodule