module real_aes_16750_n_267 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_1490, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_267);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_1490;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_267;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1172;
wire n_459;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_1185;
wire n_661;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1170;
wire n_1175;
wire n_778;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_273;
wire n_1038;
wire n_1085;
wire n_276;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp5_ASAP7_75t_L g1236 ( .A1(n_0), .A2(n_204), .B1(n_1209), .B2(n_1224), .Y(n_1236) );
CKINVDCx5p33_ASAP7_75t_R g840 ( .A(n_1), .Y(n_840) );
OAI22xp33_ASAP7_75t_L g1440 ( .A1(n_2), .A2(n_92), .B1(n_675), .B2(n_678), .Y(n_1440) );
INVxp67_ASAP7_75t_SL g1453 ( .A(n_2), .Y(n_1453) );
CKINVDCx5p33_ASAP7_75t_R g800 ( .A(n_3), .Y(n_800) );
INVx1_ASAP7_75t_L g1118 ( .A(n_4), .Y(n_1118) );
AOI221xp5_ASAP7_75t_L g1164 ( .A1(n_5), .A2(n_209), .B1(n_463), .B2(n_863), .C(n_1165), .Y(n_1164) );
INVx1_ASAP7_75t_L g1190 ( .A(n_5), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g1232 ( .A1(n_6), .A2(n_59), .B1(n_1209), .B2(n_1224), .Y(n_1232) );
INVx1_ASAP7_75t_L g1425 ( .A(n_7), .Y(n_1425) );
INVx1_ASAP7_75t_L g321 ( .A(n_8), .Y(n_321) );
OAI221xp5_ASAP7_75t_SL g412 ( .A1(n_8), .A2(n_93), .B1(n_413), .B2(n_414), .C(n_418), .Y(n_412) );
INVx1_ASAP7_75t_L g1166 ( .A(n_9), .Y(n_1166) );
AOI221xp5_ASAP7_75t_L g1192 ( .A1(n_9), .A2(n_161), .B1(n_588), .B2(n_716), .C(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g487 ( .A(n_10), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_10), .A2(n_116), .B1(n_319), .B2(n_537), .Y(n_536) );
AOI21xp33_ASAP7_75t_L g1131 ( .A1(n_11), .A2(n_627), .B(n_633), .Y(n_1131) );
INVx1_ASAP7_75t_L g1153 ( .A(n_11), .Y(n_1153) );
OAI221xp5_ASAP7_75t_L g476 ( .A1(n_12), .A2(n_220), .B1(n_413), .B2(n_414), .C(n_435), .Y(n_476) );
OA222x2_ASAP7_75t_L g552 ( .A1(n_12), .A2(n_50), .B1(n_226), .B2(n_553), .C1(n_557), .C2(n_561), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_13), .A2(n_73), .B1(n_547), .B2(n_596), .Y(n_909) );
OAI22xp33_ASAP7_75t_L g952 ( .A1(n_13), .A2(n_37), .B1(n_675), .B2(n_678), .Y(n_952) );
AOI221xp5_ASAP7_75t_L g980 ( .A1(n_14), .A2(n_241), .B1(n_348), .B2(n_981), .C(n_983), .Y(n_980) );
INVx1_ASAP7_75t_L g1001 ( .A(n_14), .Y(n_1001) );
INVx1_ASAP7_75t_L g282 ( .A(n_15), .Y(n_282) );
AND2x2_ASAP7_75t_L g323 ( .A(n_15), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g335 ( .A(n_15), .B(n_231), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_15), .B(n_292), .Y(n_515) );
AOI221xp5_ASAP7_75t_L g1027 ( .A1(n_16), .A2(n_199), .B1(n_463), .B2(n_1028), .C(n_1030), .Y(n_1027) );
INVx1_ASAP7_75t_L g1053 ( .A(n_16), .Y(n_1053) );
INVx1_ASAP7_75t_L g1065 ( .A(n_17), .Y(n_1065) );
OAI221xp5_ASAP7_75t_SL g1095 ( .A1(n_17), .A2(n_259), .B1(n_1096), .B2(n_1099), .C(n_1102), .Y(n_1095) );
INVx1_ASAP7_75t_L g594 ( .A(n_18), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_18), .A2(n_253), .B1(n_612), .B2(n_615), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_19), .A2(n_123), .B1(n_658), .B2(n_660), .Y(n_657) );
INVxp67_ASAP7_75t_SL g708 ( .A(n_19), .Y(n_708) );
INVx2_ASAP7_75t_L g1212 ( .A(n_20), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_20), .B(n_111), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_20), .B(n_1218), .Y(n_1220) );
AOI21xp5_ASAP7_75t_L g1437 ( .A1(n_21), .A2(n_411), .B(n_1438), .Y(n_1437) );
INVx1_ASAP7_75t_L g1464 ( .A(n_21), .Y(n_1464) );
INVx1_ASAP7_75t_L g837 ( .A(n_22), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g1249 ( .A1(n_23), .A2(n_34), .B1(n_1216), .B2(n_1219), .Y(n_1249) );
AOI22xp33_ASAP7_75t_L g1446 ( .A1(n_24), .A2(n_162), .B1(n_506), .B2(n_623), .Y(n_1446) );
AOI32xp33_ASAP7_75t_L g1455 ( .A1(n_24), .A2(n_318), .A3(n_1456), .B1(n_1458), .B2(n_1490), .Y(n_1455) );
XNOR2x2_ASAP7_75t_L g1159 ( .A(n_25), .B(n_1160), .Y(n_1159) );
INVx1_ASAP7_75t_L g673 ( .A(n_26), .Y(n_673) );
INVx1_ASAP7_75t_L g1126 ( .A(n_27), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1148 ( .A1(n_27), .A2(n_153), .B1(n_327), .B2(n_590), .Y(n_1148) );
AOI22xp5_ASAP7_75t_L g1235 ( .A1(n_28), .A2(n_127), .B1(n_1216), .B2(n_1219), .Y(n_1235) );
AOI22xp5_ASAP7_75t_L g1258 ( .A1(n_29), .A2(n_137), .B1(n_1209), .B2(n_1245), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_30), .B(n_861), .Y(n_1439) );
AOI221xp5_ASAP7_75t_L g1467 ( .A1(n_30), .A2(n_162), .B1(n_314), .B2(n_824), .C(n_1089), .Y(n_1467) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_31), .A2(n_183), .B1(n_672), .B2(n_861), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_31), .A2(n_147), .B1(n_884), .B2(n_890), .Y(n_889) );
AOI222xp33_ASAP7_75t_L g685 ( .A1(n_32), .A2(n_189), .B1(n_219), .B2(n_464), .C1(n_497), .C2(n_633), .Y(n_685) );
INVx1_ASAP7_75t_L g719 ( .A(n_32), .Y(n_719) );
CKINVDCx5p33_ASAP7_75t_R g747 ( .A(n_33), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_35), .B(n_1435), .Y(n_1434) );
AOI22xp33_ASAP7_75t_L g1466 ( .A1(n_35), .A2(n_264), .B1(n_588), .B2(n_715), .Y(n_1466) );
INVx1_ASAP7_75t_L g577 ( .A(n_36), .Y(n_577) );
OAI211xp5_ASAP7_75t_L g906 ( .A1(n_37), .A2(n_907), .B(n_908), .C(n_930), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_38), .A2(n_106), .B1(n_1209), .B2(n_1213), .Y(n_1208) );
INVx1_ASAP7_75t_L g1167 ( .A(n_39), .Y(n_1167) );
AOI221xp5_ASAP7_75t_L g1185 ( .A1(n_39), .A2(n_74), .B1(n_1186), .B2(n_1187), .C(n_1189), .Y(n_1185) );
AOI22xp5_ASAP7_75t_L g1244 ( .A1(n_40), .A2(n_98), .B1(n_1209), .B2(n_1245), .Y(n_1244) );
INVx1_ASAP7_75t_L g845 ( .A(n_41), .Y(n_845) );
AOI211xp5_ASAP7_75t_L g1019 ( .A1(n_42), .A2(n_625), .B(n_1020), .C(n_1022), .Y(n_1019) );
INVx1_ASAP7_75t_L g1050 ( .A(n_42), .Y(n_1050) );
OAI221xp5_ASAP7_75t_L g1176 ( .A1(n_43), .A2(n_67), .B1(n_615), .B2(n_619), .C(n_656), .Y(n_1176) );
INVxp67_ASAP7_75t_SL g1181 ( .A(n_43), .Y(n_1181) );
INVx1_ASAP7_75t_L g987 ( .A(n_44), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_45), .A2(n_78), .B1(n_863), .B2(n_999), .Y(n_1070) );
INVxp67_ASAP7_75t_SL g1104 ( .A(n_45), .Y(n_1104) );
OAI21xp33_ASAP7_75t_L g579 ( .A1(n_46), .A2(n_553), .B(n_580), .Y(n_579) );
OAI221xp5_ASAP7_75t_L g635 ( .A1(n_46), .A2(n_54), .B1(n_636), .B2(n_637), .C(n_639), .Y(n_635) );
OAI22xp33_ASAP7_75t_L g810 ( .A1(n_47), .A2(n_180), .B1(n_615), .B2(n_656), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_47), .A2(n_83), .B1(n_545), .B2(n_550), .Y(n_829) );
OAI211xp5_ASAP7_75t_SL g1114 ( .A1(n_48), .A2(n_642), .B(n_1115), .C(n_1119), .Y(n_1114) );
INVx1_ASAP7_75t_L g1138 ( .A(n_48), .Y(n_1138) );
INVx1_ASAP7_75t_L g381 ( .A(n_49), .Y(n_381) );
INVx1_ASAP7_75t_L g402 ( .A(n_49), .Y(n_402) );
INVx1_ASAP7_75t_L g474 ( .A(n_50), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_51), .A2(n_164), .B1(n_329), .B2(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g433 ( .A(n_51), .Y(n_433) );
OAI221xp5_ASAP7_75t_L g1016 ( .A1(n_52), .A2(n_247), .B1(n_615), .B2(n_619), .C(n_656), .Y(n_1016) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_52), .A2(n_132), .B1(n_547), .B2(n_596), .Y(n_1041) );
INVx1_ASAP7_75t_L g597 ( .A(n_53), .Y(n_597) );
INVxp67_ASAP7_75t_SL g647 ( .A(n_54), .Y(n_647) );
CKINVDCx5p33_ASAP7_75t_R g737 ( .A(n_55), .Y(n_737) );
CKINVDCx5p33_ASAP7_75t_R g752 ( .A(n_56), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g1215 ( .A1(n_57), .A2(n_230), .B1(n_1216), .B2(n_1219), .Y(n_1215) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_58), .A2(n_170), .B1(n_664), .B2(n_666), .C(n_668), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_58), .A2(n_225), .B1(n_713), .B2(n_715), .C(n_717), .Y(n_712) );
OAI221xp5_ASAP7_75t_L g655 ( .A1(n_60), .A2(n_246), .B1(n_615), .B2(n_619), .C(n_656), .Y(n_655) );
OAI21xp33_ASAP7_75t_SL g696 ( .A1(n_60), .A2(n_539), .B(n_561), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_61), .A2(n_240), .B1(n_658), .B2(n_660), .Y(n_937) );
INVxp67_ASAP7_75t_SL g957 ( .A(n_61), .Y(n_957) );
INVx1_ASAP7_75t_L g275 ( .A(n_62), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g1175 ( .A1(n_63), .A2(n_215), .B1(n_658), .B2(n_660), .Y(n_1175) );
INVx1_ASAP7_75t_L g1184 ( .A(n_63), .Y(n_1184) );
INVx2_ASAP7_75t_L g388 ( .A(n_64), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g1163 ( .A1(n_65), .A2(n_194), .B1(n_675), .B2(n_678), .Y(n_1163) );
INVx1_ASAP7_75t_L g1182 ( .A(n_65), .Y(n_1182) );
INVx1_ASAP7_75t_L g797 ( .A(n_66), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_66), .A2(n_228), .B1(n_329), .B2(n_358), .Y(n_823) );
INVx1_ASAP7_75t_L g1200 ( .A(n_67), .Y(n_1200) );
INVxp67_ASAP7_75t_SL g971 ( .A(n_68), .Y(n_971) );
OAI211xp5_ASAP7_75t_L g1008 ( .A1(n_68), .A2(n_619), .B(n_642), .C(n_1009), .Y(n_1008) );
CKINVDCx5p33_ASAP7_75t_R g809 ( .A(n_69), .Y(n_809) );
OAI22xp33_ASAP7_75t_L g674 ( .A1(n_70), .A2(n_72), .B1(n_675), .B2(n_678), .Y(n_674) );
INVxp67_ASAP7_75t_SL g691 ( .A(n_70), .Y(n_691) );
INVx1_ASAP7_75t_L g758 ( .A(n_71), .Y(n_758) );
INVx1_ASAP7_75t_L g695 ( .A(n_72), .Y(n_695) );
OAI221xp5_ASAP7_75t_L g936 ( .A1(n_73), .A2(n_125), .B1(n_615), .B2(n_619), .C(n_656), .Y(n_936) );
AOI221xp5_ASAP7_75t_L g1168 ( .A1(n_74), .A2(n_211), .B1(n_463), .B2(n_1169), .C(n_1170), .Y(n_1168) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_75), .A2(n_190), .B1(n_348), .B2(n_354), .C(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g434 ( .A(n_75), .Y(n_434) );
INVx1_ASAP7_75t_L g654 ( .A(n_76), .Y(n_654) );
OAI21xp33_ASAP7_75t_L g692 ( .A1(n_76), .A2(n_557), .B(n_693), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_77), .A2(n_244), .B1(n_633), .B2(n_1072), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_77), .A2(n_217), .B1(n_314), .B2(n_1089), .Y(n_1088) );
AOI221xp5_ASAP7_75t_L g1084 ( .A1(n_78), .A2(n_104), .B1(n_881), .B2(n_893), .C(n_1085), .Y(n_1084) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_79), .Y(n_481) );
INVx1_ASAP7_75t_L g973 ( .A(n_80), .Y(n_973) );
INVx1_ASAP7_75t_L g491 ( .A(n_81), .Y(n_491) );
AOI221x1_ASAP7_75t_SL g516 ( .A1(n_81), .A2(n_101), .B1(n_348), .B2(n_358), .C(n_517), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g1479 ( .A1(n_82), .A2(n_1480), .B1(n_1481), .B2(n_1482), .Y(n_1479) );
CKINVDCx20_ASAP7_75t_R g1482 ( .A(n_82), .Y(n_1482) );
OAI221xp5_ASAP7_75t_L g805 ( .A1(n_83), .A2(n_179), .B1(n_806), .B2(n_807), .C(n_808), .Y(n_805) );
OAI222xp33_ASAP7_75t_L g764 ( .A1(n_84), .A2(n_131), .B1(n_237), .B2(n_393), .C1(n_490), .C2(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g782 ( .A(n_84), .Y(n_782) );
XOR2x2_ASAP7_75t_L g1011 ( .A(n_85), .B(n_1012), .Y(n_1011) );
AOI22xp33_ASAP7_75t_SL g851 ( .A1(n_86), .A2(n_97), .B1(n_852), .B2(n_854), .Y(n_851) );
AOI221xp5_ASAP7_75t_L g880 ( .A1(n_86), .A2(n_130), .B1(n_318), .B2(n_715), .C(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g1135 ( .A(n_87), .Y(n_1135) );
AOI22xp5_ASAP7_75t_L g1225 ( .A1(n_88), .A2(n_129), .B1(n_1216), .B2(n_1219), .Y(n_1225) );
XOR2x1_ASAP7_75t_L g1420 ( .A(n_88), .B(n_1421), .Y(n_1420) );
AOI22xp33_ASAP7_75t_L g1474 ( .A1(n_88), .A2(n_1475), .B1(n_1478), .B2(n_1483), .Y(n_1474) );
AOI22xp33_ASAP7_75t_L g1241 ( .A1(n_89), .A2(n_114), .B1(n_1209), .B2(n_1224), .Y(n_1241) );
INVx1_ASAP7_75t_L g925 ( .A(n_90), .Y(n_925) );
AOI221xp5_ASAP7_75t_L g1127 ( .A1(n_91), .A2(n_145), .B1(n_629), .B2(n_770), .C(n_1128), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g1154 ( .A1(n_91), .A2(n_198), .B1(n_327), .B2(n_366), .Y(n_1154) );
INVx1_ASAP7_75t_L g1422 ( .A(n_92), .Y(n_1422) );
INVx1_ASAP7_75t_L g340 ( .A(n_93), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_94), .A2(n_234), .B1(n_603), .B2(n_604), .Y(n_975) );
AOI21xp33_ASAP7_75t_L g1004 ( .A1(n_94), .A2(n_505), .B(n_627), .Y(n_1004) );
INVx1_ASAP7_75t_L g469 ( .A(n_95), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_95), .A2(n_220), .B1(n_545), .B2(n_550), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_96), .A2(n_132), .B1(n_675), .B2(n_678), .Y(n_1026) );
OAI211xp5_ASAP7_75t_L g1034 ( .A1(n_96), .A2(n_907), .B(n_1035), .C(n_1038), .Y(n_1034) );
AOI221xp5_ASAP7_75t_L g891 ( .A1(n_97), .A2(n_210), .B1(n_892), .B2(n_893), .C(n_897), .Y(n_891) );
INVx1_ASAP7_75t_L g751 ( .A(n_99), .Y(n_751) );
AOI221xp5_ASAP7_75t_L g769 ( .A1(n_99), .A2(n_159), .B1(n_463), .B2(n_770), .C(n_773), .Y(n_769) );
OAI221xp5_ASAP7_75t_L g305 ( .A1(n_100), .A2(n_265), .B1(n_306), .B2(n_308), .C(n_313), .Y(n_305) );
INVx1_ASAP7_75t_L g372 ( .A(n_100), .Y(n_372) );
INVx1_ASAP7_75t_L g507 ( .A(n_101), .Y(n_507) );
INVx1_ASAP7_75t_L g1025 ( .A(n_102), .Y(n_1025) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_103), .Y(n_277) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_103), .B(n_275), .Y(n_1210) );
AOI22xp33_ASAP7_75t_SL g1077 ( .A1(n_104), .A2(n_175), .B1(n_374), .B2(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g1032 ( .A(n_105), .Y(n_1032) );
OAI21xp5_ASAP7_75t_SL g900 ( .A1(n_107), .A2(n_901), .B(n_902), .Y(n_900) );
INVx1_ASAP7_75t_L g959 ( .A(n_108), .Y(n_959) );
AOI22xp33_ASAP7_75t_SL g587 ( .A1(n_109), .A2(n_193), .B1(n_350), .B2(n_588), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_109), .A2(n_184), .B1(n_625), .B2(n_626), .C(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g1068 ( .A(n_110), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_111), .B(n_1212), .Y(n_1211) );
INVx1_ASAP7_75t_L g1218 ( .A(n_111), .Y(n_1218) );
AOI221xp5_ASAP7_75t_L g1441 ( .A1(n_112), .A2(n_264), .B1(n_1003), .B2(n_1442), .C(n_1445), .Y(n_1441) );
INVx1_ASAP7_75t_L g1465 ( .A(n_112), .Y(n_1465) );
AOI22xp5_ASAP7_75t_L g1257 ( .A1(n_113), .A2(n_181), .B1(n_1216), .B2(n_1219), .Y(n_1257) );
INVx1_ASAP7_75t_L g1031 ( .A(n_115), .Y(n_1031) );
INVx1_ASAP7_75t_L g498 ( .A(n_116), .Y(n_498) );
XNOR2xp5_ASAP7_75t_L g831 ( .A(n_117), .B(n_832), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g1427 ( .A1(n_118), .A2(n_257), .B1(n_658), .B2(n_660), .Y(n_1427) );
INVxp33_ASAP7_75t_L g1469 ( .A(n_118), .Y(n_1469) );
INVx1_ASAP7_75t_L g332 ( .A(n_119), .Y(n_332) );
OAI21xp33_ASAP7_75t_L g405 ( .A1(n_119), .A2(n_406), .B(n_410), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_120), .B(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g425 ( .A(n_120), .Y(n_425) );
INVx1_ASAP7_75t_L g453 ( .A(n_120), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g792 ( .A(n_121), .Y(n_792) );
INVx1_ASAP7_75t_L g759 ( .A(n_122), .Y(n_759) );
OAI22xp33_ASAP7_75t_L g767 ( .A1(n_122), .A2(n_168), .B1(n_615), .B2(n_656), .Y(n_767) );
INVxp67_ASAP7_75t_SL g688 ( .A(n_123), .Y(n_688) );
INVxp67_ASAP7_75t_SL g1130 ( .A(n_124), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_124), .A2(n_145), .B1(n_1144), .B2(n_1146), .Y(n_1143) );
INVxp67_ASAP7_75t_SL g932 ( .A(n_125), .Y(n_932) );
OAI221xp5_ASAP7_75t_L g1426 ( .A1(n_126), .A2(n_166), .B1(n_615), .B2(n_619), .C(n_656), .Y(n_1426) );
NOR2xp33_ASAP7_75t_L g1457 ( .A(n_126), .B(n_584), .Y(n_1457) );
XOR2xp5_ASAP7_75t_L g454 ( .A(n_127), .B(n_455), .Y(n_454) );
AOI221xp5_ASAP7_75t_L g926 ( .A1(n_128), .A2(n_154), .B1(n_920), .B2(n_927), .C(n_929), .Y(n_926) );
AOI221xp5_ASAP7_75t_L g948 ( .A1(n_128), .A2(n_167), .B1(n_411), .B2(n_941), .C(n_949), .Y(n_948) );
AOI221xp5_ASAP7_75t_L g862 ( .A1(n_130), .A2(n_147), .B1(n_854), .B2(n_863), .C(n_864), .Y(n_862) );
OAI221xp5_ASAP7_75t_L g755 ( .A1(n_131), .A2(n_168), .B1(n_539), .B2(n_545), .C(n_550), .Y(n_755) );
INVx1_ASAP7_75t_L g726 ( .A(n_133), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_134), .A2(n_300), .B1(n_301), .B2(n_302), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_134), .Y(n_300) );
AOI22xp33_ASAP7_75t_SL g589 ( .A1(n_135), .A2(n_254), .B1(n_364), .B2(n_590), .Y(n_589) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_135), .A2(n_214), .B1(n_411), .B2(n_625), .C(n_629), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g1242 ( .A1(n_136), .A2(n_238), .B1(n_1216), .B2(n_1219), .Y(n_1242) );
AOI22xp5_ASAP7_75t_L g1223 ( .A1(n_138), .A2(n_141), .B1(n_1209), .B2(n_1224), .Y(n_1223) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_139), .Y(n_494) );
INVx1_ASAP7_75t_L g923 ( .A(n_140), .Y(n_923) );
AOI221xp5_ASAP7_75t_L g939 ( .A1(n_140), .A2(n_266), .B1(n_940), .B2(n_941), .C(n_942), .Y(n_939) );
OAI22xp33_ASAP7_75t_L g470 ( .A1(n_142), .A2(n_151), .B1(n_471), .B2(n_472), .Y(n_470) );
INVx1_ASAP7_75t_L g570 ( .A(n_142), .Y(n_570) );
INVx1_ASAP7_75t_L g1174 ( .A(n_143), .Y(n_1174) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_144), .A2(n_195), .B1(n_364), .B2(n_365), .Y(n_363) );
INVx1_ASAP7_75t_L g447 ( .A(n_144), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g1111 ( .A1(n_146), .A2(n_1112), .B1(n_1157), .B2(n_1158), .Y(n_1111) );
INVx1_ASAP7_75t_L g1158 ( .A(n_146), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g1231 ( .A1(n_148), .A2(n_149), .B1(n_1216), .B2(n_1219), .Y(n_1231) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_150), .A2(n_660), .B1(n_795), .B2(n_798), .Y(n_794) );
INVx1_ASAP7_75t_L g816 ( .A(n_150), .Y(n_816) );
INVx1_ASAP7_75t_L g566 ( .A(n_151), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_152), .A2(n_160), .B1(n_658), .B2(n_660), .Y(n_1017) );
INVxp67_ASAP7_75t_SL g1039 ( .A(n_152), .Y(n_1039) );
AOI22xp33_ASAP7_75t_SL g1132 ( .A1(n_153), .A2(n_198), .B1(n_623), .B2(n_1133), .Y(n_1132) );
INVx1_ASAP7_75t_L g945 ( .A(n_154), .Y(n_945) );
INVx1_ASAP7_75t_L g984 ( .A(n_155), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_155), .A2(n_222), .B1(n_623), .B2(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g1120 ( .A(n_156), .Y(n_1120) );
OAI221xp5_ASAP7_75t_L g1140 ( .A1(n_156), .A2(n_197), .B1(n_550), .B2(n_1141), .C(n_1142), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_157), .A2(n_213), .B1(n_364), .B2(n_600), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_157), .A2(n_254), .B1(n_411), .B2(n_623), .Y(n_622) );
AOI221xp5_ASAP7_75t_SL g347 ( .A1(n_158), .A2(n_185), .B1(n_348), .B2(n_354), .C(n_355), .Y(n_347) );
INVx1_ASAP7_75t_L g437 ( .A(n_158), .Y(n_437) );
INVx1_ASAP7_75t_L g733 ( .A(n_159), .Y(n_733) );
INVxp67_ASAP7_75t_SL g1036 ( .A(n_160), .Y(n_1036) );
INVx1_ASAP7_75t_L g1171 ( .A(n_161), .Y(n_1171) );
BUFx3_ASAP7_75t_L g378 ( .A(n_163), .Y(n_378) );
INVx1_ASAP7_75t_L g449 ( .A(n_164), .Y(n_449) );
INVx1_ASAP7_75t_L g1121 ( .A(n_165), .Y(n_1121) );
INVxp67_ASAP7_75t_SL g1452 ( .A(n_166), .Y(n_1452) );
AOI221xp5_ASAP7_75t_L g917 ( .A1(n_167), .A2(n_207), .B1(n_824), .B2(n_918), .C(n_920), .Y(n_917) );
AOI22xp5_ASAP7_75t_L g1246 ( .A1(n_169), .A2(n_171), .B1(n_1216), .B2(n_1219), .Y(n_1246) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_170), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g1021 ( .A(n_172), .Y(n_1021) );
INVx1_ASAP7_75t_L g670 ( .A(n_173), .Y(n_670) );
INVx1_ASAP7_75t_L g988 ( .A(n_174), .Y(n_988) );
INVxp67_ASAP7_75t_SL g1105 ( .A(n_175), .Y(n_1105) );
AOI22xp5_ASAP7_75t_L g1250 ( .A1(n_176), .A2(n_232), .B1(n_1209), .B2(n_1224), .Y(n_1250) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_177), .Y(n_289) );
INVx1_ASAP7_75t_L g581 ( .A(n_178), .Y(n_581) );
OAI211xp5_ASAP7_75t_L g814 ( .A1(n_179), .A2(n_646), .B(n_815), .C(n_818), .Y(n_814) );
INVx1_ASAP7_75t_L g817 ( .A(n_180), .Y(n_817) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_182), .Y(n_791) );
AOI22xp33_ASAP7_75t_SL g882 ( .A1(n_183), .A2(n_258), .B1(n_883), .B2(n_884), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_184), .A2(n_214), .B1(n_603), .B2(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g446 ( .A(n_185), .Y(n_446) );
OAI222xp33_ASAP7_75t_L g1079 ( .A1(n_186), .A2(n_216), .B1(n_236), .B2(n_835), .C1(n_839), .C2(n_901), .Y(n_1079) );
OAI211xp5_ASAP7_75t_L g1081 ( .A1(n_186), .A2(n_1082), .B(n_1083), .C(n_1090), .Y(n_1081) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_187), .Y(n_345) );
INVx1_ASAP7_75t_L g972 ( .A(n_188), .Y(n_972) );
INVx1_ASAP7_75t_L g704 ( .A(n_189), .Y(n_704) );
INVx1_ASAP7_75t_L g450 ( .A(n_190), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g746 ( .A(n_191), .Y(n_746) );
INVx1_ASAP7_75t_L g802 ( .A(n_192), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_192), .A2(n_196), .B1(n_329), .B2(n_366), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_193), .A2(n_213), .B1(n_623), .B2(n_631), .Y(n_630) );
INVxp67_ASAP7_75t_SL g1198 ( .A(n_194), .Y(n_1198) );
INVx1_ASAP7_75t_L g443 ( .A(n_195), .Y(n_443) );
AOI221xp5_ASAP7_75t_L g789 ( .A1(n_196), .A2(n_228), .B1(n_623), .B2(n_772), .C(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g1136 ( .A(n_197), .Y(n_1136) );
INVx1_ASAP7_75t_L g1045 ( .A(n_199), .Y(n_1045) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_200), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_201), .Y(n_484) );
INVx1_ASAP7_75t_L g1023 ( .A(n_202), .Y(n_1023) );
CKINVDCx5p33_ASAP7_75t_R g796 ( .A(n_203), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g741 ( .A(n_205), .Y(n_741) );
INVxp67_ASAP7_75t_SL g757 ( .A(n_206), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_206), .A2(n_660), .B1(n_775), .B2(n_776), .Y(n_774) );
INVx1_ASAP7_75t_L g943 ( .A(n_207), .Y(n_943) );
INVx1_ASAP7_75t_L g931 ( .A(n_208), .Y(n_931) );
INVx1_ASAP7_75t_L g1194 ( .A(n_209), .Y(n_1194) );
AOI22xp33_ASAP7_75t_SL g867 ( .A1(n_210), .A2(n_258), .B1(n_852), .B2(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g1196 ( .A(n_211), .Y(n_1196) );
INVx1_ASAP7_75t_L g1431 ( .A(n_212), .Y(n_1431) );
INVxp67_ASAP7_75t_SL g1178 ( .A(n_215), .Y(n_1178) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_217), .A2(n_242), .B1(n_1074), .B2(n_1075), .Y(n_1073) );
OAI21xp5_ASAP7_75t_L g991 ( .A1(n_218), .A2(n_992), .B(n_993), .Y(n_991) );
OAI22xp5_ASAP7_75t_L g994 ( .A1(n_218), .A2(n_233), .B1(n_658), .B2(n_660), .Y(n_994) );
AOI21xp33_ASAP7_75t_L g706 ( .A1(n_219), .A2(n_318), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g968 ( .A(n_221), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_222), .A2(n_252), .B1(n_358), .B2(n_537), .Y(n_976) );
INVx1_ASAP7_75t_L g1015 ( .A(n_223), .Y(n_1015) );
INVx1_ASAP7_75t_L g872 ( .A(n_224), .Y(n_872) );
AOI21xp33_ASAP7_75t_L g680 ( .A1(n_225), .A2(n_681), .B(n_684), .Y(n_680) );
INVx1_ASAP7_75t_L g465 ( .A(n_226), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g734 ( .A(n_227), .Y(n_734) );
INVx1_ASAP7_75t_L g843 ( .A(n_229), .Y(n_843) );
INVx1_ASAP7_75t_L g1010 ( .A(n_230), .Y(n_1010) );
BUFx3_ASAP7_75t_L g292 ( .A(n_231), .Y(n_292) );
INVx1_ASAP7_75t_L g324 ( .A(n_231), .Y(n_324) );
INVxp33_ASAP7_75t_L g990 ( .A(n_233), .Y(n_990) );
INVx1_ASAP7_75t_L g997 ( .A(n_234), .Y(n_997) );
INVx1_ASAP7_75t_L g1116 ( .A(n_235), .Y(n_1116) );
INVx1_ASAP7_75t_L g761 ( .A(n_237), .Y(n_761) );
INVx2_ASAP7_75t_L g369 ( .A(n_239), .Y(n_369) );
INVx1_ASAP7_75t_L g386 ( .A(n_239), .Y(n_386) );
INVx1_ASAP7_75t_L g421 ( .A(n_239), .Y(n_421) );
INVxp67_ASAP7_75t_SL g933 ( .A(n_240), .Y(n_933) );
AOI221xp5_ASAP7_75t_L g998 ( .A1(n_241), .A2(n_252), .B1(n_374), .B2(n_629), .C(n_999), .Y(n_998) );
AOI221xp5_ASAP7_75t_L g1106 ( .A1(n_242), .A2(n_244), .B1(n_318), .B2(n_699), .C(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g1172 ( .A(n_243), .Y(n_1172) );
INVx1_ASAP7_75t_L g875 ( .A(n_245), .Y(n_875) );
INVx1_ASAP7_75t_L g694 ( .A(n_246), .Y(n_694) );
INVxp67_ASAP7_75t_SL g1037 ( .A(n_247), .Y(n_1037) );
INVx1_ASAP7_75t_L g785 ( .A(n_248), .Y(n_785) );
INVx1_ASAP7_75t_L g1067 ( .A(n_249), .Y(n_1067) );
XOR2x2_ASAP7_75t_L g650 ( .A(n_250), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g804 ( .A(n_251), .Y(n_804) );
INVx1_ASAP7_75t_L g582 ( .A(n_253), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_255), .Y(n_502) );
INVx1_ASAP7_75t_L g1124 ( .A(n_256), .Y(n_1124) );
INVxp67_ASAP7_75t_SL g1448 ( .A(n_257), .Y(n_1448) );
INVx1_ASAP7_75t_L g1064 ( .A(n_259), .Y(n_1064) );
XNOR2xp5_ASAP7_75t_L g1059 ( .A(n_260), .B(n_1060), .Y(n_1059) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_261), .Y(n_573) );
NAND2xp33_ASAP7_75t_SL g915 ( .A(n_262), .B(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g950 ( .A(n_262), .Y(n_950) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_263), .Y(n_317) );
INVx1_ASAP7_75t_L g390 ( .A(n_265), .Y(n_390) );
INVx1_ASAP7_75t_L g912 ( .A(n_266), .Y(n_912) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_293), .B(n_1202), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx3_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_278), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g1473 ( .A(n_272), .B(n_281), .Y(n_1473) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g1477 ( .A(n_274), .B(n_277), .Y(n_1477) );
INVx1_ASAP7_75t_L g1486 ( .A(n_274), .Y(n_1486) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g1488 ( .A(n_277), .B(n_1486), .Y(n_1488) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g356 ( .A(n_282), .B(n_291), .Y(n_356) );
AND2x4_ASAP7_75t_L g362 ( .A(n_282), .B(n_292), .Y(n_362) );
AND2x4_ASAP7_75t_SL g1472 ( .A(n_283), .B(n_1473), .Y(n_1472) );
INVx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x6_ASAP7_75t_L g284 ( .A(n_285), .B(n_290), .Y(n_284) );
BUFx4f_ASAP7_75t_L g703 ( .A(n_285), .Y(n_703) );
INVxp67_ASAP7_75t_L g750 ( .A(n_285), .Y(n_750) );
INVx1_ASAP7_75t_L g986 ( .A(n_285), .Y(n_986) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx4f_ASAP7_75t_L g307 ( .A(n_286), .Y(n_307) );
INVx3_ASAP7_75t_L g519 ( .A(n_286), .Y(n_519) );
INVx3_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx2_ASAP7_75t_L g312 ( .A(n_288), .Y(n_312) );
INVx2_ASAP7_75t_L g316 ( .A(n_288), .Y(n_316) );
AND2x2_ASAP7_75t_L g320 ( .A(n_288), .B(n_289), .Y(n_320) );
INVx1_ASAP7_75t_L g344 ( .A(n_288), .Y(n_344) );
AND2x2_ASAP7_75t_L g352 ( .A(n_288), .B(n_353), .Y(n_352) );
NAND2x1_ASAP7_75t_L g522 ( .A(n_288), .B(n_289), .Y(n_522) );
OR2x2_ASAP7_75t_L g311 ( .A(n_289), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g315 ( .A(n_289), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g331 ( .A(n_289), .Y(n_331) );
BUFx2_ASAP7_75t_L g339 ( .A(n_289), .Y(n_339) );
INVx2_ASAP7_75t_L g353 ( .A(n_289), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_289), .B(n_316), .Y(n_535) );
INVxp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OAI22xp33_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_962), .B1(n_963), .B2(n_1201), .Y(n_293) );
INVx1_ASAP7_75t_L g1201 ( .A(n_294), .Y(n_1201) );
BUFx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
XOR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_722), .Y(n_295) );
XNOR2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_571), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
XNOR2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_454), .Y(n_298) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_370), .Y(n_302) );
AOI21xp5_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_346), .B(n_367), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_322), .B(n_325), .Y(n_304) );
INVx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx6f_ASAP7_75t_L g1048 ( .A(n_307), .Y(n_1048) );
INVx4_ASAP7_75t_L g1191 ( .A(n_307), .Y(n_1191) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_308), .A2(n_1021), .B1(n_1044), .B2(n_1045), .Y(n_1043) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx4_ASAP7_75t_L g740 ( .A(n_309), .Y(n_740) );
INVx2_ASAP7_75t_L g1152 ( .A(n_309), .Y(n_1152) );
INVx4_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g530 ( .A(n_311), .Y(n_530) );
INVx2_ASAP7_75t_L g745 ( .A(n_311), .Y(n_745) );
BUFx3_ASAP7_75t_L g821 ( .A(n_311), .Y(n_821) );
AND2x2_ASAP7_75t_L g330 ( .A(n_312), .B(n_331), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_317), .B1(n_318), .B2(n_321), .Y(n_313) );
BUFx3_ASAP7_75t_L g884 ( .A(n_314), .Y(n_884) );
BUFx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g359 ( .A(n_315), .Y(n_359) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_315), .Y(n_366) );
BUFx3_ASAP7_75t_L g590 ( .A(n_315), .Y(n_590) );
A2O1A1Ixp33_ASAP7_75t_L g410 ( .A1(n_317), .A2(n_411), .B(n_412), .C(n_419), .Y(n_410) );
A2O1A1Ixp33_ASAP7_75t_L g326 ( .A1(n_318), .A2(n_327), .B(n_332), .C(n_333), .Y(n_326) );
BUFx3_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx3_ASAP7_75t_L g354 ( .A(n_319), .Y(n_354) );
BUFx3_ASAP7_75t_L g588 ( .A(n_319), .Y(n_588) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_319), .Y(n_714) );
AND2x6_ASAP7_75t_L g885 ( .A(n_319), .B(n_335), .Y(n_885) );
AND2x4_ASAP7_75t_SL g888 ( .A(n_319), .B(n_323), .Y(n_888) );
BUFx3_ASAP7_75t_L g892 ( .A(n_319), .Y(n_892) );
INVx1_ASAP7_75t_L g982 ( .A(n_319), .Y(n_982) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g606 ( .A(n_320), .Y(n_606) );
BUFx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_323), .B(n_421), .Y(n_560) );
AND2x2_ASAP7_75t_L g565 ( .A(n_323), .B(n_330), .Y(n_565) );
AND2x2_ASAP7_75t_L g568 ( .A(n_323), .B(n_569), .Y(n_568) );
AND2x4_ASAP7_75t_L g877 ( .A(n_323), .B(n_569), .Y(n_877) );
AND2x4_ASAP7_75t_L g879 ( .A(n_323), .B(n_366), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_336), .Y(n_325) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_329), .Y(n_364) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx3_ASAP7_75t_L g538 ( .A(n_330), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_330), .B(n_335), .Y(n_556) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NOR2x1_ASAP7_75t_L g1100 ( .A(n_334), .B(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g337 ( .A(n_335), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_335), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_335), .B(n_369), .Y(n_543) );
AOI22xp33_ASAP7_75t_SL g336 ( .A1(n_337), .A2(n_340), .B1(n_341), .B2(n_345), .Y(n_336) );
INVx1_ASAP7_75t_L g899 ( .A(n_337), .Y(n_899) );
BUFx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g549 ( .A(n_339), .Y(n_549) );
INVx1_ASAP7_75t_L g1101 ( .A(n_339), .Y(n_1101) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g550 ( .A(n_342), .B(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g596 ( .A(n_342), .B(n_551), .Y(n_596) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_345), .A2(n_390), .B1(n_391), .B2(n_397), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_357), .B1(n_360), .B2(n_363), .Y(n_346) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g603 ( .A(n_349), .Y(n_603) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_352), .Y(n_569) );
BUFx3_ASAP7_75t_L g716 ( .A(n_352), .Y(n_716) );
INVx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g897 ( .A(n_356), .Y(n_897) );
INVx2_ASAP7_75t_L g1107 ( .A(n_356), .Y(n_1107) );
AND2x4_ASAP7_75t_L g558 ( .A(n_358), .B(n_559), .Y(n_558) );
AOI332xp33_ASAP7_75t_L g815 ( .A1(n_358), .A2(n_559), .A3(n_583), .B1(n_710), .B2(n_711), .B3(n_804), .C1(n_816), .C2(n_817), .Y(n_815) );
INVx3_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx4_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x4_ASAP7_75t_L g525 ( .A(n_362), .B(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_SL g754 ( .A(n_362), .B(n_384), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_362), .B(n_526), .Y(n_824) );
INVx4_ASAP7_75t_L g881 ( .A(n_362), .Y(n_881) );
BUFx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g601 ( .A(n_366), .Y(n_601) );
INVx1_ASAP7_75t_L g511 ( .A(n_367), .Y(n_511) );
BUFx2_ASAP7_75t_L g780 ( .A(n_367), .Y(n_780) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g451 ( .A(n_368), .B(n_452), .Y(n_451) );
AND2x4_ASAP7_75t_L g514 ( .A(n_368), .B(n_515), .Y(n_514) );
BUFx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g608 ( .A(n_369), .Y(n_608) );
NAND3xp33_ASAP7_75t_SL g370 ( .A(n_371), .B(n_389), .C(n_404), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_373), .A2(n_872), .B1(n_875), .B2(n_903), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_373), .A2(n_903), .B1(n_1067), .B2(n_1068), .Y(n_1066) );
AND2x4_ASAP7_75t_L g373 ( .A(n_374), .B(n_382), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx8_ASAP7_75t_L g411 ( .A(n_375), .Y(n_411) );
INVx3_ASAP7_75t_L g475 ( .A(n_375), .Y(n_475) );
INVx2_ASAP7_75t_L g863 ( .A(n_375), .Y(n_863) );
INVx8_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2x1p5_ASAP7_75t_L g644 ( .A(n_376), .B(n_422), .Y(n_644) );
BUFx3_ASAP7_75t_L g672 ( .A(n_376), .Y(n_672) );
AND2x2_ASAP7_75t_L g676 ( .A(n_376), .B(n_677), .Y(n_676) );
BUFx3_ASAP7_75t_L g772 ( .A(n_376), .Y(n_772) );
AND2x4_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
AND2x4_ASAP7_75t_L g394 ( .A(n_377), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_378), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_378), .B(n_402), .Y(n_409) );
OR2x2_ASAP7_75t_L g432 ( .A(n_378), .B(n_380), .Y(n_432) );
AND2x4_ASAP7_75t_L g468 ( .A(n_378), .B(n_417), .Y(n_468) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVxp67_ASAP7_75t_L g395 ( .A(n_381), .Y(n_395) );
AND2x4_ASAP7_75t_L g903 ( .A(n_382), .B(n_633), .Y(n_903) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g396 ( .A(n_383), .Y(n_396) );
OR2x2_ASAP7_75t_L g398 ( .A(n_383), .B(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g406 ( .A(n_383), .B(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_387), .Y(n_383) );
OR2x2_ASAP7_75t_L g428 ( .A(n_384), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g527 ( .A(n_384), .Y(n_527) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx2_ASAP7_75t_L g551 ( .A(n_385), .Y(n_551) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g461 ( .A(n_387), .Y(n_461) );
INVx1_ASAP7_75t_L g677 ( .A(n_387), .Y(n_677) );
INVx3_ASAP7_75t_L g423 ( .A(n_388), .Y(n_423) );
NAND2xp33_ASAP7_75t_SL g429 ( .A(n_388), .B(n_425), .Y(n_429) );
BUFx3_ASAP7_75t_L g509 ( .A(n_388), .Y(n_509) );
AND2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_396), .Y(n_391) );
INVx2_ASAP7_75t_L g445 ( .A(n_392), .Y(n_445) );
INVx2_ASAP7_75t_L g806 ( .A(n_392), .Y(n_806) );
INVx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x6_ASAP7_75t_SL g658 ( .A(n_393), .B(n_659), .Y(n_658) );
BUFx2_ASAP7_75t_L g853 ( .A(n_393), .Y(n_853) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_394), .Y(n_439) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_394), .Y(n_506) );
BUFx8_ASAP7_75t_L g633 ( .A(n_394), .Y(n_633) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g901 ( .A(n_398), .B(n_596), .Y(n_901) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_399), .Y(n_435) );
INVx4_ASAP7_75t_L g489 ( .A(n_399), .Y(n_489) );
INVx3_ASAP7_75t_L g766 ( .A(n_399), .Y(n_766) );
OAI221xp5_ASAP7_75t_L g790 ( .A1(n_399), .A2(n_508), .B1(n_791), .B2(n_792), .C(n_793), .Y(n_790) );
HB1xp67_ASAP7_75t_L g1436 ( .A(n_399), .Y(n_1436) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx3_ASAP7_75t_L g418 ( .A(n_400), .Y(n_418) );
BUFx2_ASAP7_75t_L g620 ( .A(n_400), .Y(n_620) );
NAND2x1p5_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g417 ( .A(n_402), .Y(n_417) );
INVx2_ASAP7_75t_L g413 ( .A(n_403), .Y(n_413) );
AND2x4_ASAP7_75t_L g464 ( .A(n_403), .B(n_416), .Y(n_464) );
NOR2xp33_ASAP7_75t_SL g404 ( .A(n_405), .B(n_426), .Y(n_404) );
AND2x4_ASAP7_75t_L g839 ( .A(n_406), .B(n_555), .Y(n_839) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_408), .Y(n_638) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx2_ASAP7_75t_L g442 ( .A(n_409), .Y(n_442) );
INVx3_ASAP7_75t_L g617 ( .A(n_413), .Y(n_617) );
INVx2_ASAP7_75t_L g847 ( .A(n_414), .Y(n_847) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g614 ( .A(n_415), .B(n_422), .Y(n_614) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g448 ( .A1(n_418), .A2(n_431), .B1(n_449), .B2(n_450), .Y(n_448) );
OAI221xp5_ASAP7_75t_L g773 ( .A1(n_418), .A2(n_445), .B1(n_508), .B2(n_741), .C(n_746), .Y(n_773) );
OAI221xp5_ASAP7_75t_L g775 ( .A1(n_418), .A2(n_471), .B1(n_492), .B2(n_734), .C(n_747), .Y(n_775) );
OAI221xp5_ASAP7_75t_L g1030 ( .A1(n_418), .A2(n_471), .B1(n_492), .B2(n_1031), .C(n_1032), .Y(n_1030) );
OAI221xp5_ASAP7_75t_L g1165 ( .A1(n_418), .A2(n_472), .B1(n_508), .B2(n_1166), .C(n_1167), .Y(n_1165) );
OAI221xp5_ASAP7_75t_L g1170 ( .A1(n_418), .A2(n_431), .B1(n_492), .B2(n_1171), .C(n_1172), .Y(n_1170) );
AND2x2_ASAP7_75t_L g844 ( .A(n_419), .B(n_617), .Y(n_844) );
AND2x4_ASAP7_75t_L g846 ( .A(n_419), .B(n_847), .Y(n_846) );
AND2x4_ASAP7_75t_L g849 ( .A(n_419), .B(n_640), .Y(n_849) );
AND2x4_ASAP7_75t_L g419 ( .A(n_420), .B(n_422), .Y(n_419) );
OR2x2_ASAP7_75t_L g555 ( .A(n_420), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g710 ( .A(n_420), .Y(n_710) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g859 ( .A(n_421), .Y(n_859) );
INVx1_ASAP7_75t_L g478 ( .A(n_422), .Y(n_478) );
AND2x6_ASAP7_75t_L g616 ( .A(n_422), .B(n_617), .Y(n_616) );
AND2x4_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
NAND2x1p5_ASAP7_75t_L g452 ( .A(n_423), .B(n_453), .Y(n_452) );
NAND3x1_ASAP7_75t_L g858 ( .A(n_423), .B(n_453), .C(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g508 ( .A(n_425), .B(n_509), .Y(n_508) );
AND3x4_ASAP7_75t_L g866 ( .A(n_425), .B(n_509), .C(n_608), .Y(n_866) );
OAI33xp33_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_430), .A3(n_436), .B1(n_444), .B2(n_448), .B3(n_451), .Y(n_426) );
BUFx4f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx2_ASAP7_75t_L g627 ( .A(n_429), .Y(n_627) );
OAI22xp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_433), .B1(n_434), .B2(n_435), .Y(n_430) );
OAI221xp5_ASAP7_75t_L g795 ( .A1(n_431), .A2(n_492), .B1(n_620), .B2(n_796), .C(n_797), .Y(n_795) );
INVx1_ASAP7_75t_L g947 ( .A(n_431), .Y(n_947) );
BUFx4f_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx3_ASAP7_75t_L g471 ( .A(n_432), .Y(n_471) );
BUFx3_ASAP7_75t_L g490 ( .A(n_432), .Y(n_490) );
INVx2_ASAP7_75t_L g497 ( .A(n_432), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B1(n_440), .B2(n_443), .Y(n_436) );
INVx8_ASAP7_75t_L g626 ( .A(n_438), .Y(n_626) );
OAI221xp5_ASAP7_75t_L g1123 ( .A1(n_438), .A2(n_1124), .B1(n_1125), .B2(n_1126), .C(n_1127), .Y(n_1123) );
INVx5_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_SL g472 ( .A(n_439), .Y(n_472) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_439), .Y(n_483) );
INVx3_ASAP7_75t_L g799 ( .A(n_439), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_440), .A2(n_445), .B1(n_446), .B2(n_447), .Y(n_444) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx2_ASAP7_75t_L g500 ( .A(n_441), .Y(n_500) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx3_ASAP7_75t_L g485 ( .A(n_442), .Y(n_485) );
INVx3_ASAP7_75t_L g492 ( .A(n_452), .Y(n_492) );
NAND4xp75_ASAP7_75t_L g455 ( .A(n_456), .B(n_512), .C(n_552), .D(n_562), .Y(n_455) );
OAI21x1_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_479), .B(n_510), .Y(n_456) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_462), .B(n_473), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_459), .A2(n_581), .B1(n_635), .B2(n_641), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g763 ( .A1(n_459), .A2(n_643), .B1(n_758), .B2(n_764), .C(n_767), .Y(n_763) );
AOI221xp5_ASAP7_75t_L g803 ( .A1(n_459), .A2(n_643), .B1(n_804), .B2(n_805), .C(n_810), .Y(n_803) );
BUFx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g659 ( .A(n_461), .Y(n_659) );
AND2x4_ASAP7_75t_L g661 ( .A(n_461), .B(n_464), .Y(n_661) );
AOI221xp5_ASAP7_75t_SL g462 ( .A1(n_463), .A2(n_465), .B1(n_466), .B2(n_469), .C(n_470), .Y(n_462) );
BUFx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx12f_ASAP7_75t_L g623 ( .A(n_464), .Y(n_623) );
INVx5_ASAP7_75t_L g669 ( .A(n_464), .Y(n_669) );
BUFx3_ASAP7_75t_L g861 ( .A(n_464), .Y(n_861) );
BUFx2_ASAP7_75t_L g941 ( .A(n_464), .Y(n_941) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g854 ( .A(n_467), .Y(n_854) );
INVx2_ASAP7_75t_L g999 ( .A(n_467), .Y(n_999) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx3_ASAP7_75t_L g625 ( .A(n_468), .Y(n_625) );
BUFx2_ASAP7_75t_L g640 ( .A(n_468), .Y(n_640) );
AND2x2_ASAP7_75t_L g679 ( .A(n_468), .B(n_677), .Y(n_679) );
BUFx2_ASAP7_75t_L g1128 ( .A(n_468), .Y(n_1128) );
INVx1_ASAP7_75t_L g1444 ( .A(n_471), .Y(n_1444) );
A2O1A1Ixp33_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B(n_476), .C(n_477), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_475), .A2(n_577), .B1(n_597), .B2(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OR2x6_ASAP7_75t_L g619 ( .A(n_478), .B(n_620), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_486), .B1(n_493), .B2(n_501), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B1(n_484), .B2(n_485), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_481), .A2(n_494), .B1(n_518), .B2(n_520), .Y(n_517) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI221xp5_ASAP7_75t_L g528 ( .A1(n_484), .A2(n_502), .B1(n_529), .B2(n_531), .C(n_536), .Y(n_528) );
OAI221xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_488), .B1(n_490), .B2(n_491), .C(n_492), .Y(n_486) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g503 ( .A(n_489), .Y(n_503) );
INVx2_ASAP7_75t_L g667 ( .A(n_489), .Y(n_667) );
INVx2_ASAP7_75t_L g944 ( .A(n_489), .Y(n_944) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_490), .A2(n_1023), .B1(n_1024), .B2(n_1025), .Y(n_1022) );
INVx3_ASAP7_75t_L g629 ( .A(n_492), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_492), .B(n_685), .Y(n_684) );
OAI221xp5_ASAP7_75t_L g942 ( .A1(n_492), .A2(n_943), .B1(n_944), .B2(n_945), .C(n_946), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g1445 ( .A(n_492), .B(n_1446), .Y(n_1445) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B1(n_498), .B2(n_499), .Y(n_493) );
BUFx4f_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OAI221xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_503), .B1(n_504), .B2(n_507), .C(n_508), .Y(n_501) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g636 ( .A(n_506), .Y(n_636) );
INVx1_ASAP7_75t_L g665 ( .A(n_506), .Y(n_665) );
INVx2_ASAP7_75t_L g793 ( .A(n_506), .Y(n_793) );
BUFx6f_ASAP7_75t_L g940 ( .A(n_506), .Y(n_940) );
INVx2_ASAP7_75t_L g1029 ( .A(n_506), .Y(n_1029) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_508), .A2(n_669), .B1(n_670), .B2(n_671), .C(n_673), .Y(n_668) );
OAI221xp5_ASAP7_75t_L g949 ( .A1(n_508), .A2(n_925), .B1(n_944), .B2(n_950), .C(n_951), .Y(n_949) );
OAI21xp33_ASAP7_75t_L g1020 ( .A1(n_508), .A2(n_632), .B(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g1438 ( .A(n_508), .Y(n_1438) );
OAI31xp33_ASAP7_75t_L g993 ( .A1(n_510), .A2(n_994), .A3(n_995), .B(n_1008), .Y(n_993) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AOI211x1_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_516), .B(n_523), .C(n_544), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AOI31xp33_ASAP7_75t_L g586 ( .A1(n_514), .A2(n_587), .A3(n_589), .B(n_591), .Y(n_586) );
INVx2_ASAP7_75t_L g707 ( .A(n_514), .Y(n_707) );
INVx2_ASAP7_75t_L g731 ( .A(n_514), .Y(n_731) );
INVx4_ASAP7_75t_L g929 ( .A(n_514), .Y(n_929) );
INVx2_ASAP7_75t_L g979 ( .A(n_514), .Y(n_979) );
AOI222xp33_ASAP7_75t_L g1183 ( .A1(n_514), .A2(n_525), .B1(n_709), .B2(n_1184), .C1(n_1185), .C2(n_1192), .Y(n_1183) );
BUFx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx3_ASAP7_75t_L g718 ( .A(n_519), .Y(n_718) );
BUFx6f_ASAP7_75t_L g921 ( .A(n_519), .Y(n_921) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_520), .A2(n_743), .B1(n_746), .B2(n_747), .Y(n_742) );
BUFx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OR2x2_ASAP7_75t_L g561 ( .A(n_521), .B(n_560), .Y(n_561) );
OR2x2_ASAP7_75t_L g584 ( .A(n_521), .B(n_560), .Y(n_584) );
BUFx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_522), .Y(n_540) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_528), .B(n_539), .Y(n_523) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
NAND3xp33_ASAP7_75t_L g598 ( .A(n_525), .B(n_599), .C(n_602), .Y(n_598) );
AOI322xp5_ASAP7_75t_L g697 ( .A1(n_525), .A2(n_698), .A3(n_701), .B1(n_706), .B2(n_708), .C1(n_709), .C2(n_712), .Y(n_697) );
AOI322xp5_ASAP7_75t_L g974 ( .A1(n_525), .A2(n_583), .A3(n_975), .B1(n_976), .B2(n_977), .C1(n_980), .C2(n_988), .Y(n_974) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OAI221xp5_ASAP7_75t_L g1102 ( .A1(n_531), .A2(n_1103), .B1(n_1104), .B2(n_1105), .C(n_1106), .Y(n_1102) );
INVx6_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx5_ASAP7_75t_L g705 ( .A(n_532), .Y(n_705) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g720 ( .A(n_533), .Y(n_720) );
INVx2_ASAP7_75t_SL g735 ( .A(n_533), .Y(n_735) );
INVx4_ASAP7_75t_L g914 ( .A(n_533), .Y(n_914) );
INVx2_ASAP7_75t_L g928 ( .A(n_533), .Y(n_928) );
INVx8_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g883 ( .A(n_538), .Y(n_883) );
INVx1_ASAP7_75t_L g890 ( .A(n_538), .Y(n_890) );
INVx2_ASAP7_75t_SL g1089 ( .A(n_538), .Y(n_1089) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_539), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g1149 ( .A1(n_539), .A2(n_1150), .B(n_1151), .Y(n_1149) );
OR2x6_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
INVx4_ASAP7_75t_L g739 ( .A(n_540), .Y(n_739) );
BUFx4f_ASAP7_75t_L g822 ( .A(n_540), .Y(n_822) );
BUFx6f_ASAP7_75t_L g827 ( .A(n_540), .Y(n_827) );
BUFx4f_ASAP7_75t_L g1044 ( .A(n_540), .Y(n_1044) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2x2_ASAP7_75t_L g547 ( .A(n_542), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g593 ( .A(n_547), .Y(n_593) );
HB1xp67_ASAP7_75t_L g1141 ( .A(n_547), .Y(n_1141) );
INVx2_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g564 ( .A(n_551), .Y(n_564) );
INVxp67_ASAP7_75t_L g836 ( .A(n_551), .Y(n_836) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g711 ( .A(n_556), .Y(n_711) );
INVxp67_ASAP7_75t_L g1451 ( .A(n_557), .Y(n_1451) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_558), .A2(n_581), .B1(n_582), .B2(n_583), .Y(n_580) );
AOI222xp33_ASAP7_75t_L g756 ( .A1(n_558), .A2(n_583), .B1(n_709), .B2(n_757), .C1(n_758), .C2(n_759), .Y(n_756) );
AOI222xp33_ASAP7_75t_L g930 ( .A1(n_558), .A2(n_583), .B1(n_709), .B2(n_931), .C1(n_932), .C2(n_933), .Y(n_930) );
AOI222xp33_ASAP7_75t_L g970 ( .A1(n_558), .A2(n_593), .B1(n_595), .B2(n_971), .C1(n_972), .C2(n_973), .Y(n_970) );
AOI222xp33_ASAP7_75t_L g1035 ( .A1(n_558), .A2(n_583), .B1(n_709), .B2(n_1015), .C1(n_1036), .C2(n_1037), .Y(n_1035) );
AOI222xp33_ASAP7_75t_L g1137 ( .A1(n_558), .A2(n_583), .B1(n_709), .B2(n_1118), .C1(n_1121), .C2(n_1138), .Y(n_1137) );
AOI222xp33_ASAP7_75t_L g1180 ( .A1(n_558), .A2(n_593), .B1(n_595), .B2(n_1174), .C1(n_1181), .C2(n_1182), .Y(n_1180) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AOI22xp33_ASAP7_75t_SL g562 ( .A1(n_563), .A2(n_566), .B1(n_567), .B2(n_570), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_563), .B(n_577), .Y(n_576) );
AOI211xp5_ASAP7_75t_L g690 ( .A1(n_563), .A2(n_691), .B(n_692), .C(n_696), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_563), .B(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_563), .B(n_809), .Y(n_813) );
INVx3_ASAP7_75t_L g907 ( .A(n_563), .Y(n_907) );
AOI211x1_ASAP7_75t_L g967 ( .A1(n_563), .A2(n_968), .B(n_969), .C(n_991), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_563), .A2(n_1116), .B1(n_1135), .B2(n_1156), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_563), .B(n_1198), .Y(n_1197) );
AO211x2_ASAP7_75t_L g1421 ( .A1(n_563), .A2(n_1422), .B(n_1423), .C(n_1449), .Y(n_1421) );
AND2x4_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AND2x4_ASAP7_75t_L g567 ( .A(n_564), .B(n_568), .Y(n_567) );
BUFx6f_ASAP7_75t_L g874 ( .A(n_565), .Y(n_874) );
INVx1_ASAP7_75t_L g1092 ( .A(n_565), .Y(n_1092) );
INVx1_ASAP7_75t_L g646 ( .A(n_567), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_567), .B(n_688), .Y(n_687) );
NAND2xp33_ASAP7_75t_SL g781 ( .A(n_567), .B(n_782), .Y(n_781) );
HB1xp67_ASAP7_75t_L g958 ( .A(n_567), .Y(n_958) );
INVx1_ASAP7_75t_L g992 ( .A(n_567), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_567), .B(n_1039), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1447 ( .A(n_567), .B(n_1448), .Y(n_1447) );
BUFx6f_ASAP7_75t_L g700 ( .A(n_569), .Y(n_700) );
INVx2_ASAP7_75t_L g896 ( .A(n_569), .Y(n_896) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_649), .B1(n_650), .B2(n_721), .Y(n_571) );
INVx1_ASAP7_75t_L g721 ( .A(n_572), .Y(n_721) );
OAI21x1_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_574), .B(n_648), .Y(n_572) );
NAND4xp25_ASAP7_75t_L g648 ( .A(n_573), .B(n_576), .C(n_578), .D(n_607), .Y(n_648) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND3xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .C(n_607), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_579), .B(n_585), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g1199 ( .A1(n_583), .A2(n_591), .B(n_1200), .Y(n_1199) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND3xp33_ASAP7_75t_SL g585 ( .A(n_586), .B(n_592), .C(n_598), .Y(n_585) );
NOR3xp33_ASAP7_75t_L g818 ( .A(n_591), .B(n_819), .C(n_829), .Y(n_818) );
NOR3xp33_ASAP7_75t_L g908 ( .A(n_591), .B(n_909), .C(n_910), .Y(n_908) );
AOI21xp33_ASAP7_75t_L g989 ( .A1(n_591), .A2(n_709), .B(n_990), .Y(n_989) );
OR3x1_ASAP7_75t_L g1040 ( .A(n_591), .B(n_1041), .C(n_1042), .Y(n_1040) );
AOI21xp33_ASAP7_75t_L g1468 ( .A1(n_591), .A2(n_709), .B(n_1469), .Y(n_1468) );
AOI22xp33_ASAP7_75t_SL g592 ( .A1(n_593), .A2(n_594), .B1(n_595), .B2(n_597), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_593), .A2(n_595), .B1(n_694), .B2(n_695), .Y(n_693) );
AOI222xp33_ASAP7_75t_L g1450 ( .A1(n_593), .A2(n_595), .B1(n_1425), .B2(n_1451), .C1(n_1452), .C2(n_1453), .Y(n_1450) );
INVx2_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g1087 ( .A(n_605), .Y(n_1087) );
INVx1_ASAP7_75t_L g1146 ( .A(n_605), .Y(n_1146) );
BUFx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_608), .A2(n_609), .B1(n_645), .B2(n_647), .Y(n_607) );
INVx2_ASAP7_75t_SL g686 ( .A(n_608), .Y(n_686) );
INVx1_ASAP7_75t_L g812 ( .A(n_608), .Y(n_812) );
NAND3xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_621), .C(n_634), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_618), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g656 ( .A(n_614), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_614), .A2(n_616), .B1(n_972), .B2(n_988), .Y(n_1009) );
AOI221xp5_ASAP7_75t_L g1119 ( .A1(n_614), .A2(n_616), .B1(n_618), .B2(n_1120), .C(n_1121), .Y(n_1119) );
INVx4_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NOR3xp33_ASAP7_75t_L g768 ( .A(n_618), .B(n_769), .C(n_774), .Y(n_768) );
NOR3xp33_ASAP7_75t_L g788 ( .A(n_618), .B(n_789), .C(n_794), .Y(n_788) );
CKINVDCx5p33_ASAP7_75t_R g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g683 ( .A(n_620), .Y(n_683) );
INVx1_ASAP7_75t_L g1003 ( .A(n_620), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B1(n_628), .B2(n_630), .Y(n_621) );
BUFx2_ASAP7_75t_L g868 ( .A(n_623), .Y(n_868) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx3_ASAP7_75t_L g777 ( .A(n_633), .Y(n_777) );
INVx2_ASAP7_75t_SL g951 ( .A(n_633), .Y(n_951) );
OAI221xp5_ASAP7_75t_L g996 ( .A1(n_637), .A2(n_806), .B1(n_987), .B2(n_997), .C(n_998), .Y(n_996) );
CKINVDCx8_ASAP7_75t_R g637 ( .A(n_638), .Y(n_637) );
INVx3_ASAP7_75t_L g778 ( .A(n_638), .Y(n_778) );
INVx3_ASAP7_75t_L g801 ( .A(n_638), .Y(n_801) );
INVx1_ASAP7_75t_L g1024 ( .A(n_638), .Y(n_1024) );
INVx3_ASAP7_75t_L g1125 ( .A(n_638), .Y(n_1125) );
BUFx2_ASAP7_75t_L g1078 ( .A(n_640), .Y(n_1078) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI211xp5_ASAP7_75t_SL g653 ( .A1(n_643), .A2(n_654), .B(n_655), .C(n_657), .Y(n_653) );
AOI211xp5_ASAP7_75t_SL g935 ( .A1(n_643), .A2(n_931), .B(n_936), .C(n_937), .Y(n_935) );
AOI211xp5_ASAP7_75t_L g1014 ( .A1(n_643), .A2(n_1015), .B(n_1016), .C(n_1017), .Y(n_1014) );
AOI211xp5_ASAP7_75t_SL g1173 ( .A1(n_643), .A2(n_1174), .B(n_1175), .C(n_1176), .Y(n_1173) );
AOI211xp5_ASAP7_75t_SL g1424 ( .A1(n_643), .A2(n_1425), .B(n_1426), .C(n_1427), .Y(n_1424) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OR2x6_ASAP7_75t_L g835 ( .A(n_644), .B(n_836), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_645), .B(n_1178), .Y(n_1177) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NOR2x1_ASAP7_75t_L g651 ( .A(n_652), .B(n_689), .Y(n_651) );
A2O1A1Ixp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_662), .B(n_686), .C(n_687), .Y(n_652) );
CKINVDCx5p33_ASAP7_75t_R g1117 ( .A(n_658), .Y(n_1117) );
INVx3_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_661), .A2(n_1116), .B1(n_1117), .B2(n_1118), .Y(n_1115) );
NOR3xp33_ASAP7_75t_SL g662 ( .A(n_663), .B(n_674), .C(n_680), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g1072 ( .A(n_669), .Y(n_1072) );
INVx2_ASAP7_75t_L g1075 ( .A(n_669), .Y(n_1075) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_670), .A2(n_718), .B1(n_719), .B2(n_720), .Y(n_717) );
INVx2_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_672), .B(n_809), .Y(n_808) );
BUFx3_ASAP7_75t_L g1006 ( .A(n_672), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_673), .A2(n_703), .B1(n_704), .B2(n_705), .Y(n_702) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_676), .A2(n_679), .B1(n_968), .B2(n_973), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_676), .A2(n_679), .B1(n_1135), .B2(n_1136), .Y(n_1134) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_697), .Y(n_689) );
BUFx3_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_703), .A2(n_733), .B1(n_734), .B2(n_735), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g1463 ( .A1(n_703), .A2(n_705), .B1(n_1464), .B2(n_1465), .Y(n_1463) );
OAI33xp33_ASAP7_75t_L g1042 ( .A1(n_707), .A2(n_753), .A3(n_1043), .B1(n_1046), .B2(n_1049), .B3(n_1052), .Y(n_1042) );
AND2x4_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
BUFx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
BUFx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g1145 ( .A(n_716), .Y(n_1145) );
INVx1_ASAP7_75t_L g1188 ( .A(n_716), .Y(n_1188) );
OAI22xp5_ASAP7_75t_L g1052 ( .A1(n_718), .A2(n_735), .B1(n_1025), .B2(n_1053), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_720), .A2(n_1023), .B1(n_1032), .B2(n_1047), .Y(n_1046) );
XNOR2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_830), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
XNOR2x1_ASAP7_75t_L g724 ( .A(n_725), .B(n_783), .Y(n_724) );
XNOR2x1_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_728), .B(n_762), .Y(n_727) );
NAND3xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_756), .C(n_760), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_755), .Y(n_729) );
OAI33xp33_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_732), .A3(n_736), .B1(n_742), .B2(n_748), .B3(n_753), .Y(n_730) );
OAI22xp5_ASAP7_75t_SL g819 ( .A1(n_731), .A2(n_820), .B1(n_824), .B2(n_825), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_735), .A2(n_749), .B1(n_751), .B2(n_752), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g1193 ( .A1(n_735), .A2(n_1194), .B1(n_1195), .B2(n_1196), .Y(n_1193) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_738), .B1(n_740), .B2(n_741), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_737), .A2(n_752), .B1(n_777), .B2(n_778), .Y(n_776) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g919 ( .A(n_739), .Y(n_919) );
INVx1_ASAP7_75t_L g1051 ( .A(n_739), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g1049 ( .A1(n_743), .A2(n_1031), .B1(n_1050), .B2(n_1051), .Y(n_1049) );
INVx4_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
BUFx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g826 ( .A(n_745), .Y(n_826) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
A2O1A1Ixp33_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_768), .B(n_779), .C(n_781), .Y(n_762) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g807 ( .A(n_766), .Y(n_807) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
BUFx2_ASAP7_75t_L g1133 ( .A(n_772), .Y(n_1133) );
INVx1_ASAP7_75t_L g1074 ( .A(n_777), .Y(n_1074) );
AOI21xp5_ASAP7_75t_L g869 ( .A1(n_779), .A2(n_870), .B(n_900), .Y(n_869) );
INVx1_ASAP7_75t_L g1033 ( .A(n_779), .Y(n_1033) );
A2O1A1Ixp33_ASAP7_75t_L g1161 ( .A1(n_779), .A2(n_1162), .B(n_1173), .C(n_1177), .Y(n_1161) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g1113 ( .A1(n_780), .A2(n_1114), .B(n_1122), .Y(n_1113) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
XNOR2x1_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
OR2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_814), .Y(n_786) );
A2O1A1Ixp33_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_803), .B(n_811), .C(n_813), .Y(n_787) );
OAI221xp5_ASAP7_75t_L g825 ( .A1(n_791), .A2(n_796), .B1(n_826), .B2(n_827), .C(n_828), .Y(n_825) );
OAI221xp5_ASAP7_75t_L g820 ( .A1(n_792), .A2(n_800), .B1(n_821), .B2(n_822), .C(n_823), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_800), .B1(n_801), .B2(n_802), .Y(n_798) );
OAI211xp5_ASAP7_75t_L g1129 ( .A1(n_807), .A2(n_1130), .B(n_1131), .C(n_1132), .Y(n_1129) );
A2O1A1Ixp33_ASAP7_75t_SL g1423 ( .A1(n_811), .A2(n_1424), .B(n_1428), .C(n_1447), .Y(n_1423) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
BUFx2_ASAP7_75t_L g955 ( .A(n_812), .Y(n_955) );
INVx2_ASAP7_75t_L g916 ( .A(n_821), .Y(n_916) );
OAI221xp5_ASAP7_75t_L g922 ( .A1(n_822), .A2(n_923), .B1(n_924), .B2(n_925), .C(n_926), .Y(n_922) );
INVx1_ASAP7_75t_L g1147 ( .A(n_824), .Y(n_1147) );
OAI22xp5_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_904), .B1(n_960), .B2(n_961), .Y(n_830) );
INVx1_ASAP7_75t_L g961 ( .A(n_831), .Y(n_961) );
NAND2xp67_ASAP7_75t_L g832 ( .A(n_833), .B(n_869), .Y(n_832) );
AOI221xp5_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_837), .B1(n_838), .B2(n_840), .C(n_841), .Y(n_833) );
INVx3_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
AOI221xp5_ASAP7_75t_L g878 ( .A1(n_837), .A2(n_879), .B1(n_880), .B2(n_882), .C(n_885), .Y(n_878) );
INVx8_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
NAND3xp33_ASAP7_75t_SL g841 ( .A(n_842), .B(n_848), .C(n_850), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_844), .B1(n_845), .B2(n_846), .Y(n_842) );
AOI222xp33_ASAP7_75t_L g886 ( .A1(n_843), .A2(n_845), .B1(n_887), .B2(n_889), .C1(n_891), .C2(n_898), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_844), .A2(n_846), .B1(n_1064), .B2(n_1065), .Y(n_1063) );
INVx3_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
NOR3xp33_ASAP7_75t_L g1061 ( .A(n_849), .B(n_1062), .C(n_1079), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_851), .A2(n_855), .B1(n_862), .B2(n_867), .Y(n_850) );
INVx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
AND2x2_ASAP7_75t_L g855 ( .A(n_856), .B(n_860), .Y(n_855) );
BUFx2_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx3_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx3_ASAP7_75t_L g1076 ( .A(n_858), .Y(n_1076) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
AOI33xp33_ASAP7_75t_L g1069 ( .A1(n_865), .A2(n_1070), .A3(n_1071), .B1(n_1073), .B2(n_1076), .B3(n_1077), .Y(n_1069) );
BUFx3_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
NAND3xp33_ASAP7_75t_SL g870 ( .A(n_871), .B(n_878), .C(n_886), .Y(n_870) );
AOI22xp5_ASAP7_75t_L g871 ( .A1(n_872), .A2(n_873), .B1(n_875), .B2(n_876), .Y(n_871) );
HB1xp67_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
BUFx6f_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g1094 ( .A(n_877), .Y(n_1094) );
INVx3_ASAP7_75t_L g1082 ( .A(n_879), .Y(n_1082) );
AOI21xp5_ASAP7_75t_SL g1083 ( .A1(n_885), .A2(n_1084), .B(n_1088), .Y(n_1083) );
BUFx3_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx2_ASAP7_75t_L g1098 ( .A(n_888), .Y(n_1098) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
HB1xp67_ASAP7_75t_L g1462 ( .A(n_895), .Y(n_1462) );
INVx2_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g960 ( .A(n_904), .Y(n_960) );
XOR2x2_ASAP7_75t_L g904 ( .A(n_905), .B(n_959), .Y(n_904) );
NOR2x1_ASAP7_75t_SL g905 ( .A(n_906), .B(n_934), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_911), .B(n_922), .Y(n_910) );
OAI211xp5_ASAP7_75t_L g911 ( .A1(n_912), .A2(n_913), .B(n_915), .C(n_917), .Y(n_911) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g983 ( .A1(n_914), .A2(n_984), .B1(n_985), .B2(n_987), .Y(n_983) );
OAI22xp5_ASAP7_75t_L g1189 ( .A1(n_914), .A2(n_1172), .B1(n_1190), .B2(n_1191), .Y(n_1189) );
INVx3_ASAP7_75t_L g924 ( .A(n_916), .Y(n_924) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
OAI221xp5_ASAP7_75t_L g1151 ( .A1(n_919), .A2(n_1124), .B1(n_1152), .B2(n_1153), .C(n_1154), .Y(n_1151) );
INVx2_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVxp33_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx2_ASAP7_75t_SL g1459 ( .A(n_929), .Y(n_1459) );
A2O1A1Ixp33_ASAP7_75t_SL g934 ( .A1(n_935), .A2(n_938), .B(n_953), .C(n_956), .Y(n_934) );
NOR3xp33_ASAP7_75t_L g938 ( .A(n_939), .B(n_948), .C(n_952), .Y(n_938) );
INVx1_ASAP7_75t_L g1432 ( .A(n_940), .Y(n_1432) );
INVx2_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g1169 ( .A(n_951), .Y(n_1169) );
OAI21xp5_ASAP7_75t_L g1080 ( .A1(n_953), .A2(n_1081), .B(n_1095), .Y(n_1080) );
INVx2_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_957), .B(n_958), .Y(n_956) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
XNOR2xp5_ASAP7_75t_L g963 ( .A(n_964), .B(n_1109), .Y(n_963) );
AOI22xp5_ASAP7_75t_L g964 ( .A1(n_965), .A2(n_1056), .B1(n_1057), .B2(n_1108), .Y(n_964) );
INVx1_ASAP7_75t_L g1108 ( .A(n_965), .Y(n_1108) );
AOI22xp5_ASAP7_75t_L g965 ( .A1(n_966), .A2(n_1011), .B1(n_1054), .B2(n_1055), .Y(n_965) );
INVx1_ASAP7_75t_L g1054 ( .A(n_966), .Y(n_1054) );
XOR2x2_ASAP7_75t_L g966 ( .A(n_967), .B(n_1010), .Y(n_966) );
NAND3xp33_ASAP7_75t_L g969 ( .A(n_970), .B(n_974), .C(n_989), .Y(n_969) );
INVx1_ASAP7_75t_L g1150 ( .A(n_977), .Y(n_1150) );
INVx1_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
BUFx6f_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
INVx1_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g1186 ( .A(n_982), .Y(n_1186) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g1195 ( .A(n_986), .Y(n_1195) );
INVx1_ASAP7_75t_L g1156 ( .A(n_992), .Y(n_1156) );
NAND3xp33_ASAP7_75t_L g995 ( .A(n_996), .B(n_1000), .C(n_1007), .Y(n_995) );
OAI211xp5_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1002), .B(n_1004), .C(n_1005), .Y(n_1000) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
INVx2_ASAP7_75t_L g1055 ( .A(n_1011), .Y(n_1055) );
AOI211x1_ASAP7_75t_L g1012 ( .A1(n_1013), .A2(n_1033), .B(n_1034), .C(n_1040), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1018), .Y(n_1013) );
NOR3xp33_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1026), .C(n_1027), .Y(n_1018) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
INVx3_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
INVx2_ASAP7_75t_L g1103 ( .A(n_1048), .Y(n_1103) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
HB1xp67_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1080), .Y(n_1060) );
NAND3xp33_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1066), .C(n_1069), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_1067), .A2(n_1068), .B1(n_1091), .B2(n_1093), .Y(n_1090) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
INVx2_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
INVx4_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
INVx2_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
XOR2x2_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1159), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1112), .Y(n_1157) );
NAND4xp25_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1137), .C(n_1139), .D(n_1155), .Y(n_1112) );
NAND3xp33_ASAP7_75t_L g1122 ( .A(n_1123), .B(n_1129), .C(n_1134), .Y(n_1122) );
NOR2xp33_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1149), .Y(n_1139) );
NAND3xp33_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1147), .C(n_1148), .Y(n_1142) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
OR2x2_ASAP7_75t_L g1160 ( .A(n_1161), .B(n_1179), .Y(n_1160) );
NOR3xp33_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1164), .C(n_1168), .Y(n_1162) );
NAND4xp25_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1183), .C(n_1197), .D(n_1199), .Y(n_1179) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
OAI221xp5_ASAP7_75t_L g1202 ( .A1(n_1203), .A2(n_1416), .B1(n_1419), .B2(n_1470), .C(n_1474), .Y(n_1202) );
AND3x1_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1353), .C(n_1390), .Y(n_1203) );
AOI211xp5_ASAP7_75t_SL g1204 ( .A1(n_1205), .A2(n_1226), .B(n_1280), .C(n_1329), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1207), .B(n_1221), .Y(n_1206) );
INVx3_ASAP7_75t_L g1301 ( .A(n_1207), .Y(n_1301) );
A2O1A1Ixp33_ASAP7_75t_L g1319 ( .A1(n_1207), .A2(n_1320), .B(n_1321), .C(n_1322), .Y(n_1319) );
NAND2xp5_ASAP7_75t_L g1382 ( .A(n_1207), .B(n_1279), .Y(n_1382) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1215), .Y(n_1207) );
AND2x6_ASAP7_75t_L g1209 ( .A(n_1210), .B(n_1211), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1210), .B(n_1214), .Y(n_1213) );
AND2x4_ASAP7_75t_L g1216 ( .A(n_1210), .B(n_1217), .Y(n_1216) );
AND2x6_ASAP7_75t_L g1219 ( .A(n_1210), .B(n_1220), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1210), .B(n_1214), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1210), .B(n_1214), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1217 ( .A(n_1212), .B(n_1218), .Y(n_1217) );
INVx2_ASAP7_75t_L g1418 ( .A(n_1219), .Y(n_1418) );
HB1xp67_ASAP7_75t_L g1485 ( .A(n_1220), .Y(n_1485) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1221), .Y(n_1292) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1221), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1221), .B(n_1261), .Y(n_1321) );
NAND2xp5_ASAP7_75t_L g1327 ( .A(n_1221), .B(n_1328), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1361 ( .A(n_1221), .B(n_1243), .Y(n_1361) );
NAND3xp33_ASAP7_75t_L g1367 ( .A(n_1221), .B(n_1337), .C(n_1368), .Y(n_1367) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1222), .B(n_1279), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_1222), .B(n_1294), .Y(n_1293) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1222), .Y(n_1298) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1222), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1222), .B(n_1243), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1223), .B(n_1225), .Y(n_1222) );
OAI211xp5_ASAP7_75t_SL g1226 ( .A1(n_1227), .A2(n_1237), .B(n_1251), .C(n_1268), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1229), .B(n_1233), .Y(n_1228) );
NOR2xp33_ASAP7_75t_L g1362 ( .A(n_1229), .B(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1230), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1230), .B(n_1256), .Y(n_1265) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1230), .Y(n_1274) );
OR2x2_ASAP7_75t_L g1295 ( .A(n_1230), .B(n_1255), .Y(n_1295) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_1230), .B(n_1234), .Y(n_1299) );
NAND2xp5_ASAP7_75t_L g1306 ( .A(n_1230), .B(n_1233), .Y(n_1306) );
NAND2x1_ASAP7_75t_L g1230 ( .A(n_1231), .B(n_1232), .Y(n_1230) );
OR2x2_ASAP7_75t_L g1263 ( .A(n_1233), .B(n_1264), .Y(n_1263) );
OR2x2_ASAP7_75t_L g1272 ( .A(n_1233), .B(n_1273), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_1233), .B(n_1276), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1233), .B(n_1265), .Y(n_1325) );
OR2x2_ASAP7_75t_L g1333 ( .A(n_1233), .B(n_1295), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1352 ( .A(n_1233), .B(n_1313), .Y(n_1352) );
NAND2xp5_ASAP7_75t_L g1374 ( .A(n_1233), .B(n_1254), .Y(n_1374) );
INVx2_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1234), .B(n_1248), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1234), .B(n_1267), .Y(n_1266) );
AOI22xp5_ASAP7_75t_L g1268 ( .A1(n_1234), .A2(n_1269), .B1(n_1271), .B2(n_1275), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1318 ( .A(n_1234), .B(n_1259), .Y(n_1318) );
NOR2xp33_ASAP7_75t_L g1335 ( .A(n_1234), .B(n_1336), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1234), .B(n_1255), .Y(n_1347) );
OR2x2_ASAP7_75t_L g1381 ( .A(n_1234), .B(n_1295), .Y(n_1381) );
OR2x2_ASAP7_75t_L g1386 ( .A(n_1234), .B(n_1256), .Y(n_1386) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1234), .B(n_1256), .Y(n_1406) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1236), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1247), .Y(n_1237) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1238), .Y(n_1328) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1238), .Y(n_1402) );
NAND2xp5_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1243), .Y(n_1238) );
INVx2_ASAP7_75t_L g1261 ( .A(n_1239), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1239), .B(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
OR2x2_ASAP7_75t_L g1270 ( .A(n_1240), .B(n_1243), .Y(n_1270) );
INVx2_ASAP7_75t_SL g1278 ( .A(n_1240), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1240), .B(n_1276), .Y(n_1294) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_1240), .B(n_1279), .Y(n_1343) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_1240), .B(n_1282), .Y(n_1370) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1241), .B(n_1242), .Y(n_1240) );
CKINVDCx5p33_ASAP7_75t_R g1279 ( .A(n_1243), .Y(n_1279) );
AOI221xp5_ASAP7_75t_L g1281 ( .A1(n_1243), .A2(n_1254), .B1(n_1282), .B2(n_1285), .C(n_1289), .Y(n_1281) );
AOI221xp5_ASAP7_75t_L g1302 ( .A1(n_1243), .A2(n_1256), .B1(n_1303), .B2(n_1307), .C(n_1310), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1392 ( .A(n_1243), .B(n_1248), .Y(n_1392) );
NAND2xp5_ASAP7_75t_L g1409 ( .A(n_1243), .B(n_1410), .Y(n_1409) );
AND2x4_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1246), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1247), .B(n_1254), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1247), .B(n_1305), .Y(n_1304) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1247), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1247), .B(n_1347), .Y(n_1346) );
OAI211xp5_ASAP7_75t_L g1355 ( .A1(n_1247), .A2(n_1356), .B(n_1358), .C(n_1360), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1388 ( .A(n_1247), .B(n_1389), .Y(n_1388) );
OR2x2_ASAP7_75t_L g1408 ( .A(n_1247), .B(n_1306), .Y(n_1408) );
CKINVDCx5p33_ASAP7_75t_R g1247 ( .A(n_1248), .Y(n_1247) );
INVx3_ASAP7_75t_L g1276 ( .A(n_1248), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1248), .B(n_1292), .Y(n_1291) );
NAND2xp5_ASAP7_75t_L g1412 ( .A(n_1248), .B(n_1287), .Y(n_1412) );
AND2x4_ASAP7_75t_SL g1248 ( .A(n_1249), .B(n_1250), .Y(n_1248) );
OAI22xp33_ASAP7_75t_L g1251 ( .A1(n_1252), .A2(n_1261), .B1(n_1262), .B2(n_1266), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1253), .B(n_1261), .Y(n_1252) );
NAND2xp5_ASAP7_75t_L g1253 ( .A(n_1254), .B(n_1260), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1323 ( .A(n_1254), .B(n_1324), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1255), .B(n_1259), .Y(n_1254) );
OAI322xp33_ASAP7_75t_L g1289 ( .A1(n_1255), .A2(n_1261), .A3(n_1290), .B1(n_1293), .B2(n_1295), .C1(n_1296), .C2(n_1299), .Y(n_1289) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
OR2x2_ASAP7_75t_L g1273 ( .A(n_1256), .B(n_1274), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1258), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1260), .B(n_1313), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1376 ( .A(n_1260), .B(n_1265), .Y(n_1376) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1261), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1358 ( .A(n_1261), .B(n_1359), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_1261), .B(n_1376), .Y(n_1375) );
NAND2xp5_ASAP7_75t_L g1398 ( .A(n_1261), .B(n_1271), .Y(n_1398) );
AND2x2_ASAP7_75t_L g1415 ( .A(n_1261), .B(n_1292), .Y(n_1415) );
O2A1O1Ixp33_ASAP7_75t_L g1399 ( .A1(n_1262), .A2(n_1400), .B(n_1402), .C(n_1403), .Y(n_1399) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
OR2x2_ASAP7_75t_L g1283 ( .A(n_1264), .B(n_1284), .Y(n_1283) );
OAI22xp5_ASAP7_75t_SL g1391 ( .A1(n_1264), .A2(n_1296), .B1(n_1392), .B2(n_1393), .Y(n_1391) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1296 ( .A(n_1269), .B(n_1297), .Y(n_1296) );
AOI322xp5_ASAP7_75t_L g1317 ( .A1(n_1269), .A2(n_1291), .A3(n_1318), .B1(n_1319), .B2(n_1323), .C1(n_1325), .C2(n_1326), .Y(n_1317) );
INVx2_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1414 ( .A(n_1271), .B(n_1276), .Y(n_1414) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1273), .Y(n_1313) );
NOR2xp33_ASAP7_75t_L g1357 ( .A(n_1273), .B(n_1342), .Y(n_1357) );
NOR2xp33_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1277), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1276), .B(n_1309), .Y(n_1308) );
CKINVDCx14_ASAP7_75t_R g1340 ( .A(n_1276), .Y(n_1340) );
NOR2xp33_ASAP7_75t_L g1364 ( .A(n_1276), .B(n_1287), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_1276), .B(n_1278), .Y(n_1368) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1277), .Y(n_1309) );
OR2x2_ASAP7_75t_L g1277 ( .A(n_1278), .B(n_1279), .Y(n_1277) );
INVx2_ASAP7_75t_L g1287 ( .A(n_1278), .Y(n_1287) );
A2O1A1Ixp33_ASAP7_75t_L g1372 ( .A1(n_1278), .A2(n_1373), .B(n_1375), .C(n_1377), .Y(n_1372) );
A2O1A1Ixp33_ASAP7_75t_L g1404 ( .A1(n_1278), .A2(n_1345), .B(n_1405), .C(n_1407), .Y(n_1404) );
NAND2xp5_ASAP7_75t_L g1330 ( .A(n_1279), .B(n_1301), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1279), .B(n_1339), .Y(n_1338) );
OAI221xp5_ASAP7_75t_SL g1280 ( .A1(n_1281), .A2(n_1300), .B1(n_1302), .B2(n_1314), .C(n_1317), .Y(n_1280) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1284), .Y(n_1324) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1287), .B(n_1288), .Y(n_1286) );
NOR2xp33_ASAP7_75t_L g1394 ( .A(n_1287), .B(n_1395), .Y(n_1394) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1288), .Y(n_1322) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1294), .Y(n_1350) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1295), .Y(n_1337) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
CKINVDCx14_ASAP7_75t_R g1354 ( .A(n_1300), .Y(n_1354) );
OAI221xp5_ASAP7_75t_L g1378 ( .A1(n_1300), .A2(n_1379), .B1(n_1382), .B2(n_1383), .C(n_1384), .Y(n_1378) );
OAI31xp33_ASAP7_75t_SL g1390 ( .A1(n_1300), .A2(n_1391), .A3(n_1394), .B(n_1397), .Y(n_1390) );
CKINVDCx14_ASAP7_75t_R g1300 ( .A(n_1301), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1301), .B(n_1316), .Y(n_1315) );
AOI322xp5_ASAP7_75t_L g1334 ( .A1(n_1303), .A2(n_1335), .A3(n_1338), .B1(n_1340), .B2(n_1341), .C1(n_1344), .C2(n_1346), .Y(n_1334) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1309), .B(n_1312), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1383 ( .A(n_1309), .B(n_1380), .Y(n_1383) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
NOR2xp33_ASAP7_75t_L g1336 ( .A(n_1313), .B(n_1337), .Y(n_1336) );
CKINVDCx14_ASAP7_75t_R g1314 ( .A(n_1315), .Y(n_1314) );
OR2x2_ASAP7_75t_L g1342 ( .A(n_1316), .B(n_1343), .Y(n_1342) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1318), .Y(n_1411) );
OAI211xp5_ASAP7_75t_SL g1397 ( .A1(n_1322), .A2(n_1398), .B(n_1399), .C(n_1413), .Y(n_1397) );
NAND2xp5_ASAP7_75t_L g1401 ( .A(n_1324), .B(n_1337), .Y(n_1401) );
NOR2xp33_ASAP7_75t_L g1393 ( .A(n_1325), .B(n_1365), .Y(n_1393) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_1325), .B(n_1332), .Y(n_1396) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
OAI211xp5_ASAP7_75t_SL g1329 ( .A1(n_1330), .A2(n_1331), .B(n_1334), .C(n_1348), .Y(n_1329) );
INVxp67_ASAP7_75t_SL g1377 ( .A(n_1330), .Y(n_1377) );
INVxp67_ASAP7_75t_L g1359 ( .A(n_1331), .Y(n_1359) );
OR2x2_ASAP7_75t_L g1331 ( .A(n_1332), .B(n_1333), .Y(n_1331) );
INVx2_ASAP7_75t_L g1365 ( .A(n_1333), .Y(n_1365) );
AOI221xp5_ASAP7_75t_SL g1360 ( .A1(n_1338), .A2(n_1361), .B1(n_1362), .B2(n_1365), .C(n_1366), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1348 ( .A(n_1339), .B(n_1349), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1379 ( .A(n_1340), .B(n_1380), .Y(n_1379) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1343), .Y(n_1389) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1345), .Y(n_1371) );
NOR2xp33_ASAP7_75t_L g1349 ( .A(n_1350), .B(n_1351), .Y(n_1349) );
INVx2_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
AOI211xp5_ASAP7_75t_L g1353 ( .A1(n_1354), .A2(n_1355), .B(n_1369), .C(n_1378), .Y(n_1353) );
INVxp67_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
OAI21xp5_ASAP7_75t_L g1384 ( .A1(n_1365), .A2(n_1385), .B(n_1387), .Y(n_1384) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
OAI21xp5_ASAP7_75t_L g1369 ( .A1(n_1370), .A2(n_1371), .B(n_1372), .Y(n_1369) );
OAI21xp33_ASAP7_75t_L g1413 ( .A1(n_1373), .A2(n_1414), .B(n_1415), .Y(n_1413) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
NAND2xp5_ASAP7_75t_SL g1403 ( .A(n_1404), .B(n_1409), .Y(n_1403) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
NOR2xp33_ASAP7_75t_L g1410 ( .A(n_1411), .B(n_1412), .Y(n_1410) );
CKINVDCx20_ASAP7_75t_R g1416 ( .A(n_1417), .Y(n_1416) );
CKINVDCx20_ASAP7_75t_R g1417 ( .A(n_1418), .Y(n_1417) );
HB1xp67_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
HB1xp67_ASAP7_75t_L g1481 ( .A(n_1421), .Y(n_1481) );
NOR3xp33_ASAP7_75t_L g1428 ( .A(n_1429), .B(n_1440), .C(n_1441), .Y(n_1428) );
NOR3xp33_ASAP7_75t_L g1429 ( .A(n_1430), .B(n_1433), .C(n_1439), .Y(n_1429) );
NOR2xp33_ASAP7_75t_L g1430 ( .A(n_1431), .B(n_1432), .Y(n_1430) );
NOR2xp33_ASAP7_75t_L g1461 ( .A(n_1431), .B(n_1457), .Y(n_1461) );
NAND2xp5_ASAP7_75t_L g1433 ( .A(n_1434), .B(n_1437), .Y(n_1433) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1443), .Y(n_1442) );
INVx2_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
NAND3xp33_ASAP7_75t_L g1449 ( .A(n_1450), .B(n_1454), .C(n_1468), .Y(n_1449) );
AOI22xp5_ASAP7_75t_L g1454 ( .A1(n_1455), .A2(n_1460), .B1(n_1466), .B2(n_1467), .Y(n_1454) );
AOI22xp5_ASAP7_75t_L g1460 ( .A1(n_1456), .A2(n_1461), .B1(n_1462), .B2(n_1463), .Y(n_1460) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
BUFx3_ASAP7_75t_L g1471 ( .A(n_1472), .Y(n_1471) );
BUFx2_ASAP7_75t_SL g1475 ( .A(n_1476), .Y(n_1475) );
BUFx3_ASAP7_75t_L g1476 ( .A(n_1477), .Y(n_1476) );
INVxp33_ASAP7_75t_SL g1478 ( .A(n_1479), .Y(n_1478) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1481), .Y(n_1480) );
HB1xp67_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
OAI21xp5_ASAP7_75t_L g1484 ( .A1(n_1485), .A2(n_1486), .B(n_1487), .Y(n_1484) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
endmodule