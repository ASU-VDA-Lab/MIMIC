module fake_jpeg_11435_n_645 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_645);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_645;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_SL g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_63),
.Y(n_175)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_66),
.Y(n_149)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_68),
.Y(n_213)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_70),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_42),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_73),
.B(n_77),
.Y(n_133)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_74),
.Y(n_211)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_76),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_39),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_78),
.B(n_81),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_79),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_82),
.B(n_84),
.Y(n_156)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_38),
.B(n_18),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_38),
.B(n_18),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_85),
.B(n_93),
.Y(n_162)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_87),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_88),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_91),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_92),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_39),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx6_ASAP7_75t_SL g95 ( 
.A(n_42),
.Y(n_95)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_95),
.Y(n_203)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_96),
.B(n_97),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_39),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_98),
.Y(n_178)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_100),
.Y(n_168)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_102),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g198 ( 
.A(n_103),
.Y(n_198)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_19),
.Y(n_104)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_31),
.Y(n_106)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_107),
.Y(n_191)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_32),
.Y(n_108)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_108),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_60),
.B(n_17),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_109),
.B(n_110),
.Y(n_183)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_22),
.Y(n_110)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_112),
.Y(n_202)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_32),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_113),
.Y(n_216)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_32),
.Y(n_115)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_115),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_17),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_117),
.B(n_119),
.Y(n_204)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_29),
.Y(n_118)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_24),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_46),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_120),
.B(n_121),
.Y(n_206)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_24),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_32),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_122),
.B(n_124),
.Y(n_217)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_49),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g154 ( 
.A(n_123),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_46),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_19),
.Y(n_125)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_46),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_54),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g127 ( 
.A(n_42),
.Y(n_127)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_52),
.Y(n_129)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_127),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_136),
.B(n_158),
.Y(n_222)
);

BUFx12_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_148),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_33),
.C(n_58),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_157),
.B(n_159),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_83),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_107),
.B(n_44),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_161),
.B(n_32),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_108),
.B(n_33),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_166),
.B(n_162),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_113),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_170),
.B(n_174),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_115),
.Y(n_174)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_61),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_179),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_92),
.B(n_103),
.Y(n_184)
);

NAND2x1_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_208),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_79),
.B(n_59),
.C(n_58),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_185),
.B(n_66),
.Y(n_240)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_64),
.Y(n_186)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_186),
.Y(n_218)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_75),
.Y(n_187)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_89),
.Y(n_188)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_188),
.Y(n_252)
);

BUFx16f_ASAP7_75t_L g193 ( 
.A(n_88),
.Y(n_193)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_91),
.Y(n_195)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_195),
.Y(n_258)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_98),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_111),
.Y(n_197)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_112),
.Y(n_199)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_199),
.Y(n_236)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_66),
.A2(n_37),
.B(n_23),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_201),
.B(n_54),
.Y(n_266)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_116),
.Y(n_207)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

NAND2x1_ASAP7_75t_L g208 ( 
.A(n_123),
.B(n_47),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_86),
.Y(n_209)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_68),
.Y(n_210)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_210),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_71),
.Y(n_212)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_76),
.Y(n_214)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_214),
.Y(n_264)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_87),
.Y(n_215)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

O2A1O1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_217),
.A2(n_47),
.B(n_50),
.C(n_35),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_219),
.B(n_240),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_175),
.B(n_40),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_220),
.B(n_225),
.Y(n_317)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_150),
.Y(n_221)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_221),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_150),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_223),
.B(n_229),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_167),
.A2(n_80),
.B1(n_41),
.B2(n_34),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_228),
.A2(n_247),
.B1(n_279),
.B2(n_281),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_176),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_133),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_233),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_183),
.B(n_37),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_234),
.B(n_237),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_183),
.B(n_25),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_133),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g295 ( 
.A(n_241),
.B(n_259),
.C(n_265),
.Y(n_295)
);

AND2x2_ASAP7_75t_SL g244 ( 
.A(n_130),
.B(n_105),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_244),
.B(n_230),
.C(n_248),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_156),
.B(n_88),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_246),
.B(n_260),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_167),
.A2(n_41),
.B1(n_34),
.B2(n_54),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_184),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_248),
.Y(n_339)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_165),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_249),
.Y(n_318)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_211),
.Y(n_250)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_250),
.Y(n_304)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_176),
.Y(n_251)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_251),
.Y(n_306)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_193),
.Y(n_253)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_253),
.Y(n_331)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_206),
.Y(n_254)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_254),
.Y(n_316)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_141),
.Y(n_257)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_257),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_204),
.B(n_44),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_156),
.B(n_105),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_162),
.B(n_27),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_261),
.B(n_266),
.Y(n_302)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_206),
.Y(n_262)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_262),
.Y(n_321)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_180),
.Y(n_263)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_204),
.B(n_25),
.Y(n_265)
);

CKINVDCx11_ASAP7_75t_R g267 ( 
.A(n_203),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_267),
.B(n_269),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_134),
.Y(n_268)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_268),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_216),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_200),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_270),
.Y(n_294)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_182),
.Y(n_272)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_272),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_273),
.B(n_276),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_134),
.Y(n_274)
);

INVx6_ASAP7_75t_L g320 ( 
.A(n_274),
.Y(n_320)
);

OA22x2_ASAP7_75t_L g275 ( 
.A1(n_208),
.A2(n_114),
.B1(n_55),
.B2(n_41),
.Y(n_275)
);

AOI22x1_ASAP7_75t_L g346 ( 
.A1(n_275),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_166),
.B(n_23),
.Y(n_276)
);

INVx6_ASAP7_75t_SL g277 ( 
.A(n_217),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_277),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_132),
.B(n_142),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_286),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_154),
.A2(n_34),
.B1(n_52),
.B2(n_55),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_163),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_154),
.A2(n_55),
.B1(n_59),
.B2(n_57),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_137),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_282),
.Y(n_315)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_143),
.Y(n_283)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_283),
.Y(n_328)
);

INVx11_ASAP7_75t_L g284 ( 
.A(n_140),
.Y(n_284)
);

BUFx8_ASAP7_75t_L g327 ( 
.A(n_284),
.Y(n_327)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_171),
.Y(n_285)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_285),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_216),
.B(n_57),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_160),
.Y(n_287)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_287),
.Y(n_345)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_169),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_288),
.Y(n_343)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_191),
.Y(n_289)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_289),
.Y(n_329)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_163),
.Y(n_290)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_290),
.Y(n_337)
);

OAI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_138),
.A2(n_50),
.B1(n_27),
.B2(n_45),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_291),
.A2(n_293),
.B1(n_168),
.B2(n_164),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_135),
.B(n_45),
.Y(n_292)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_292),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_155),
.A2(n_36),
.B1(n_35),
.B2(n_17),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_238),
.B(n_36),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_299),
.B(n_305),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_301),
.B(n_307),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_233),
.B(n_205),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_220),
.A2(n_189),
.B1(n_192),
.B2(n_146),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_308),
.A2(n_314),
.B1(n_332),
.B2(n_231),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_219),
.A2(n_138),
.B1(n_146),
.B2(n_189),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_313),
.A2(n_322),
.B1(n_268),
.B2(n_224),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_278),
.A2(n_192),
.B1(n_173),
.B2(n_178),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_244),
.B(n_168),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_319),
.B(n_338),
.C(n_270),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_275),
.A2(n_178),
.B1(n_164),
.B2(n_202),
.Y(n_322)
);

BUFx24_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

INVx13_ASAP7_75t_L g388 ( 
.A(n_323),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_244),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_324),
.B(n_340),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_230),
.B(n_151),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_325),
.B(n_330),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_242),
.B(n_172),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_279),
.A2(n_173),
.B1(n_202),
.B2(n_131),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_257),
.A2(n_139),
.B1(n_153),
.B2(n_145),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_335),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_243),
.B(n_177),
.C(n_152),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_222),
.Y(n_340)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_236),
.Y(n_344)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_344),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_346),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_218),
.B(n_227),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_347),
.B(n_350),
.Y(n_372)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_239),
.Y(n_349)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_349),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_226),
.B(n_147),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_235),
.B(n_144),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_290),
.Y(n_373)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_318),
.Y(n_355)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_355),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_325),
.B(n_275),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_357),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_302),
.B(n_245),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_358),
.B(n_316),
.Y(n_409)
);

INVx6_ASAP7_75t_SL g361 ( 
.A(n_323),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_361),
.Y(n_408)
);

INVx6_ASAP7_75t_L g363 ( 
.A(n_298),
.Y(n_363)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_363),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_351),
.A2(n_131),
.B1(n_291),
.B2(n_231),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_364),
.A2(n_367),
.B1(n_383),
.B2(n_362),
.Y(n_410)
);

AND2x6_ASAP7_75t_L g369 ( 
.A(n_323),
.B(n_228),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_369),
.B(n_374),
.Y(n_423)
);

AND2x2_ASAP7_75t_SL g370 ( 
.A(n_301),
.B(n_288),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_371),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_249),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_373),
.B(n_377),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_347),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_342),
.B(n_282),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_375),
.B(n_378),
.Y(n_412)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_350),
.Y(n_376)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_376),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_305),
.B(n_252),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_333),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_303),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_379),
.B(n_381),
.Y(n_403)
);

INVx3_ASAP7_75t_SL g380 ( 
.A(n_298),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g407 ( 
.A1(n_380),
.A2(n_397),
.B1(n_399),
.B2(n_315),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_353),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_326),
.B(n_252),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_382),
.B(n_393),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_351),
.A2(n_258),
.B1(n_280),
.B2(n_274),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_332),
.A2(n_255),
.B1(n_258),
.B2(n_264),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_384),
.Y(n_405)
);

BUFx24_ASAP7_75t_SL g385 ( 
.A(n_297),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_385),
.B(n_390),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_308),
.A2(n_255),
.B1(n_264),
.B2(n_256),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_386),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_319),
.Y(n_400)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_330),
.Y(n_389)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_389),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_300),
.B(n_232),
.Y(n_390)
);

INVx13_ASAP7_75t_L g391 ( 
.A(n_331),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_391),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_312),
.A2(n_281),
.B(n_247),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_392),
.A2(n_359),
.B(n_357),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_341),
.B(n_232),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_317),
.B(n_190),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_394),
.A2(n_371),
.B(n_377),
.Y(n_430)
);

AND2x6_ASAP7_75t_L g395 ( 
.A(n_295),
.B(n_284),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_395),
.B(n_398),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_396),
.A2(n_320),
.B1(n_294),
.B2(n_329),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_336),
.A2(n_314),
.B1(n_346),
.B2(n_318),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_306),
.B(n_253),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_SL g399 ( 
.A1(n_352),
.A2(n_256),
.B1(n_149),
.B2(n_224),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_400),
.B(n_402),
.C(n_417),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_370),
.B(n_299),
.C(n_338),
.Y(n_402)
);

AO22x1_ASAP7_75t_L g404 ( 
.A1(n_376),
.A2(n_313),
.B1(n_322),
.B2(n_307),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_404),
.B(n_409),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_407),
.A2(n_431),
.B(n_405),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_410),
.A2(n_414),
.B1(n_429),
.B2(n_434),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_367),
.A2(n_321),
.B1(n_310),
.B2(n_339),
.Y(n_414)
);

AO22x1_ASAP7_75t_SL g415 ( 
.A1(n_389),
.A2(n_337),
.B1(n_328),
.B2(n_309),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_415),
.B(n_418),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_370),
.B(n_387),
.C(n_354),
.Y(n_417)
);

OAI32xp33_ASAP7_75t_L g418 ( 
.A1(n_368),
.A2(n_348),
.A3(n_304),
.B1(n_352),
.B2(n_315),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_419),
.A2(n_420),
.B1(n_424),
.B2(n_426),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_354),
.A2(n_294),
.B1(n_320),
.B2(n_296),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_370),
.B(n_311),
.C(n_309),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_421),
.B(n_373),
.C(n_365),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_371),
.A2(n_343),
.B1(n_331),
.B2(n_296),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_422),
.A2(n_435),
.B(n_392),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_354),
.A2(n_311),
.B1(n_328),
.B2(n_334),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_396),
.A2(n_334),
.B1(n_345),
.B2(n_343),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_361),
.A2(n_327),
.B(n_345),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_428),
.A2(n_388),
.B(n_398),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_362),
.A2(n_327),
.B1(n_15),
.B2(n_210),
.Y(n_429)
);

AND2x2_ASAP7_75t_SL g471 ( 
.A(n_430),
.B(n_365),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_360),
.A2(n_327),
.B1(n_15),
.B2(n_46),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_368),
.A2(n_198),
.B(n_181),
.Y(n_435)
);

INVx11_ASAP7_75t_L g441 ( 
.A(n_408),
.Y(n_441)
);

BUFx2_ASAP7_75t_SL g498 ( 
.A(n_441),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_403),
.B(n_374),
.Y(n_442)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_442),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_412),
.Y(n_443)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_443),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_444),
.B(n_471),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_403),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_445),
.B(n_451),
.Y(n_475)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_415),
.Y(n_446)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_446),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_427),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_447),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_423),
.A2(n_437),
.B1(n_438),
.B2(n_432),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_448),
.A2(n_406),
.B1(n_435),
.B2(n_421),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_437),
.A2(n_357),
.B1(n_381),
.B2(n_372),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_452),
.A2(n_453),
.B(n_467),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_431),
.A2(n_369),
.B(n_388),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_454),
.B(n_474),
.C(n_450),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_401),
.B(n_372),
.Y(n_455)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_455),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_416),
.B(n_356),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_456),
.B(n_466),
.Y(n_479)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_415),
.Y(n_457)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_457),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_401),
.B(n_356),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_458),
.B(n_460),
.Y(n_484)
);

CKINVDCx14_ASAP7_75t_R g459 ( 
.A(n_416),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_459),
.B(n_430),
.Y(n_476)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_432),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_425),
.B(n_379),
.Y(n_461)
);

NAND3xp33_ASAP7_75t_L g493 ( 
.A(n_461),
.B(n_468),
.C(n_469),
.Y(n_493)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_438),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_462),
.B(n_463),
.Y(n_488)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_427),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_424),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_465),
.Y(n_504)
);

AOI322xp5_ASAP7_75t_L g466 ( 
.A1(n_414),
.A2(n_395),
.A3(n_358),
.B1(n_388),
.B2(n_383),
.C1(n_382),
.C2(n_375),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_409),
.B(n_390),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_418),
.B(n_366),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_420),
.B(n_366),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_470),
.B(n_472),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_433),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_413),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_473),
.B(n_363),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_417),
.B(n_394),
.C(n_355),
.Y(n_474)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_476),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_445),
.B(n_436),
.Y(n_480)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_480),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_481),
.B(n_492),
.C(n_502),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_456),
.B(n_436),
.Y(n_482)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_482),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_453),
.A2(n_411),
.B(n_405),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_483),
.A2(n_486),
.B(n_494),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_485),
.A2(n_444),
.B1(n_470),
.B2(n_449),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_464),
.A2(n_406),
.B(n_428),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_450),
.B(n_400),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_487),
.B(n_452),
.Y(n_526)
);

AOI22x1_ASAP7_75t_L g489 ( 
.A1(n_440),
.A2(n_411),
.B1(n_404),
.B2(n_406),
.Y(n_489)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_489),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_461),
.B(n_402),
.Y(n_491)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_491),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_394),
.C(n_422),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_448),
.A2(n_404),
.B1(n_413),
.B2(n_433),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_499),
.B(n_472),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_454),
.B(n_419),
.C(n_426),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_442),
.B(n_363),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_503),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_451),
.B(n_380),
.C(n_391),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_505),
.B(n_487),
.C(n_502),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_468),
.B(n_391),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_467),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_446),
.A2(n_380),
.B1(n_198),
.B2(n_181),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_508),
.A2(n_467),
.B(n_441),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_494),
.A2(n_464),
.B1(n_469),
.B2(n_440),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_512),
.A2(n_514),
.B1(n_516),
.B2(n_531),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_480),
.A2(n_457),
.B1(n_449),
.B2(n_455),
.Y(n_514)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_498),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_515),
.Y(n_540)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_517),
.Y(n_544)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_519),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_496),
.A2(n_439),
.B1(n_471),
.B2(n_458),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_520),
.A2(n_521),
.B1(n_523),
.B2(n_504),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_496),
.A2(n_439),
.B1(n_471),
.B2(n_462),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_522),
.B(n_484),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_500),
.A2(n_471),
.B1(n_460),
.B2(n_466),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_524),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_490),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_525),
.B(n_530),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_526),
.B(n_488),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_481),
.B(n_473),
.C(n_463),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_528),
.B(n_535),
.C(n_538),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_SL g529 ( 
.A(n_479),
.B(n_148),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_SL g560 ( 
.A(n_529),
.B(n_488),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_486),
.A2(n_0),
.B(n_2),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_475),
.A2(n_500),
.B1(n_477),
.B2(n_497),
.Y(n_531)
);

HAxp5_ASAP7_75t_SL g532 ( 
.A(n_507),
.B(n_495),
.CON(n_532),
.SN(n_532)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_532),
.A2(n_507),
.B(n_495),
.Y(n_539)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_477),
.Y(n_533)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_533),
.Y(n_547)
);

NOR3xp33_ASAP7_75t_SL g534 ( 
.A(n_493),
.B(n_0),
.C(n_3),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_534),
.B(n_478),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_492),
.B(n_0),
.C(n_3),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_485),
.B(n_0),
.C(n_4),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_539),
.B(n_557),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_528),
.B(n_478),
.Y(n_542)
);

NAND3xp33_ASAP7_75t_L g576 ( 
.A(n_542),
.B(n_552),
.C(n_530),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_522),
.B(n_505),
.C(n_507),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_543),
.B(n_554),
.C(n_556),
.Y(n_567)
);

A2O1A1Ixp33_ASAP7_75t_SL g549 ( 
.A1(n_527),
.A2(n_483),
.B(n_489),
.C(n_475),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_549),
.B(n_510),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_550),
.B(n_563),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_511),
.B(n_536),
.Y(n_551)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_551),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_537),
.B(n_497),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_509),
.B(n_503),
.C(n_489),
.Y(n_554)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_555),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_509),
.B(n_484),
.C(n_490),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_523),
.B(n_508),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_558),
.B(n_563),
.Y(n_583)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_517),
.Y(n_559)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_559),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_560),
.B(n_562),
.Y(n_579)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_533),
.Y(n_561)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_561),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_526),
.B(n_504),
.C(n_501),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_SL g564 ( 
.A(n_557),
.B(n_518),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_564),
.B(n_568),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_553),
.A2(n_520),
.B1(n_521),
.B2(n_527),
.Y(n_566)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_566),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_556),
.B(n_514),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_540),
.Y(n_572)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_572),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_546),
.B(n_515),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_573),
.B(n_576),
.Y(n_598)
);

OAI21x1_ASAP7_75t_SL g589 ( 
.A1(n_575),
.A2(n_584),
.B(n_547),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_554),
.B(n_512),
.Y(n_577)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_577),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_544),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_578),
.B(n_580),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_548),
.A2(n_513),
.B1(n_538),
.B2(n_534),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_543),
.B(n_510),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_581),
.B(n_562),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_583),
.B(n_545),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_541),
.B(n_501),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g608 ( 
.A(n_586),
.B(n_579),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_587),
.B(n_9),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_583),
.B(n_541),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_588),
.B(n_593),
.Y(n_604)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_589),
.Y(n_606)
);

NOR2xp67_ASAP7_75t_L g590 ( 
.A(n_571),
.B(n_531),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_590),
.A2(n_591),
.B(n_596),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_575),
.A2(n_558),
.B(n_524),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_567),
.B(n_549),
.C(n_529),
.Y(n_593)
);

OAI321xp33_ASAP7_75t_L g595 ( 
.A1(n_582),
.A2(n_549),
.A3(n_499),
.B1(n_532),
.B2(n_560),
.C(n_535),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_595),
.A2(n_574),
.B1(n_566),
.B2(n_569),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_567),
.B(n_549),
.C(n_5),
.Y(n_596)
);

A2O1A1Ixp33_ASAP7_75t_L g597 ( 
.A1(n_575),
.A2(n_4),
.B(n_7),
.C(n_8),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_597),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_SL g599 ( 
.A1(n_570),
.A2(n_8),
.B(n_9),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_599),
.B(n_596),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_570),
.A2(n_578),
.B(n_565),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_SL g611 ( 
.A1(n_600),
.A2(n_572),
.B(n_10),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_588),
.B(n_581),
.C(n_571),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_605),
.B(n_610),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_607),
.B(n_611),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_608),
.B(n_592),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_586),
.B(n_587),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_609),
.B(n_608),
.C(n_604),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_585),
.B(n_579),
.C(n_574),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_SL g612 ( 
.A1(n_598),
.A2(n_9),
.B(n_10),
.Y(n_612)
);

AOI21x1_ASAP7_75t_SL g619 ( 
.A1(n_612),
.A2(n_594),
.B(n_599),
.Y(n_619)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_613),
.Y(n_618)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_615),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_600),
.B(n_11),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_616),
.B(n_597),
.Y(n_621)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_619),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_620),
.B(n_626),
.Y(n_632)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_621),
.Y(n_630)
);

NOR2xp67_ASAP7_75t_L g624 ( 
.A(n_605),
.B(n_602),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_624),
.B(n_613),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_610),
.B(n_601),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_625),
.B(n_627),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_609),
.B(n_591),
.C(n_593),
.Y(n_627)
);

BUFx12_ASAP7_75t_L g629 ( 
.A(n_619),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_629),
.B(n_618),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_623),
.A2(n_606),
.B1(n_614),
.B2(n_603),
.Y(n_631)
);

AO21x1_ASAP7_75t_L g636 ( 
.A1(n_631),
.A2(n_617),
.B(n_623),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_634),
.A2(n_627),
.B(n_616),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_635),
.B(n_637),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_SL g639 ( 
.A1(n_636),
.A2(n_638),
.B1(n_633),
.B2(n_630),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_632),
.B(n_622),
.Y(n_637)
);

XOR2xp5_ASAP7_75t_L g641 ( 
.A(n_639),
.B(n_628),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_641),
.B(n_640),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_642),
.B(n_629),
.C(n_12),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_643),
.B(n_12),
.C(n_13),
.Y(n_644)
);

XOR2xp5_ASAP7_75t_L g645 ( 
.A(n_644),
.B(n_13),
.Y(n_645)
);


endmodule