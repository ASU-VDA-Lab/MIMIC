module fake_jpeg_103_n_603 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_603);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_603;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_18),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_6),
.Y(n_55)
);

INVx11_ASAP7_75t_SL g56 ( 
.A(n_4),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_13),
.B(n_9),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_58),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_18),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_59),
.B(n_73),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g195 ( 
.A(n_61),
.Y(n_195)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_63),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_65),
.Y(n_157)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_68),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_69),
.Y(n_174)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_72),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_10),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_74),
.Y(n_151)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_76),
.Y(n_197)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_23),
.B(n_10),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_78),
.B(n_88),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_79),
.Y(n_201)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_80),
.Y(n_196)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_81),
.Y(n_169)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_86),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_20),
.B(n_10),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_89),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_23),
.B(n_18),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_47),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_91),
.Y(n_181)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_92),
.Y(n_168)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_23),
.B(n_10),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_95),
.B(n_101),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_96),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_97),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_98),
.Y(n_220)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_20),
.B(n_9),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_102),
.Y(n_219)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_103),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_43),
.B(n_17),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_104),
.B(n_124),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_106),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_107),
.Y(n_214)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_108),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_110),
.Y(n_173)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_30),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_111),
.Y(n_210)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_41),
.Y(n_114)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_114),
.Y(n_178)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_28),
.Y(n_115)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_19),
.Y(n_116)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_19),
.Y(n_117)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_39),
.Y(n_118)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_118),
.Y(n_200)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_31),
.Y(n_119)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_28),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_120),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_31),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_48),
.B1(n_54),
.B2(n_43),
.Y(n_146)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_30),
.Y(n_122)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_122),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_39),
.Y(n_123)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_123),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_40),
.B(n_11),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_32),
.Y(n_125)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_125),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_32),
.Y(n_126)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_28),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_41),
.Y(n_149)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_28),
.Y(n_128)
);

BUFx2_ASAP7_75t_R g166 ( 
.A(n_128),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_78),
.A2(n_52),
.B1(n_55),
.B2(n_38),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_138),
.A2(n_153),
.B1(n_162),
.B2(n_177),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_124),
.A2(n_60),
.B1(n_69),
.B2(n_68),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_141),
.A2(n_146),
.B1(n_155),
.B2(n_179),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_64),
.B(n_41),
.C(n_55),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_142),
.B(n_17),
.Y(n_242)
);

OR2x4_ASAP7_75t_L g147 ( 
.A(n_61),
.B(n_48),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_147),
.B(n_194),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_149),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_105),
.A2(n_52),
.B1(n_24),
.B2(n_38),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_76),
.A2(n_54),
.B1(n_24),
.B2(n_36),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_79),
.A2(n_53),
.B1(n_44),
.B2(n_32),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_106),
.A2(n_107),
.B1(n_86),
.B2(n_102),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_71),
.A2(n_36),
.B1(n_45),
.B2(n_35),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_80),
.B(n_45),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_180),
.B(n_186),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_125),
.A2(n_53),
.B1(n_44),
.B2(n_33),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_182),
.A2(n_218),
.B1(n_0),
.B2(n_1),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_83),
.B(n_42),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_116),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_188),
.B(n_198),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_120),
.A2(n_98),
.B1(n_109),
.B2(n_33),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_190),
.A2(n_207),
.B1(n_1),
.B2(n_2),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_117),
.B(n_42),
.Y(n_194)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_118),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_123),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_199),
.B(n_202),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_65),
.B(n_35),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_126),
.B(n_53),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_215),
.Y(n_226)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_72),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_205),
.B(n_213),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_120),
.A2(n_44),
.B1(n_33),
.B2(n_28),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_94),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_92),
.B(n_29),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_99),
.B(n_29),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_1),
.Y(n_234)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_128),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_217),
.B(n_195),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_100),
.A2(n_29),
.B1(n_1),
.B2(n_2),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_221),
.Y(n_310)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_223),
.Y(n_325)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_224),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_225),
.A2(n_273),
.B1(n_222),
.B2(n_275),
.Y(n_311)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_227),
.Y(n_340)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_228),
.Y(n_343)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_229),
.Y(n_315)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_230),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_155),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_231),
.A2(n_248),
.B1(n_252),
.B2(n_254),
.Y(n_308)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_232),
.Y(n_313)
);

OA22x2_ASAP7_75t_L g300 ( 
.A1(n_233),
.A2(n_231),
.B1(n_261),
.B2(n_274),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_234),
.B(n_247),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_149),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_235),
.Y(n_322)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_161),
.Y(n_236)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_236),
.Y(n_321)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_197),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_237),
.Y(n_312)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_140),
.Y(n_238)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_238),
.Y(n_352)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_239),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_139),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_240),
.B(n_241),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_139),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_242),
.B(n_262),
.C(n_250),
.Y(n_317)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_170),
.Y(n_243)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_243),
.Y(n_351)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_176),
.Y(n_244)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_244),
.Y(n_355)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_245),
.Y(n_347)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_246),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_164),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_129),
.A2(n_12),
.B1(n_13),
.B2(n_17),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_133),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_249),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_154),
.A2(n_12),
.B1(n_3),
.B2(n_4),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_250),
.B(n_268),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_173),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_251),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_178),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_211),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_253),
.B(n_259),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_212),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_130),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_255),
.B(n_261),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_175),
.B(n_5),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_256),
.B(n_265),
.Y(n_320)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_197),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_257),
.Y(n_341)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_201),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_258),
.Y(n_342)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

BUFx2_ASAP7_75t_SL g260 ( 
.A(n_166),
.Y(n_260)
);

INVx13_ASAP7_75t_L g318 ( 
.A(n_260),
.Y(n_318)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_182),
.Y(n_261)
);

AND2x2_ASAP7_75t_SL g262 ( 
.A(n_143),
.B(n_5),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_206),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_263),
.B(n_278),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_165),
.B(n_5),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_144),
.B(n_5),
.Y(n_267)
);

AND2x2_ASAP7_75t_SL g309 ( 
.A(n_267),
.B(n_269),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_150),
.A2(n_136),
.B1(n_131),
.B2(n_160),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_172),
.B(n_169),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_130),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_271),
.B(n_274),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_207),
.A2(n_190),
.B(n_185),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_272),
.A2(n_291),
.B(n_264),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_201),
.A2(n_209),
.B1(n_133),
.B2(n_163),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_273),
.A2(n_275),
.B1(n_249),
.B2(n_237),
.Y(n_304)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_218),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_209),
.A2(n_174),
.B1(n_163),
.B2(n_214),
.Y(n_275)
);

INVx11_ASAP7_75t_L g276 ( 
.A(n_185),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_276),
.A2(n_224),
.B1(n_230),
.B2(n_229),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_145),
.B(n_151),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_277),
.B(n_286),
.Y(n_326)
);

AOI32xp33_ASAP7_75t_L g278 ( 
.A1(n_204),
.A2(n_208),
.A3(n_158),
.B1(n_192),
.B2(n_156),
.Y(n_278)
);

INVx8_ASAP7_75t_L g280 ( 
.A(n_152),
.Y(n_280)
);

NOR2x1_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_297),
.Y(n_305)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_135),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_281),
.B(n_284),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_162),
.A2(n_181),
.B1(n_137),
.B2(n_148),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_282),
.A2(n_295),
.B1(n_276),
.B2(n_223),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_156),
.A2(n_192),
.B1(n_167),
.B2(n_210),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_283),
.A2(n_285),
.B1(n_290),
.B2(n_292),
.Y(n_302)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_196),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_210),
.A2(n_173),
.B1(n_184),
.B2(n_204),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_174),
.B(n_157),
.Y(n_286)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_157),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_288),
.B(n_258),
.Y(n_354)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_196),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_289),
.B(n_294),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_132),
.A2(n_159),
.B1(n_168),
.B2(n_134),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_159),
.B(n_132),
.Y(n_291)
);

AND2x2_ASAP7_75t_SL g335 ( 
.A(n_291),
.B(n_294),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_168),
.A2(n_134),
.B1(n_183),
.B2(n_152),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_183),
.B(n_134),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_219),
.A2(n_155),
.B1(n_146),
.B2(n_104),
.Y(n_295)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_219),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_298),
.B(n_291),
.Y(n_338)
);

A2O1A1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_226),
.A2(n_256),
.B(n_234),
.C(n_296),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_299),
.B(n_247),
.Y(n_366)
);

OAI21xp33_ASAP7_75t_SL g367 ( 
.A1(n_300),
.A2(n_330),
.B(n_247),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_301),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_304),
.A2(n_345),
.B1(n_341),
.B2(n_342),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_266),
.A2(n_226),
.B1(n_272),
.B2(n_222),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_306),
.A2(n_311),
.B1(n_314),
.B2(n_339),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_286),
.A2(n_296),
.B1(n_279),
.B2(n_277),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_317),
.B(n_309),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_242),
.B(n_265),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_323),
.B(n_334),
.C(n_289),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_262),
.A2(n_268),
.B1(n_267),
.B2(n_287),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_327),
.A2(n_280),
.B1(n_334),
.B2(n_299),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_269),
.B(n_262),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_335),
.B(n_336),
.Y(n_383)
);

NAND3xp33_ASAP7_75t_SL g337 ( 
.A(n_293),
.B(n_269),
.C(n_227),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_337),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_338),
.B(n_251),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_221),
.A2(n_228),
.B1(n_245),
.B2(n_239),
.Y(n_339)
);

AOI22x1_ASAP7_75t_L g345 ( 
.A1(n_267),
.A2(n_297),
.B1(n_238),
.B2(n_288),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_270),
.A2(n_236),
.B1(n_243),
.B2(n_244),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_346),
.A2(n_344),
.B1(n_353),
.B2(n_351),
.Y(n_392)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_354),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_356),
.B(n_377),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_357),
.B(n_366),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_329),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_358),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_314),
.B(n_281),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_360),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_232),
.C(n_284),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_362),
.B(n_376),
.C(n_388),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_326),
.B(n_246),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_364),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_326),
.B(n_253),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_320),
.B(n_259),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_365),
.B(n_368),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_367),
.A2(n_390),
.B(n_350),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_320),
.B(n_257),
.Y(n_368)
);

OAI21xp33_ASAP7_75t_SL g417 ( 
.A1(n_369),
.A2(n_315),
.B(n_316),
.Y(n_417)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_340),
.Y(n_371)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_371),
.Y(n_404)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_340),
.Y(n_372)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_372),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_327),
.B(n_263),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_373),
.B(n_389),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_374),
.Y(n_429)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_310),
.Y(n_375)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_375),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_309),
.B(n_335),
.C(n_317),
.Y(n_376)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_310),
.Y(n_378)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_378),
.Y(n_415)
);

OAI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_330),
.A2(n_311),
.B1(n_324),
.B2(n_332),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_379),
.A2(n_392),
.B1(n_399),
.B2(n_319),
.Y(n_402)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_352),
.Y(n_380)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_380),
.Y(n_416)
);

AOI32xp33_ASAP7_75t_L g381 ( 
.A1(n_348),
.A2(n_322),
.A3(n_324),
.B1(n_309),
.B2(n_335),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_381),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_349),
.A2(n_333),
.B1(n_348),
.B2(n_304),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_382),
.A2(n_384),
.B1(n_385),
.B2(n_394),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_308),
.A2(n_300),
.B1(n_303),
.B2(n_322),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_300),
.A2(n_303),
.B1(n_345),
.B2(n_338),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_303),
.B(n_354),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_391),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_328),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_387),
.B(n_397),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_346),
.B(n_343),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_325),
.B(n_343),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_305),
.A2(n_345),
.B(n_302),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_325),
.B(n_344),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_305),
.B(n_307),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_313),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_300),
.A2(n_341),
.B1(n_342),
.B2(n_347),
.Y(n_394)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_351),
.Y(n_396)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_396),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_315),
.B(n_316),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_355),
.Y(n_398)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_398),
.Y(n_431)
);

OAI22xp33_ASAP7_75t_SL g399 ( 
.A1(n_302),
.A2(n_352),
.B1(n_313),
.B2(n_347),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_391),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_400),
.B(n_359),
.Y(n_452)
);

NOR2x1_ASAP7_75t_L g401 ( 
.A(n_383),
.B(n_355),
.Y(n_401)
);

A2O1A1Ixp33_ASAP7_75t_L g465 ( 
.A1(n_401),
.A2(n_408),
.B(n_409),
.C(n_403),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_402),
.A2(n_412),
.B(n_420),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_411),
.B(n_419),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_SL g412 ( 
.A(n_383),
.B(n_331),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_417),
.A2(n_426),
.B1(n_418),
.B2(n_431),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_370),
.B(n_321),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_377),
.B(n_321),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_362),
.C(n_386),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_363),
.B(n_312),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_423),
.B(n_424),
.Y(n_445)
);

CKINVDCx14_ASAP7_75t_R g424 ( 
.A(n_393),
.Y(n_424)
);

OAI32xp33_ASAP7_75t_L g426 ( 
.A1(n_383),
.A2(n_350),
.A3(n_312),
.B1(n_329),
.B2(n_318),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_426),
.B(n_427),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_364),
.B(n_312),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_356),
.B(n_318),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_430),
.B(n_434),
.C(n_378),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_384),
.A2(n_385),
.B1(n_374),
.B2(n_394),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_433),
.A2(n_425),
.B1(n_424),
.B2(n_402),
.Y(n_446)
);

XNOR2x1_ASAP7_75t_L g434 ( 
.A(n_376),
.B(n_331),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_416),
.Y(n_436)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_436),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_429),
.A2(n_382),
.B1(n_370),
.B2(n_390),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_437),
.A2(n_467),
.B1(n_468),
.B2(n_405),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_401),
.Y(n_439)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_439),
.Y(n_498)
);

CKINVDCx14_ASAP7_75t_R g440 ( 
.A(n_408),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_440),
.B(n_452),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_400),
.A2(n_361),
.B1(n_368),
.B2(n_365),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_441),
.A2(n_446),
.B1(n_448),
.B2(n_449),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_410),
.Y(n_442)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_442),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_443),
.B(n_460),
.C(n_462),
.Y(n_470)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_413),
.Y(n_444)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_444),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_425),
.A2(n_373),
.B1(n_387),
.B2(n_392),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_433),
.A2(n_388),
.B1(n_359),
.B2(n_372),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_450),
.B(n_430),
.Y(n_477)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_413),
.Y(n_451)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_451),
.Y(n_495)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_415),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_453),
.B(n_454),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_410),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_409),
.A2(n_395),
.B1(n_371),
.B2(n_375),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_455),
.A2(n_404),
.B1(n_414),
.B2(n_416),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_380),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_457),
.B(n_458),
.Y(n_491)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_415),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_423),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_459),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_421),
.B(n_396),
.C(n_398),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_427),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_461),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_421),
.B(n_358),
.C(n_395),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_420),
.A2(n_358),
.B(n_432),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_463),
.A2(n_464),
.B(n_465),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_412),
.A2(n_401),
.B(n_405),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_418),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_466),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_406),
.A2(n_403),
.B1(n_419),
.B2(n_411),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_450),
.B(n_434),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_471),
.B(n_478),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_473),
.A2(n_482),
.B1(n_487),
.B2(n_497),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_443),
.B(n_434),
.C(n_435),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_476),
.B(n_477),
.C(n_493),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_443),
.B(n_435),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_446),
.A2(n_417),
.B1(n_406),
.B2(n_422),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_460),
.B(n_422),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_484),
.B(n_486),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_460),
.B(n_431),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_441),
.A2(n_404),
.B1(n_414),
.B2(n_407),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_488),
.A2(n_489),
.B1(n_457),
.B2(n_438),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_448),
.A2(n_449),
.B1(n_456),
.B2(n_468),
.Y(n_489)
);

XNOR2x1_ASAP7_75t_L g490 ( 
.A(n_465),
.B(n_437),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_490),
.B(n_496),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_436),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_492),
.B(n_481),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_462),
.B(n_454),
.C(n_442),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_462),
.B(n_464),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_456),
.A2(n_440),
.B1(n_461),
.B2(n_459),
.Y(n_497)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_483),
.Y(n_502)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_502),
.Y(n_525)
);

CKINVDCx14_ASAP7_75t_R g503 ( 
.A(n_480),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_503),
.Y(n_528)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_483),
.Y(n_504)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_504),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_478),
.B(n_465),
.C(n_463),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_505),
.B(n_496),
.C(n_477),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_469),
.A2(n_447),
.B(n_445),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_507),
.B(n_511),
.Y(n_537)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_508),
.Y(n_532)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_491),
.Y(n_510)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_510),
.Y(n_541)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_491),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_494),
.Y(n_512)
);

INVxp33_ASAP7_75t_SL g536 ( 
.A(n_512),
.Y(n_536)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_480),
.Y(n_513)
);

INVx11_ASAP7_75t_L g531 ( 
.A(n_513),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_473),
.A2(n_445),
.B1(n_452),
.B2(n_455),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_514),
.A2(n_517),
.B1(n_479),
.B2(n_489),
.Y(n_535)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_494),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_515),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_488),
.B(n_467),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_516),
.B(n_519),
.Y(n_542)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_495),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_518),
.A2(n_522),
.B1(n_523),
.B2(n_479),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_493),
.B(n_438),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_486),
.B(n_447),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_520),
.B(n_484),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_472),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_521),
.A2(n_475),
.B1(n_474),
.B2(n_495),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_485),
.A2(n_444),
.B1(n_451),
.B2(n_453),
.Y(n_522)
);

INVx6_ASAP7_75t_L g523 ( 
.A(n_472),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_527),
.B(n_505),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_529),
.A2(n_506),
.B1(n_514),
.B2(n_502),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_501),
.B(n_470),
.C(n_476),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_530),
.B(n_539),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_SL g533 ( 
.A(n_520),
.B(n_471),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_500),
.B(n_470),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_534),
.B(n_499),
.Y(n_550)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_535),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_501),
.B(n_469),
.C(n_498),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_540),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g543 ( 
.A(n_532),
.B(n_511),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_543),
.B(n_551),
.Y(n_561)
);

CKINVDCx14_ASAP7_75t_R g544 ( 
.A(n_537),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_544),
.A2(n_552),
.B1(n_556),
.B2(n_541),
.Y(n_562)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_538),
.Y(n_546)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_546),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_530),
.B(n_499),
.C(n_500),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_548),
.B(n_549),
.Y(n_559)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_532),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_550),
.B(n_554),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_534),
.B(n_539),
.C(n_527),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_535),
.A2(n_497),
.B1(n_518),
.B2(n_516),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_537),
.A2(n_507),
.B(n_504),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_555),
.A2(n_541),
.B1(n_524),
.B2(n_525),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_529),
.A2(n_506),
.B1(n_510),
.B2(n_522),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_557),
.B(n_526),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_558),
.B(n_565),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_547),
.B(n_542),
.C(n_533),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_560),
.B(n_564),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_562),
.B(n_490),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_554),
.A2(n_528),
.B(n_540),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_563),
.A2(n_553),
.B(n_536),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_551),
.B(n_542),
.C(n_509),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_548),
.B(n_509),
.C(n_524),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_567),
.B(n_538),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_553),
.B(n_521),
.Y(n_568)
);

NOR2xp67_ASAP7_75t_L g573 ( 
.A(n_568),
.B(n_552),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_550),
.B(n_482),
.C(n_487),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_569),
.B(n_556),
.C(n_555),
.Y(n_575)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_571),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_573),
.B(n_574),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_559),
.B(n_545),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_575),
.B(n_579),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_570),
.B(n_557),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_576),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_561),
.B(n_523),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_577),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_580),
.B(n_581),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_566),
.B(n_475),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_576),
.B(n_565),
.C(n_558),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_586),
.B(n_575),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_SL g587 ( 
.A1(n_572),
.A2(n_580),
.B(n_578),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_SL g590 ( 
.A1(n_587),
.A2(n_564),
.B(n_560),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_590),
.B(n_589),
.C(n_585),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_591),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_586),
.B(n_570),
.Y(n_592)
);

NOR3xp33_ASAP7_75t_L g595 ( 
.A(n_592),
.B(n_593),
.C(n_594),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_588),
.B(n_579),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_584),
.B(n_567),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_597),
.A2(n_589),
.B(n_582),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_598),
.A2(n_599),
.B(n_595),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_596),
.B(n_585),
.C(n_583),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_600),
.B(n_517),
.C(n_515),
.Y(n_601)
);

MAJx2_ASAP7_75t_L g602 ( 
.A(n_601),
.B(n_512),
.C(n_531),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_602),
.B(n_531),
.Y(n_603)
);


endmodule