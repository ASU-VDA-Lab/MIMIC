module fake_jpeg_1303_n_691 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_691);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_691;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_540;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_398;
wire n_583;
wire n_56;
wire n_240;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_553;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_61),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_62),
.B(n_76),
.Y(n_141)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_64),
.Y(n_162)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_65),
.Y(n_172)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g209 ( 
.A(n_66),
.Y(n_209)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_67),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_70),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_71),
.Y(n_160)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_72),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_19),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_73),
.B(n_100),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_75),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_26),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_77),
.Y(n_174)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_78),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g229 ( 
.A(n_79),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_83),
.Y(n_175)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_84),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_85),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_86),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_87),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_88),
.Y(n_187)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_89),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_90),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_91),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_93),
.Y(n_166)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_94),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_55),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_95),
.B(n_116),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_98),
.Y(n_183)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_99),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_20),
.B(n_18),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_101),
.Y(n_180)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_102),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_104),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_46),
.B(n_17),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_105),
.B(n_108),
.Y(n_164)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_106),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_20),
.B(n_17),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

CKINVDCx9p33_ASAP7_75t_R g210 ( 
.A(n_109),
.Y(n_210)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_33),
.Y(n_114)
);

INVx11_ASAP7_75t_L g161 ( 
.A(n_114),
.Y(n_161)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_55),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_22),
.Y(n_118)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_118),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_21),
.B(n_0),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_119),
.B(n_48),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_121),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_22),
.Y(n_122)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_33),
.Y(n_123)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_123),
.Y(n_221)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_124),
.Y(n_217)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_33),
.Y(n_125)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_49),
.Y(n_126)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_126),
.Y(n_224)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_53),
.Y(n_127)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_127),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_24),
.Y(n_128)
);

INVx11_ASAP7_75t_L g212 ( 
.A(n_128),
.Y(n_212)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_129),
.Y(n_230)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_24),
.Y(n_130)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_53),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_52),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_54),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_132),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_90),
.A2(n_58),
.B1(n_54),
.B2(n_35),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_142),
.A2(n_152),
.B1(n_184),
.B2(n_0),
.Y(n_277)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_81),
.Y(n_150)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_150),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_91),
.A2(n_97),
.B1(n_120),
.B2(n_113),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_72),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_155),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_165),
.Y(n_242)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_67),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_171),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_79),
.B(n_21),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_178),
.B(n_198),
.Y(n_250)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_79),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_181),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_89),
.A2(n_58),
.B1(n_54),
.B2(n_40),
.Y(n_184)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_70),
.Y(n_186)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_80),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_188),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_86),
.B(n_35),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_190),
.Y(n_285)
);

CKINVDCx12_ASAP7_75t_R g192 ( 
.A(n_74),
.Y(n_192)
);

CKINVDCx12_ASAP7_75t_R g290 ( 
.A(n_192),
.Y(n_290)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_101),
.Y(n_195)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_195),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_93),
.Y(n_196)
);

INVx11_ASAP7_75t_L g307 ( 
.A(n_196),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_81),
.B(n_40),
.Y(n_198)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_82),
.A2(n_39),
.B(n_48),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_201),
.B(n_202),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_82),
.B(n_39),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_114),
.Y(n_204)
);

NAND2xp33_ASAP7_75t_SL g314 ( 
.A(n_204),
.B(n_9),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_99),
.B(n_41),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_205),
.B(n_218),
.Y(n_291)
);

INVx6_ASAP7_75t_SL g206 ( 
.A(n_123),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_206),
.Y(n_301)
);

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_96),
.Y(n_208)
);

INVx5_ASAP7_75t_L g293 ( 
.A(n_208),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_117),
.B(n_41),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_32),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_128),
.B(n_34),
.Y(n_218)
);

INVx11_ASAP7_75t_L g219 ( 
.A(n_128),
.Y(n_219)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_45),
.Y(n_249)
);

INVx11_ASAP7_75t_L g222 ( 
.A(n_118),
.Y(n_222)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_122),
.B(n_28),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_223),
.B(n_226),
.Y(n_302)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_59),
.Y(n_225)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_68),
.B(n_34),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_69),
.B(n_32),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_231),
.B(n_182),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_232),
.B(n_237),
.Y(n_363)
);

AND2x2_ASAP7_75t_SL g233 ( 
.A(n_214),
.B(n_52),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_233),
.Y(n_376)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_136),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_234),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_141),
.B(n_28),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_162),
.B(n_30),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_238),
.B(n_243),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g239 ( 
.A1(n_190),
.A2(n_45),
.B(n_43),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_239),
.B(n_289),
.Y(n_325)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_172),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_241),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_164),
.B(n_30),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_L g244 ( 
.A1(n_142),
.A2(n_132),
.B1(n_111),
.B2(n_103),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_244),
.A2(n_277),
.B1(n_158),
.B2(n_154),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_249),
.B(n_294),
.Y(n_320)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_150),
.Y(n_251)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_251),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_252),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_215),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_253),
.Y(n_351)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_174),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_254),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_255),
.Y(n_364)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_219),
.Y(n_256)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_256),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_258),
.Y(n_347)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_133),
.Y(n_259)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_259),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_152),
.A2(n_88),
.B1(n_85),
.B2(n_83),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_260),
.A2(n_266),
.B1(n_295),
.B2(n_311),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_176),
.B(n_43),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_261),
.B(n_271),
.Y(n_322)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_166),
.Y(n_262)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_262),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_133),
.Y(n_263)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_263),
.Y(n_365)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_212),
.Y(n_264)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_264),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_210),
.A2(n_24),
.B1(n_52),
.B2(n_58),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_265),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_144),
.A2(n_52),
.B1(n_75),
.B2(n_2),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_185),
.Y(n_267)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_267),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_148),
.Y(n_269)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_269),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_183),
.B(n_52),
.Y(n_271)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_148),
.Y(n_272)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_272),
.Y(n_339)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_222),
.Y(n_273)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_273),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_189),
.B(n_193),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_274),
.B(n_282),
.Y(n_338)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_191),
.Y(n_275)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_275),
.Y(n_350)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_151),
.Y(n_276)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_276),
.Y(n_355)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_154),
.Y(n_278)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_278),
.Y(n_358)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_228),
.Y(n_279)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_279),
.Y(n_361)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_230),
.Y(n_280)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_280),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_134),
.B(n_1),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_281),
.Y(n_368)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_197),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_147),
.B(n_2),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_283),
.B(n_286),
.Y(n_356)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_168),
.Y(n_284)
);

INVx11_ASAP7_75t_L g337 ( 
.A(n_284),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_229),
.B(n_3),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_229),
.B(n_170),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_287),
.B(n_292),
.Y(n_359)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_157),
.Y(n_289)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_217),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_170),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_144),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_207),
.B(n_5),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_296),
.B(n_297),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_146),
.B(n_5),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_224),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_298),
.B(n_300),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_199),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_299),
.B(n_306),
.Y(n_367)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_135),
.Y(n_300)
);

INVx5_ASAP7_75t_SL g303 ( 
.A(n_199),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_303),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_180),
.B(n_7),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_304),
.B(n_305),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_139),
.B(n_7),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_194),
.B(n_8),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_153),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_308),
.B(n_310),
.Y(n_369)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_177),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_309),
.B(n_312),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_204),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_175),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_311)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_221),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_313),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_314),
.A2(n_200),
.B(n_145),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_194),
.B(n_10),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_315),
.A2(n_290),
.B1(n_303),
.B2(n_301),
.Y(n_331)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_209),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_317),
.Y(n_345)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_159),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_321),
.Y(n_396)
);

AO22x1_ASAP7_75t_L g323 ( 
.A1(n_285),
.A2(n_213),
.B1(n_203),
.B2(n_161),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_323),
.B(n_336),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_331),
.B(n_378),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_242),
.B(n_140),
.C(n_160),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_333),
.B(n_335),
.C(n_370),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_334),
.A2(n_342),
.B1(n_352),
.B2(n_353),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_281),
.B(n_200),
.Y(n_335)
);

OA22x2_ASAP7_75t_L g336 ( 
.A1(n_260),
.A2(n_167),
.B1(n_173),
.B2(n_163),
.Y(n_336)
);

O2A1O1Ixp33_ASAP7_75t_L g341 ( 
.A1(n_268),
.A2(n_167),
.B(n_149),
.C(n_145),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_341),
.B(n_371),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_233),
.A2(n_211),
.B1(n_163),
.B2(n_137),
.Y(n_342)
);

AOI32xp33_ASAP7_75t_L g346 ( 
.A1(n_302),
.A2(n_209),
.A3(n_211),
.B1(n_196),
.B2(n_137),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_346),
.B(n_143),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_244),
.A2(n_187),
.B1(n_175),
.B2(n_179),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g425 ( 
.A1(n_349),
.A2(n_372),
.B1(n_353),
.B2(n_366),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_233),
.A2(n_156),
.B1(n_187),
.B2(n_179),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_311),
.A2(n_156),
.B1(n_158),
.B2(n_173),
.Y(n_353)
);

MAJx2_ASAP7_75t_L g370 ( 
.A(n_291),
.B(n_250),
.C(n_249),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_314),
.B(n_239),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_245),
.A2(n_149),
.B1(n_138),
.B2(n_169),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_235),
.B(n_208),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_265),
.A2(n_138),
.B1(n_208),
.B2(n_182),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_379),
.A2(n_380),
.B1(n_366),
.B2(n_352),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_266),
.A2(n_182),
.B1(n_169),
.B2(n_168),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_345),
.Y(n_381)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_381),
.Y(n_433)
);

OR2x2_ASAP7_75t_SL g382 ( 
.A(n_376),
.B(n_235),
.Y(n_382)
);

NOR2x1_ASAP7_75t_L g472 ( 
.A(n_382),
.B(n_143),
.Y(n_472)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_345),
.Y(n_383)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_383),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_325),
.A2(n_245),
.B1(n_313),
.B2(n_262),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_384),
.A2(n_411),
.B(n_423),
.Y(n_461)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_350),
.Y(n_385)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_385),
.Y(n_443)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_350),
.Y(n_386)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_386),
.Y(n_448)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_326),
.Y(n_388)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_388),
.Y(n_450)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_357),
.Y(n_389)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_389),
.Y(n_449)
);

INVx13_ASAP7_75t_L g390 ( 
.A(n_354),
.Y(n_390)
);

BUFx5_ASAP7_75t_L g435 ( 
.A(n_390),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_334),
.A2(n_272),
.B1(n_259),
.B2(n_278),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_391),
.A2(n_414),
.B1(n_330),
.B2(n_339),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_335),
.B(n_248),
.C(n_246),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_392),
.B(n_421),
.C(n_355),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_395),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_360),
.B(n_317),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_397),
.B(n_406),
.Y(n_459)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_326),
.Y(n_398)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_398),
.Y(n_456)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_361),
.Y(n_399)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_399),
.Y(n_464)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_361),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_400),
.B(n_403),
.Y(n_462)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_377),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g404 ( 
.A1(n_343),
.A2(n_275),
.B1(n_257),
.B2(n_288),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_404),
.A2(n_409),
.B1(n_425),
.B2(n_429),
.Y(n_454)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_377),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_405),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_363),
.B(n_270),
.Y(n_406)
);

INVx13_ASAP7_75t_L g407 ( 
.A(n_354),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g468 ( 
.A1(n_407),
.A2(n_410),
.B1(n_412),
.B2(n_415),
.Y(n_468)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_319),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_408),
.B(n_420),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_362),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_321),
.B(n_273),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_357),
.Y(n_412)
);

INVx3_ASAP7_75t_SL g413 ( 
.A(n_362),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_413),
.B(n_419),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_371),
.A2(n_252),
.B1(n_258),
.B2(n_255),
.Y(n_414)
);

INVx13_ASAP7_75t_L g415 ( 
.A(n_337),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_322),
.B(n_270),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_416),
.B(n_418),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_417),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_338),
.B(n_288),
.Y(n_418)
);

INVx5_ASAP7_75t_L g419 ( 
.A(n_351),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_339),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_333),
.B(n_276),
.C(n_289),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_327),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_422),
.B(n_430),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_378),
.A2(n_295),
.B(n_293),
.Y(n_423)
);

CKINVDCx14_ASAP7_75t_R g424 ( 
.A(n_325),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_424),
.Y(n_432)
);

INVx13_ASAP7_75t_L g426 ( 
.A(n_337),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_426),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_359),
.B(n_143),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_427),
.B(n_355),
.Y(n_469)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_325),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_428),
.A2(n_323),
.B1(n_369),
.B2(n_373),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_342),
.A2(n_307),
.B1(n_247),
.B2(n_256),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_344),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_393),
.A2(n_375),
.B1(n_320),
.B2(n_373),
.Y(n_436)
);

AO21x2_ASAP7_75t_L g513 ( 
.A1(n_436),
.A2(n_467),
.B(n_403),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_396),
.A2(n_341),
.B(n_367),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_438),
.A2(n_441),
.B(n_472),
.Y(n_502)
);

AO22x1_ASAP7_75t_L g444 ( 
.A1(n_402),
.A2(n_373),
.B1(n_323),
.B2(n_336),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_444),
.B(n_451),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_446),
.A2(n_453),
.B1(n_386),
.B2(n_399),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_387),
.B(n_370),
.Y(n_447)
);

XNOR2x1_ASAP7_75t_L g479 ( 
.A(n_447),
.B(n_457),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_381),
.B(n_356),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_383),
.B(n_368),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_452),
.B(n_455),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_396),
.A2(n_374),
.B1(n_336),
.B2(n_358),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_392),
.B(n_411),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_411),
.B(n_368),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_458),
.B(n_401),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_387),
.B(n_332),
.C(n_318),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_460),
.B(n_408),
.C(n_422),
.Y(n_480)
);

XOR2x2_ASAP7_75t_L g463 ( 
.A(n_394),
.B(n_382),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_463),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_423),
.A2(n_374),
.B(n_236),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_465),
.A2(n_251),
.B(n_236),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_421),
.B(n_331),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_466),
.B(n_411),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_393),
.A2(n_336),
.B1(n_358),
.B2(n_330),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_469),
.B(n_473),
.Y(n_488)
);

OAI21xp33_ASAP7_75t_L g482 ( 
.A1(n_472),
.A2(n_401),
.B(n_402),
.Y(n_482)
);

NAND3xp33_ASAP7_75t_L g473 ( 
.A(n_397),
.B(n_348),
.C(n_324),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_462),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_474),
.B(n_484),
.Y(n_538)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_462),
.Y(n_476)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_476),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_480),
.B(n_483),
.C(n_491),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_SL g521 ( 
.A(n_481),
.B(n_432),
.Y(n_521)
);

NOR3xp33_ASAP7_75t_L g537 ( 
.A(n_482),
.B(n_502),
.C(n_507),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_447),
.B(n_457),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_462),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_434),
.Y(n_485)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_485),
.Y(n_525)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_486),
.Y(n_549)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_449),
.Y(n_487)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_487),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_439),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_489),
.B(n_497),
.Y(n_547)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_449),
.Y(n_490)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_490),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_460),
.B(n_384),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_461),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_492),
.B(n_512),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_466),
.B(n_388),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_493),
.B(n_498),
.C(n_511),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_441),
.B(n_438),
.Y(n_494)
);

OAI22xp33_ASAP7_75t_SL g539 ( 
.A1(n_494),
.A2(n_470),
.B1(n_450),
.B2(n_445),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_461),
.A2(n_402),
.B(n_409),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_495),
.A2(n_413),
.B(n_431),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_433),
.A2(n_442),
.B1(n_455),
.B2(n_453),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_496),
.A2(n_442),
.B1(n_444),
.B2(n_467),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_469),
.B(n_385),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_463),
.B(n_398),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_499),
.B(n_505),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_440),
.B(n_348),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_500),
.B(n_501),
.Y(n_514)
);

INVx8_ASAP7_75t_L g501 ( 
.A(n_440),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_451),
.B(n_348),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_503),
.B(n_509),
.Y(n_516)
);

OAI22x1_ASAP7_75t_L g504 ( 
.A1(n_458),
.A2(n_414),
.B1(n_390),
.B2(n_407),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_504),
.A2(n_506),
.B(n_471),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_444),
.A2(n_391),
.B1(n_419),
.B2(n_420),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_434),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_443),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_508),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_436),
.B(n_410),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_443),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_510),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_452),
.B(n_400),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_433),
.B(n_405),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_513),
.A2(n_465),
.B1(n_446),
.B2(n_432),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_515),
.A2(n_533),
.B1(n_540),
.B2(n_505),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_501),
.B(n_459),
.Y(n_517)
);

CKINVDCx16_ASAP7_75t_R g575 ( 
.A(n_517),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_480),
.B(n_439),
.Y(n_518)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_518),
.Y(n_562)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_519),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_SL g566 ( 
.A(n_521),
.B(n_481),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_487),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_522),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_488),
.B(n_478),
.Y(n_523)
);

NOR3xp33_ASAP7_75t_L g583 ( 
.A(n_523),
.B(n_528),
.C(n_535),
.Y(n_583)
);

OAI32xp33_ASAP7_75t_L g524 ( 
.A1(n_475),
.A2(n_437),
.A3(n_448),
.B1(n_464),
.B2(n_456),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_524),
.B(n_527),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_512),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_478),
.B(n_437),
.Y(n_528)
);

OA22x2_ASAP7_75t_L g529 ( 
.A1(n_513),
.A2(n_468),
.B1(n_454),
.B2(n_448),
.Y(n_529)
);

OA21x2_ASAP7_75t_L g556 ( 
.A1(n_529),
.A2(n_544),
.B(n_504),
.Y(n_556)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_475),
.Y(n_531)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_531),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_496),
.A2(n_470),
.B1(n_445),
.B2(n_464),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_477),
.B(n_456),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_539),
.A2(n_435),
.B1(n_426),
.B2(n_415),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_476),
.B(n_450),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_541),
.B(n_545),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_511),
.B(n_431),
.Y(n_543)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_543),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_486),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_513),
.A2(n_430),
.B1(n_417),
.B2(n_413),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_546),
.A2(n_508),
.B1(n_510),
.B2(n_507),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_479),
.B(n_340),
.C(n_389),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_551),
.B(n_493),
.C(n_483),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_555),
.B(n_558),
.C(n_576),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_556),
.A2(n_561),
.B1(n_569),
.B2(n_571),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_548),
.B(n_498),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_557),
.B(n_574),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_542),
.B(n_479),
.C(n_491),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_559),
.A2(n_532),
.B1(n_519),
.B2(n_520),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_541),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_560),
.B(n_563),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_514),
.A2(n_513),
.B1(n_477),
.B2(n_494),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_547),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_566),
.B(n_572),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_SL g607 ( 
.A1(n_567),
.A2(n_582),
.B1(n_550),
.B2(n_534),
.Y(n_607)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_526),
.Y(n_568)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_568),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_531),
.A2(n_513),
.B1(n_495),
.B2(n_485),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_545),
.A2(n_506),
.B1(n_492),
.B2(n_502),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_542),
.B(n_412),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_526),
.Y(n_573)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_573),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_548),
.B(n_340),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_551),
.B(n_490),
.C(n_324),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_536),
.B(n_527),
.Y(n_577)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_577),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_536),
.B(n_430),
.Y(n_578)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_578),
.Y(n_595)
);

BUFx24_ASAP7_75t_SL g579 ( 
.A(n_538),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_SL g598 ( 
.A(n_579),
.B(n_581),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_515),
.A2(n_417),
.B1(n_435),
.B2(n_347),
.Y(n_580)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_580),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_543),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_562),
.A2(n_537),
.B(n_530),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_584),
.A2(n_585),
.B1(n_599),
.B2(n_603),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_574),
.B(n_521),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_587),
.B(n_588),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_572),
.B(n_530),
.C(n_520),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_555),
.B(n_544),
.C(n_525),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_590),
.B(n_596),
.C(n_602),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_576),
.B(n_525),
.C(n_532),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_557),
.B(n_516),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_597),
.B(n_608),
.Y(n_611)
);

CKINVDCx14_ASAP7_75t_R g599 ( 
.A(n_553),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_558),
.B(n_532),
.C(n_533),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_552),
.A2(n_569),
.B1(n_564),
.B2(n_553),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_SL g604 ( 
.A1(n_552),
.A2(n_549),
.B1(n_546),
.B2(n_529),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_604),
.B(n_606),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_565),
.B(n_529),
.C(n_540),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_605),
.B(n_556),
.C(n_529),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_566),
.B(n_524),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_607),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_565),
.B(n_549),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_590),
.B(n_573),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_614),
.B(n_624),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_615),
.B(n_600),
.Y(n_635)
);

CKINVDCx14_ASAP7_75t_R g616 ( 
.A(n_593),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_616),
.B(n_629),
.Y(n_636)
);

OAI322xp33_ASAP7_75t_L g617 ( 
.A1(n_598),
.A2(n_570),
.A3(n_583),
.B1(n_564),
.B2(n_577),
.C1(n_568),
.C2(n_556),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_SL g637 ( 
.A(n_617),
.B(n_623),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_SL g619 ( 
.A(n_602),
.B(n_575),
.C(n_570),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_619),
.B(n_622),
.Y(n_648)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_589),
.Y(n_620)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_620),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_586),
.B(n_567),
.C(n_582),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_621),
.B(n_628),
.C(n_631),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_594),
.A2(n_578),
.B(n_550),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_596),
.B(n_554),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_609),
.B(n_534),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_591),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_SL g647 ( 
.A(n_625),
.B(n_10),
.Y(n_647)
);

AOI321xp33_ASAP7_75t_L g627 ( 
.A1(n_606),
.A2(n_328),
.A3(n_522),
.B1(n_365),
.B2(n_347),
.C(n_307),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_SL g640 ( 
.A1(n_627),
.A2(n_585),
.B(n_622),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_586),
.B(n_522),
.C(n_328),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_595),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_603),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_630),
.B(n_592),
.Y(n_641)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_609),
.B(n_329),
.C(n_365),
.Y(n_631)
);

NOR2xp67_ASAP7_75t_L g632 ( 
.A(n_614),
.B(n_588),
.Y(n_632)
);

NOR3xp33_ASAP7_75t_L g660 ( 
.A(n_632),
.B(n_647),
.C(n_649),
.Y(n_660)
);

XNOR2x1_ASAP7_75t_L g653 ( 
.A(n_635),
.B(n_646),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_613),
.A2(n_605),
.B1(n_601),
.B2(n_604),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_SL g650 ( 
.A1(n_638),
.A2(n_613),
.B1(n_615),
.B2(n_611),
.Y(n_650)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_621),
.B(n_592),
.Y(n_639)
);

XNOR2xp5_ASAP7_75t_L g652 ( 
.A(n_639),
.B(n_642),
.Y(n_652)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_640),
.Y(n_656)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_641),
.Y(n_659)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_610),
.B(n_364),
.Y(n_642)
);

XOR2xp5_ASAP7_75t_L g643 ( 
.A(n_610),
.B(n_364),
.Y(n_643)
);

XNOR2xp5_ASAP7_75t_L g654 ( 
.A(n_643),
.B(n_624),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_612),
.B(n_329),
.C(n_351),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_645),
.B(n_631),
.C(n_247),
.Y(n_655)
);

XOR2x2_ASAP7_75t_SL g646 ( 
.A(n_618),
.B(n_240),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_628),
.B(n_253),
.Y(n_649)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_650),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_SL g651 ( 
.A1(n_648),
.A2(n_626),
.B1(n_612),
.B2(n_627),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_651),
.B(n_654),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_655),
.B(n_633),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_637),
.A2(n_240),
.B(n_264),
.Y(n_657)
);

OAI21x1_ASAP7_75t_L g665 ( 
.A1(n_657),
.A2(n_644),
.B(n_643),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_SL g658 ( 
.A1(n_635),
.A2(n_269),
.B1(n_263),
.B2(n_293),
.Y(n_658)
);

MAJx2_ASAP7_75t_L g673 ( 
.A(n_658),
.B(n_12),
.C(n_13),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_648),
.A2(n_284),
.B1(n_169),
.B2(n_168),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_661),
.B(n_662),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_636),
.A2(n_196),
.B1(n_11),
.B2(n_12),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_L g663 ( 
.A1(n_638),
.A2(n_10),
.B(n_11),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_SL g670 ( 
.A1(n_663),
.A2(n_642),
.B(n_634),
.Y(n_670)
);

NAND3xp33_ASAP7_75t_L g674 ( 
.A(n_665),
.B(n_663),
.C(n_655),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_656),
.A2(n_634),
.B(n_639),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_666),
.A2(n_668),
.B(n_653),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_SL g668 ( 
.A1(n_659),
.A2(n_646),
.B(n_645),
.Y(n_668)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_670),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_SL g675 ( 
.A(n_671),
.B(n_672),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_660),
.B(n_633),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_673),
.B(n_14),
.Y(n_677)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_674),
.Y(n_681)
);

NAND3xp33_ASAP7_75t_L g676 ( 
.A(n_669),
.B(n_653),
.C(n_658),
.Y(n_676)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_676),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_677),
.B(n_679),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_SL g684 ( 
.A1(n_678),
.A2(n_667),
.B(n_652),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_SL g679 ( 
.A(n_664),
.B(n_652),
.Y(n_679)
);

AOI322xp5_ASAP7_75t_L g686 ( 
.A1(n_684),
.A2(n_680),
.A3(n_675),
.B1(n_667),
.B2(n_654),
.C1(n_16),
.C2(n_15),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_682),
.Y(n_685)
);

MAJIxp5_ASAP7_75t_L g687 ( 
.A(n_685),
.B(n_686),
.C(n_681),
.Y(n_687)
);

BUFx24_ASAP7_75t_SL g688 ( 
.A(n_687),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_688),
.B(n_683),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_689),
.A2(n_14),
.B(n_15),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_SL g691 ( 
.A1(n_690),
.A2(n_15),
.B(n_16),
.Y(n_691)
);


endmodule