module fake_jpeg_22780_n_221 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_221);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_221;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_33),
.B(n_34),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_39),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_24),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_1),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_43),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_2),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_31),
.B1(n_24),
.B2(n_22),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_46),
.A2(n_66),
.B1(n_69),
.B2(n_3),
.Y(n_97)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_17),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_51),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_17),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_32),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_16),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_20),
.Y(n_75)
);

CKINVDCx12_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_23),
.B1(n_21),
.B2(n_25),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_57),
.A2(n_26),
.B1(n_15),
.B2(n_16),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_30),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_64),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_65),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_22),
.B1(n_23),
.B2(n_32),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_51),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_23),
.B1(n_29),
.B2(n_19),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_42),
.A2(n_25),
.B1(n_29),
.B2(n_19),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_20),
.B1(n_28),
.B2(n_26),
.Y(n_80)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_75),
.B(n_87),
.Y(n_128)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_62),
.B1(n_71),
.B2(n_52),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_81),
.B(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_30),
.Y(n_82)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_16),
.C(n_30),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_101),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_85),
.A2(n_86),
.B1(n_95),
.B2(n_9),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_26),
.B1(n_15),
.B2(n_16),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_30),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_3),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_60),
.A2(n_16),
.B(n_26),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_53),
.B(n_64),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_70),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_92),
.B(n_9),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_47),
.B(n_16),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_15),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_98),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_15),
.B1(n_4),
.B2(n_5),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_3),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_4),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_7),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_45),
.B(n_5),
.C(n_6),
.Y(n_101)
);

NOR2x1_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_55),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_104),
.B(n_120),
.Y(n_136)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_127),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_112),
.B1(n_117),
.B2(n_122),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_111),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_62),
.B(n_58),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_52),
.B(n_64),
.C(n_65),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_5),
.B(n_6),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_115),
.B(n_99),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_80),
.A2(n_65),
.B1(n_49),
.B2(n_8),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_6),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_123),
.B(n_126),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_9),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_10),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_120),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_11),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_110),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

AOI221xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_115),
.B1(n_125),
.B2(n_98),
.C(n_117),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_77),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_150),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_77),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_127),
.A2(n_86),
.B1(n_83),
.B2(n_91),
.Y(n_139)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

CKINVDCx12_ASAP7_75t_R g140 ( 
.A(n_104),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_144),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_102),
.A2(n_91),
.B1(n_89),
.B2(n_74),
.Y(n_143)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_128),
.B(n_75),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_148),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_110),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_147),
.Y(n_167)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_151),
.A2(n_119),
.B(n_125),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_148),
.A2(n_102),
.B1(n_109),
.B2(n_121),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_130),
.B1(n_131),
.B2(n_96),
.Y(n_179)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_157),
.A2(n_165),
.B(n_131),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_121),
.C(n_113),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_161),
.C(n_113),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_149),
.C(n_151),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_129),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_162),
.Y(n_174)
);

AOI221xp5_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_150),
.B1(n_133),
.B2(n_134),
.C(n_137),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_122),
.B(n_72),
.C(n_76),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_173),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_166),
.A2(n_135),
.B(n_146),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_172),
.B1(n_177),
.B2(n_165),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_143),
.B(n_136),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_175),
.C(n_182),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_155),
.B1(n_168),
.B2(n_161),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_155),
.A2(n_130),
.B(n_139),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_179),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_167),
.B(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_159),
.B(n_142),
.Y(n_181)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

AO221x1_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_156),
.B1(n_141),
.B2(n_116),
.C(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_185),
.Y(n_199)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_176),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_187),
.A2(n_188),
.B1(n_173),
.B2(n_153),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_164),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_192),
.A2(n_154),
.B1(n_177),
.B2(n_175),
.Y(n_194)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

NOR3xp33_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_174),
.C(n_178),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_195),
.B(n_201),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_200),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_182),
.C(n_160),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_197),
.B(n_198),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_172),
.C(n_171),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_164),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_157),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_191),
.B(n_193),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_202),
.A2(n_138),
.B(n_183),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_199),
.A2(n_183),
.B1(n_189),
.B2(n_187),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_208),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_200),
.C(n_201),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_211),
.Y(n_213)
);

AOI322xp5_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_195),
.A3(n_107),
.B1(n_101),
.B2(n_49),
.C1(n_114),
.C2(n_74),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_207),
.A2(n_76),
.B(n_114),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_212),
.A2(n_203),
.B(n_208),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_214),
.A2(n_206),
.B(n_13),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_74),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_11),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_217),
.B1(n_84),
.B2(n_13),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_217),
.A2(n_213),
.B(n_206),
.Y(n_218)
);

NAND2xp33_ASAP7_75t_R g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_84),
.Y(n_221)
);


endmodule