module fake_jpeg_21190_n_302 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_302);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_265;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_23),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_11),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_30),
.Y(n_46)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_39),
.B(n_37),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_47),
.A2(n_30),
.B(n_22),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_41),
.B1(n_33),
.B2(n_24),
.Y(n_69)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_62),
.B(n_73),
.Y(n_117)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_63),
.B(n_67),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_21),
.B(n_33),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_64),
.A2(n_104),
.B(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_25),
.B(n_33),
.C(n_13),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_68),
.B(n_79),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_69),
.A2(n_78),
.B1(n_86),
.B2(n_91),
.Y(n_127)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_70),
.B(n_81),
.Y(n_124)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_48),
.B(n_26),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_72),
.B(n_75),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_36),
.Y(n_73)
);

AO22x1_ASAP7_75t_SL g74 ( 
.A1(n_51),
.A2(n_34),
.B1(n_31),
.B2(n_35),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_97),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_26),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_45),
.B1(n_18),
.B2(n_44),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_54),
.B(n_28),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_77),
.B(n_80),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_14),
.B1(n_44),
.B2(n_29),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_59),
.B(n_24),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_27),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_36),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_92),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_38),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_96),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_50),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_85),
.B(n_89),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_35),
.B1(n_45),
.B2(n_31),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_50),
.B(n_28),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_88),
.B(n_95),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_59),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_93),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_31),
.B1(n_34),
.B2(n_42),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_42),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_47),
.B(n_29),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_38),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_48),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_27),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_98),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_47),
.A2(n_34),
.B1(n_32),
.B2(n_25),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_99),
.A2(n_18),
.B1(n_22),
.B2(n_30),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_47),
.B(n_27),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_100),
.Y(n_135)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_56),
.B(n_27),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_47),
.B(n_27),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_68),
.A2(n_32),
.B1(n_43),
.B2(n_12),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_106),
.A2(n_81),
.B1(n_61),
.B2(n_82),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_38),
.C(n_30),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_105),
.C(n_84),
.Y(n_150)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_71),
.B(n_38),
.Y(n_131)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_84),
.B(n_96),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_62),
.B(n_43),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_73),
.Y(n_146)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_137),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_138),
.A2(n_69),
.B1(n_91),
.B2(n_64),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_141),
.A2(n_154),
.B1(n_166),
.B2(n_121),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_74),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_142),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_87),
.Y(n_143)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_79),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_145),
.B(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_94),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_151),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_129),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_96),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_87),
.Y(n_152)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

AO21x1_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_163),
.B(n_131),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_108),
.A2(n_100),
.B1(n_95),
.B2(n_74),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_85),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_89),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_140),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_119),
.A2(n_102),
.B1(n_63),
.B2(n_70),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_127),
.B1(n_121),
.B2(n_110),
.Y(n_181)
);

BUFx12_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_30),
.B(n_18),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_118),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_164),
.A2(n_116),
.B(n_113),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_108),
.A2(n_90),
.B1(n_93),
.B2(n_66),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_112),
.B(n_114),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_167),
.B(n_115),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_150),
.C(n_148),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_156),
.C(n_159),
.Y(n_199)
);

OAI32xp33_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_112),
.A3(n_120),
.B1(n_122),
.B2(n_133),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_194),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_107),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_173),
.B(n_179),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_161),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_180),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_129),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_181),
.A2(n_185),
.B1(n_192),
.B2(n_125),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_183),
.A2(n_189),
.B1(n_196),
.B2(n_160),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_142),
.A2(n_127),
.B1(n_110),
.B2(n_138),
.Y(n_185)
);

FAx1_ASAP7_75t_SL g187 ( 
.A(n_167),
.B(n_152),
.CI(n_155),
.CON(n_187),
.SN(n_187)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_191),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_143),
.A2(n_137),
.B1(n_130),
.B2(n_116),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_141),
.A2(n_166),
.B1(n_144),
.B2(n_159),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_190),
.A2(n_147),
.B(n_139),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_142),
.A2(n_136),
.B1(n_113),
.B2(n_114),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_153),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_144),
.A2(n_125),
.B1(n_131),
.B2(n_123),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_186),
.Y(n_197)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_208),
.C(n_218),
.Y(n_233)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_201),
.Y(n_226)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_194),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_209),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_205),
.A2(n_206),
.B1(n_12),
.B2(n_19),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_175),
.A2(n_161),
.B1(n_147),
.B2(n_164),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_211),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_153),
.C(n_163),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_184),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_210),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_109),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_213),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_165),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_189),
.A2(n_128),
.B1(n_118),
.B2(n_124),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_162),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_183),
.A2(n_128),
.B1(n_158),
.B2(n_111),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_178),
.A2(n_162),
.B1(n_12),
.B2(n_19),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_187),
.Y(n_225)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_205),
.A2(n_174),
.B1(n_175),
.B2(n_180),
.Y(n_227)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_169),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_229),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_193),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_173),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_232),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_179),
.Y(n_232)
);

AOI322xp5_ASAP7_75t_SL g235 ( 
.A1(n_208),
.A2(n_172),
.A3(n_196),
.B1(n_192),
.B2(n_170),
.C1(n_190),
.C2(n_174),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_220),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_203),
.A2(n_168),
.B1(n_162),
.B2(n_19),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_236),
.A2(n_240),
.B1(n_17),
.B2(n_1),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_168),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_237),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_12),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_232),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_199),
.C(n_212),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_250),
.C(n_253),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_234),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_246),
.B(n_247),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_223),
.A2(n_198),
.B(n_206),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_249),
.B(n_251),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_213),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_230),
.B(n_219),
.Y(n_253)
);

OA21x2_ASAP7_75t_L g255 ( 
.A1(n_236),
.A2(n_198),
.B(n_217),
.Y(n_255)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_239),
.A2(n_207),
.B1(n_197),
.B2(n_11),
.Y(n_256)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_256),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_30),
.C(n_19),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_241),
.C(n_231),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_0),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_254),
.A2(n_239),
.B1(n_240),
.B2(n_227),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_263),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_252),
.A2(n_255),
.B1(n_242),
.B2(n_253),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_266),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_248),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_SL g267 ( 
.A1(n_255),
.A2(n_226),
.B(n_224),
.C(n_222),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_267),
.A2(n_247),
.B1(n_17),
.B2(n_2),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_250),
.B(n_252),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_222),
.C(n_17),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_244),
.C(n_17),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_271),
.A2(n_245),
.B1(n_257),
.B2(n_9),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_276),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_274),
.A2(n_260),
.B1(n_261),
.B2(n_268),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_270),
.A2(n_244),
.B(n_9),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_265),
.B(n_4),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_0),
.C(n_1),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_280),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_2),
.C(n_3),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_278),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_286),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_286),
.B1(n_267),
.B2(n_281),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_285),
.Y(n_293)
);

OAI21x1_ASAP7_75t_L g285 ( 
.A1(n_277),
.A2(n_267),
.B(n_269),
.Y(n_285)
);

O2A1O1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_277),
.A2(n_267),
.B(n_261),
.C(n_264),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_259),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_287),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_263),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_289),
.B(n_291),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_292),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_292),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_274),
.Y(n_298)
);

OAI21x1_ASAP7_75t_SL g297 ( 
.A1(n_294),
.A2(n_290),
.B(n_293),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_297),
.A2(n_298),
.B(n_295),
.Y(n_299)
);

NOR3xp33_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_3),
.C(n_4),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g301 ( 
.A(n_300),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_3),
.B(n_5),
.Y(n_302)
);


endmodule