module fake_jpeg_10421_n_200 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_200);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_6),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_34),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_28),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_60),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_17),
.B1(n_19),
.B2(n_18),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_54),
.B1(n_17),
.B2(n_35),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_55),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_17),
.B1(n_19),
.B2(n_18),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_19),
.B(n_25),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_17),
.B1(n_28),
.B2(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_30),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_62),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_0),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_63),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_75),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_29),
.Y(n_70)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_74),
.B1(n_46),
.B2(n_44),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_29),
.Y(n_72)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_29),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_26),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_52),
.B(n_35),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_53),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_59),
.B1(n_62),
.B2(n_21),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_16),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_22),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_47),
.B1(n_46),
.B2(n_44),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_82),
.A2(n_74),
.B1(n_73),
.B2(n_72),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_83),
.A2(n_74),
.B1(n_67),
.B2(n_48),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_90),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_95),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_78),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_99),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_77),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_92),
.B(n_100),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_64),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_47),
.B1(n_56),
.B2(n_59),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_70),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_64),
.B1(n_76),
.B2(n_71),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_22),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_80),
.C(n_77),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_68),
.C(n_93),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_104),
.A2(n_119),
.B1(n_86),
.B2(n_94),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_107),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_112),
.Y(n_126)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_115),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_96),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_110),
.B(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_65),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_117),
.Y(n_134)
);

AOI322xp5_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_48),
.A3(n_68),
.B1(n_61),
.B2(n_81),
.C1(n_77),
.C2(n_22),
.Y(n_117)
);

AO22x1_ASAP7_75t_SL g119 ( 
.A1(n_85),
.A2(n_63),
.B1(n_30),
.B2(n_61),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_105),
.B(n_85),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_125),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_120),
.Y(n_122)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_129),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_99),
.Y(n_124)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

AO22x2_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_106),
.B1(n_116),
.B2(n_107),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_127),
.A2(n_128),
.B(n_106),
.Y(n_139)
);

NAND2x1_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_93),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_94),
.C(n_86),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_130),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_84),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_137),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_103),
.B(n_16),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_139),
.A2(n_140),
.B(n_141),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_108),
.B(n_112),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_132),
.A2(n_111),
.B(n_109),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_129),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_142),
.A2(n_148),
.B(n_134),
.Y(n_159)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

OAI321xp33_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_104),
.A3(n_111),
.B1(n_16),
.B2(n_31),
.C(n_26),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_145),
.B(n_147),
.Y(n_162)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_131),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_144),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_158),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_126),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_156),
.C(n_157),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_136),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_123),
.C(n_133),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_159),
.A2(n_162),
.B(n_154),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_143),
.A2(n_92),
.B1(n_31),
.B2(n_26),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_20),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_24),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_41),
.C(n_63),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_41),
.C(n_30),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_SL g166 ( 
.A(n_154),
.B(n_142),
.C(n_150),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_166),
.A2(n_171),
.B(n_159),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_165),
.A2(n_146),
.B1(n_164),
.B2(n_160),
.Y(n_167)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_160),
.A2(n_138),
.B1(n_24),
.B2(n_21),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_169),
.A2(n_20),
.B1(n_2),
.B2(n_3),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_170),
.B(n_27),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_155),
.C(n_156),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_174),
.A2(n_161),
.B(n_24),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_27),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_20),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_176),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_179),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_182),
.Y(n_186)
);

AOI322xp5_ASAP7_75t_L g184 ( 
.A1(n_181),
.A2(n_172),
.A3(n_173),
.B1(n_14),
.B2(n_13),
.C1(n_11),
.C2(n_7),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_157),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_1),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_184),
.A2(n_178),
.B1(n_13),
.B2(n_11),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_168),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_168),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_189),
.B(n_176),
.Y(n_190)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_190),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_191),
.B(n_193),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_188),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_192),
.A2(n_186),
.B(n_187),
.Y(n_194)
);

AOI322xp5_ASAP7_75t_L g197 ( 
.A1(n_194),
.A2(n_185),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_1),
.C2(n_7),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_198),
.B1(n_196),
.B2(n_5),
.Y(n_199)
);

AOI322xp5_ASAP7_75t_L g198 ( 
.A1(n_195),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_8),
.C1(n_188),
.C2(n_178),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_4),
.Y(n_200)
);


endmodule