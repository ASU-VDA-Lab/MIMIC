module real_jpeg_17614_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_0),
.A2(n_6),
.B1(n_42),
.B2(n_46),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_0),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_0),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_0),
.B(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_0),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_0),
.B(n_103),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_0),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_0),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_0),
.B(n_116),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_1),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_1),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_1),
.B(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_1),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_1),
.B(n_207),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_1),
.B(n_229),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_2),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_2),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_2),
.B(n_187),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_3),
.Y(n_108)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_3),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_4),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_4),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_4),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_4),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_4),
.Y(n_298)
);

AND2x4_ASAP7_75t_SL g115 ( 
.A(n_5),
.B(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_5),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_6),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_6),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_6),
.B(n_191),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_6),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_7),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_7),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_7),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_7),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_7),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_7),
.B(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_7),
.B(n_354),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_8),
.Y(n_230)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_9),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_9),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_9),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_9),
.Y(n_193)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_9),
.Y(n_336)
);

NAND2x1_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_29),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_10),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_10),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_10),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_10),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_10),
.B(n_226),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_10),
.B(n_37),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_11),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_11),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_11),
.B(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_11),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_11),
.B(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_12),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_12),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_12),
.B(n_131),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_12),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_12),
.B(n_211),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_12),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_12),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_12),
.B(n_323),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_13),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_13),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_14),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g121 ( 
.A(n_15),
.Y(n_121)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_15),
.Y(n_181)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g113 ( 
.A(n_16),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_217),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_215),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_169),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_20),
.B(n_169),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_95),
.C(n_135),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_22),
.A2(n_23),
.B1(n_95),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_62),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_24),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_40),
.C(n_50),
.Y(n_24)
);

XNOR2x2_ASAP7_75t_L g270 ( 
.A(n_25),
.B(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_28),
.B(n_33),
.C(n_36),
.Y(n_64)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_35),
.Y(n_308)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_39),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_40),
.A2(n_41),
.B1(n_50),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_41),
.A2(n_238),
.B(n_244),
.Y(n_237)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_45),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_49),
.Y(n_208)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_50),
.Y(n_272)
);

MAJx2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_56),
.C(n_59),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_51),
.A2(n_52),
.B1(n_59),
.B2(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_51),
.A2(n_52),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_56),
.B(n_140),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_59),
.Y(n_141)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_72),
.B1(n_93),
.B2(n_94),
.Y(n_62)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

XNOR2x1_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

MAJx2_ASAP7_75t_L g202 ( 
.A(n_64),
.B(n_66),
.C(n_70),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_66),
.A2(n_67),
.B1(n_231),
.B2(n_232),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_67),
.B(n_224),
.C(n_231),
.Y(n_223)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_72),
.B(n_94),
.C(n_171),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_85),
.C(n_89),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.C(n_81),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_74),
.B(n_78),
.C(n_81),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_74),
.B(n_81),
.Y(n_250)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_74),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_77),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_78),
.B(n_250),
.Y(n_249)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_80),
.Y(n_211)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_84),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_91),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_92),
.Y(n_243)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_95),
.Y(n_279)
);

XOR2x2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_123),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_109),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_97),
.B(n_109),
.C(n_124),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.C(n_105),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_98),
.A2(n_105),
.B1(n_106),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_98),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_102),
.B(n_167),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_105),
.B(n_259),
.C(n_262),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_105),
.A2(n_106),
.B1(n_259),
.B2(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_110),
.B(n_115),
.C(n_119),
.Y(n_184)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_118),
.B1(n_119),
.B2(n_122),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_115),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_115),
.A2(n_122),
.B1(n_177),
.B2(n_182),
.Y(n_176)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_120),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_125),
.B(n_130),
.C(n_132),
.Y(n_212)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_136),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_162),
.C(n_166),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_137),
.B(n_274),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.C(n_152),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2x1_ASAP7_75t_L g265 ( 
.A(n_139),
.B(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_142),
.B(n_152),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_148),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_143),
.B(n_148),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_150),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.C(n_158),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_153),
.A2(n_156),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_153),
.Y(n_255)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_156),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_156),
.A2(n_256),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_156),
.B(n_331),
.C(n_337),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_158),
.B(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_162),
.B(n_166),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_199),
.B1(n_213),
.B2(n_214),
.Y(n_172)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_173),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_183),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_177),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_180),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx6_ASAP7_75t_L g324 ( 
.A(n_188),
.Y(n_324)
);

XNOR2x1_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.Y(n_189)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_197),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_212),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_387),
.Y(n_218)
);

NAND3xp33_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_275),
.C(n_280),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_267),
.Y(n_220)
);

NOR2xp67_ASAP7_75t_SL g390 ( 
.A(n_221),
.B(n_267),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_251),
.C(n_265),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_222),
.B(n_385),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_236),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_223),
.B(n_237),
.C(n_249),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_224),
.B(n_376),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_225),
.B(n_228),
.Y(n_321)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_225),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_225),
.A2(n_340),
.B1(n_341),
.B2(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_249),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_252),
.B(n_265),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_257),
.C(n_263),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_253),
.B(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_258),
.B(n_264),
.Y(n_371)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_259),
.Y(n_317)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_262),
.B(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_273),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_270),
.C(n_273),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_276),
.Y(n_389)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_277),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_382),
.B(n_386),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_367),
.B(n_381),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_325),
.B(n_366),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_312),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g366 ( 
.A(n_284),
.B(n_312),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_299),
.C(n_306),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_286),
.B(n_362),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_288),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_290),
.C(n_294),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_294),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_299),
.A2(n_300),
.B1(n_306),
.B2(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_301),
.B(n_303),
.Y(n_338)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_306),
.Y(n_363)
);

AO22x1_ASAP7_75t_SL g306 ( 
.A1(n_307),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_306)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_307),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_309),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_310),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_311),
.B(n_353),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_318),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_314),
.B(n_318),
.C(n_380),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_315),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJx2_ASAP7_75t_L g378 ( 
.A(n_319),
.B(n_321),
.C(n_322),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_360),
.B(n_365),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_342),
.B(n_359),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_339),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_339),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_329),
.A2(n_330),
.B1(n_337),
.B2(n_338),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_341),
.Y(n_351)
);

AOI21x1_ASAP7_75t_SL g342 ( 
.A1(n_343),
.A2(n_352),
.B(n_358),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_350),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_350),
.Y(n_358)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_361),
.B(n_364),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_361),
.B(n_364),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_368),
.B(n_379),
.Y(n_367)
);

NOR2xp67_ASAP7_75t_L g381 ( 
.A(n_368),
.B(n_379),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_370),
.B1(n_372),
.B2(n_373),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_374),
.C(n_378),
.Y(n_383)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_374),
.A2(n_375),
.B1(n_377),
.B2(n_378),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_383),
.B(n_384),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.C(n_390),
.Y(n_387)
);


endmodule