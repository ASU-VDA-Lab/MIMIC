module fake_netlist_5_662_n_1163 (n_137, n_210, n_168, n_260, n_164, n_191, n_286, n_91, n_208, n_82, n_122, n_194, n_282, n_142, n_176, n_10, n_214, n_140, n_24, n_248, n_124, n_86, n_136, n_146, n_268, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_241, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_281, n_207, n_240, n_114, n_57, n_96, n_37, n_189, n_220, n_291, n_165, n_111, n_229, n_108, n_231, n_257, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_249, n_271, n_284, n_46, n_233, n_21, n_94, n_203, n_245, n_274, n_205, n_113, n_38, n_123, n_139, n_105, n_280, n_246, n_80, n_4, n_179, n_125, n_35, n_269, n_167, n_128, n_73, n_234, n_277, n_17, n_92, n_19, n_267, n_149, n_120, n_285, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_254, n_14, n_225, n_84, n_23, n_202, n_130, n_266, n_272, n_219, n_157, n_258, n_265, n_29, n_79, n_193, n_293, n_131, n_151, n_47, n_173, n_192, n_244, n_251, n_25, n_53, n_160, n_198, n_223, n_288, n_247, n_188, n_190, n_8, n_201, n_292, n_158, n_263, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_264, n_283, n_109, n_112, n_212, n_85, n_159, n_163, n_276, n_95, n_119, n_183, n_185, n_243, n_239, n_275, n_175, n_252, n_169, n_59, n_262, n_26, n_255, n_133, n_238, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_290, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_242, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_259, n_273, n_287, n_270, n_222, n_230, n_81, n_118, n_28, n_89, n_279, n_70, n_115, n_68, n_93, n_253, n_261, n_72, n_174, n_186, n_199, n_289, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_256, n_48, n_204, n_50, n_250, n_52, n_278, n_88, n_110, n_216, n_1163);

input n_137;
input n_210;
input n_168;
input n_260;
input n_164;
input n_191;
input n_286;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_282;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_268;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_241;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_281;
input n_207;
input n_240;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_291;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_257;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_249;
input n_271;
input n_284;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_245;
input n_274;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_280;
input n_246;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_269;
input n_167;
input n_128;
input n_73;
input n_234;
input n_277;
input n_17;
input n_92;
input n_19;
input n_267;
input n_149;
input n_120;
input n_285;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_254;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_266;
input n_272;
input n_219;
input n_157;
input n_258;
input n_265;
input n_29;
input n_79;
input n_193;
input n_293;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_244;
input n_251;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_288;
input n_247;
input n_188;
input n_190;
input n_8;
input n_201;
input n_292;
input n_158;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_264;
input n_283;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_276;
input n_95;
input n_119;
input n_183;
input n_185;
input n_243;
input n_239;
input n_275;
input n_175;
input n_252;
input n_169;
input n_59;
input n_262;
input n_26;
input n_255;
input n_133;
input n_238;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_290;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_242;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_259;
input n_273;
input n_287;
input n_270;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_279;
input n_70;
input n_115;
input n_68;
input n_93;
input n_253;
input n_261;
input n_72;
input n_174;
input n_186;
input n_199;
input n_289;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_256;
input n_48;
input n_204;
input n_50;
input n_250;
input n_52;
input n_278;
input n_88;
input n_110;
input n_216;

output n_1163;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_1141;
wire n_785;
wire n_316;
wire n_855;
wire n_389;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_912;
wire n_968;
wire n_315;
wire n_523;
wire n_913;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_1161;
wire n_678;
wire n_664;
wire n_697;
wire n_376;
wire n_503;
wire n_967;
wire n_1150;
wire n_605;
wire n_776;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_620;
wire n_351;
wire n_643;
wire n_367;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_1157;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_501;
wire n_823;
wire n_983;
wire n_1128;
wire n_725;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_688;
wire n_581;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_690;
wire n_1013;
wire n_583;
wire n_718;
wire n_671;
wire n_819;
wire n_302;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_372;
wire n_443;
wire n_677;
wire n_864;
wire n_859;
wire n_1110;
wire n_951;
wire n_1121;
wire n_821;
wire n_714;
wire n_447;
wire n_433;
wire n_314;
wire n_604;
wire n_368;
wire n_321;
wire n_909;
wire n_625;
wire n_949;
wire n_854;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_946;
wire n_417;
wire n_932;
wire n_1048;
wire n_612;
wire n_1001;
wire n_498;
wire n_385;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_1152;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_640;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_739;
wire n_508;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_947;
wire n_820;
wire n_936;
wire n_373;
wire n_757;
wire n_1090;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_1107;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1032;
wire n_1143;
wire n_804;
wire n_867;
wire n_1124;
wire n_537;
wire n_1158;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_756;
wire n_1145;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_394;
wire n_579;
wire n_992;
wire n_1049;
wire n_1153;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_1154;
wire n_883;
wire n_1135;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_1108;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_1016;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_918;
wire n_942;
wire n_381;
wire n_1147;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_1096;
wire n_1095;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_570;
wire n_457;
wire n_514;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_1148;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_339;
wire n_1146;
wire n_882;
wire n_398;
wire n_1149;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_1020;
wire n_662;
wire n_459;
wire n_1062;
wire n_646;
wire n_962;
wire n_400;
wire n_930;
wire n_436;
wire n_580;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_922;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_816;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_528;
wire n_479;
wire n_510;
wire n_680;
wire n_974;
wire n_395;
wire n_553;
wire n_432;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_1159;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_928;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_1151;
wire n_1134;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_517;
wire n_342;
wire n_482;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_866;
wire n_573;
wire n_796;
wire n_969;
wire n_1069;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_1061;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_477;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_770;
wire n_844;
wire n_1031;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_1028;
wire n_383;
wire n_711;
wire n_834;
wire n_781;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_1101;
wire n_585;
wire n_349;
wire n_1106;
wire n_616;
wire n_953;
wire n_601;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1116;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_1131;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_513;
wire n_425;
wire n_407;
wire n_527;
wire n_707;
wire n_710;
wire n_795;
wire n_832;
wire n_695;
wire n_857;
wire n_1072;
wire n_656;
wire n_560;
wire n_340;
wire n_1094;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_495;
wire n_487;
wire n_665;
wire n_602;
wire n_574;
wire n_437;
wire n_403;
wire n_453;
wire n_421;
wire n_879;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_1156;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_404;
wire n_686;
wire n_366;
wire n_572;
wire n_754;
wire n_712;
wire n_847;
wire n_1136;
wire n_815;
wire n_596;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_529;
wire n_735;
wire n_702;
wire n_822;
wire n_412;
wire n_679;
wire n_327;
wire n_1109;
wire n_657;
wire n_895;
wire n_644;
wire n_728;
wire n_1037;
wire n_1160;
wire n_1080;
wire n_1162;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_352;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_811;
wire n_766;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_803;
wire n_868;
wire n_1092;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_1138;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_1155;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_200),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_103),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_78),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_42),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_12),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_242),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_293),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_220),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_130),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_163),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_66),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_53),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_184),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_264),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_256),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_221),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_289),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_262),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_96),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_97),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_290),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_72),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_147),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_121),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_150),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_161),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_233),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_260),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_5),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_156),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_230),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_8),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_28),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_291),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_111),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_23),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_216),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_40),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_18),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_159),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_255),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_104),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_112),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_12),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_201),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_286),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_168),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_283),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_253),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_117),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_154),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_120),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_190),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_287),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_76),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_10),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_186),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_236),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_34),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_285),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_118),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_52),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_65),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_162),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_81),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_228),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_124),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_199),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_160),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_189),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_69),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_13),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_158),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_136),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_27),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_277),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_175),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_11),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_234),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_237),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_246),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_127),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_169),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_170),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_185),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_7),
.Y(n_380)
);

BUFx10_ASAP7_75t_L g381 ( 
.A(n_110),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_40),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_261),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_203),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_140),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_142),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_62),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_241),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_240),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_31),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_113),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_263),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_92),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_75),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_101),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_55),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_74),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_210),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_257),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_207),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_24),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_212),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_122),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_141),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_63),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_31),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_279),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_0),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_144),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_94),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_114),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_179),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_22),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_16),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_32),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_178),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_254),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_281),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g419 ( 
.A(n_5),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_205),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_232),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_244),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_93),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_134),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_128),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_24),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_98),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_250),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_271),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_165),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_208),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_282),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_231),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_21),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_85),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_34),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_79),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_204),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_82),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_50),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_173),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_229),
.Y(n_442)
);

BUFx10_ASAP7_75t_L g443 ( 
.A(n_64),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_239),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_276),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_102),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_213),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_174),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_60),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_148),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_71),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_206),
.Y(n_452)
);

CKINVDCx14_ASAP7_75t_R g453 ( 
.A(n_164),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_149),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_275),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_191),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_109),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_197),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_44),
.Y(n_459)
);

BUFx5_ASAP7_75t_L g460 ( 
.A(n_155),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_225),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_0),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_267),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_19),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_292),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_167),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_23),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_46),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_198),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_273),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_196),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_138),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_157),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_26),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_108),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_129),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_238),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_28),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_252),
.Y(n_479)
);

BUFx10_ASAP7_75t_L g480 ( 
.A(n_187),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_84),
.Y(n_481)
);

AND2x6_ASAP7_75t_L g482 ( 
.A(n_358),
.B(n_41),
.Y(n_482)
);

INVx4_ASAP7_75t_L g483 ( 
.A(n_358),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_416),
.B(n_1),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_383),
.B(n_1),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_308),
.B(n_2),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_358),
.Y(n_487)
);

BUFx8_ASAP7_75t_SL g488 ( 
.A(n_401),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_416),
.B(n_2),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_460),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_358),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_329),
.B(n_348),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_326),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_433),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_464),
.B(n_295),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_349),
.B(n_3),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_384),
.B(n_3),
.Y(n_497)
);

BUFx8_ASAP7_75t_SL g498 ( 
.A(n_297),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_369),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_372),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_433),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_353),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_433),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_433),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_353),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_391),
.B(n_4),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_403),
.B(n_4),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_436),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_476),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_464),
.B(n_6),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_409),
.B(n_6),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_303),
.B(n_472),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_294),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_382),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_303),
.B(n_7),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_472),
.B(n_8),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_476),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_476),
.Y(n_518)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_476),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_308),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_334),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_334),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_323),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_296),
.B(n_386),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_412),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_381),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_299),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_295),
.B(n_9),
.Y(n_528)
);

INVx5_ASAP7_75t_L g529 ( 
.A(n_381),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_412),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_470),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_441),
.B(n_9),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_470),
.B(n_10),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_319),
.B(n_11),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_460),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_393),
.B(n_13),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_361),
.B(n_14),
.Y(n_537)
);

BUFx12f_ASAP7_75t_L g538 ( 
.A(n_443),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_361),
.B(n_14),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_301),
.B(n_15),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_397),
.B(n_15),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_390),
.Y(n_542)
);

BUFx8_ASAP7_75t_SL g543 ( 
.A(n_309),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_413),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_415),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_434),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_327),
.Y(n_547)
);

INVx5_ASAP7_75t_L g548 ( 
.A(n_443),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_475),
.B(n_16),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_480),
.Y(n_550)
);

INVx5_ASAP7_75t_L g551 ( 
.A(n_480),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_302),
.B(n_17),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_453),
.B(n_17),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_313),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_453),
.B(n_18),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_300),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_330),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_304),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_298),
.B(n_19),
.Y(n_559)
);

BUFx8_ASAP7_75t_L g560 ( 
.A(n_436),
.Y(n_560)
);

AND2x6_ASAP7_75t_L g561 ( 
.A(n_314),
.B(n_43),
.Y(n_561)
);

BUFx12f_ASAP7_75t_L g562 ( 
.A(n_332),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_317),
.B(n_20),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_460),
.B(n_20),
.Y(n_564)
);

INVx5_ASAP7_75t_L g565 ( 
.A(n_419),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_460),
.B(n_21),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_318),
.B(n_22),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_305),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_320),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_460),
.B(n_25),
.Y(n_570)
);

NAND2xp33_ASAP7_75t_L g571 ( 
.A(n_333),
.B(n_25),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_306),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_322),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_460),
.B(n_26),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_336),
.B(n_27),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_343),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_467),
.Y(n_577)
);

BUFx8_ASAP7_75t_SL g578 ( 
.A(n_316),
.Y(n_578)
);

CKINVDCx6p67_ASAP7_75t_R g579 ( 
.A(n_324),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_346),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_347),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_352),
.Y(n_582)
);

NOR2x1_ASAP7_75t_L g583 ( 
.A(n_462),
.B(n_45),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_338),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_350),
.B(n_29),
.Y(n_585)
);

OAI22xp33_ASAP7_75t_SL g586 ( 
.A1(n_485),
.A2(n_380),
.B1(n_406),
.B2(n_366),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_524),
.B(n_354),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_494),
.Y(n_588)
);

OAI22xp33_ASAP7_75t_SL g589 ( 
.A1(n_492),
.A2(n_555),
.B1(n_553),
.B2(n_489),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_494),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_494),
.Y(n_591)
);

AO22x2_ASAP7_75t_L g592 ( 
.A1(n_510),
.A2(n_478),
.B1(n_426),
.B2(n_356),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_495),
.B(n_307),
.Y(n_593)
);

INVx8_ASAP7_75t_L g594 ( 
.A(n_498),
.Y(n_594)
);

OAI22xp33_ASAP7_75t_L g595 ( 
.A1(n_484),
.A2(n_414),
.B1(n_474),
.B2(n_408),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_528),
.A2(n_359),
.B1(n_362),
.B2(n_335),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_503),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_503),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_487),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_513),
.B(n_374),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_503),
.Y(n_601)
);

OAI22xp33_ASAP7_75t_SL g602 ( 
.A1(n_585),
.A2(n_378),
.B1(n_385),
.B2(n_375),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_537),
.A2(n_363),
.B1(n_417),
.B2(n_410),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_487),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_547),
.B(n_310),
.Y(n_605)
);

OR2x6_ASAP7_75t_L g606 ( 
.A(n_562),
.B(n_387),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_527),
.B(n_388),
.Y(n_607)
);

AO22x2_ASAP7_75t_L g608 ( 
.A1(n_486),
.A2(n_539),
.B1(n_549),
.B2(n_552),
.Y(n_608)
);

OAI22xp33_ASAP7_75t_L g609 ( 
.A1(n_529),
.A2(n_435),
.B1(n_438),
.B2(n_429),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_532),
.A2(n_465),
.B1(n_456),
.B2(n_454),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_571),
.A2(n_341),
.B1(n_312),
.B2(n_315),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_496),
.A2(n_321),
.B1(n_325),
.B2(n_311),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_491),
.Y(n_613)
);

AO22x2_ASAP7_75t_L g614 ( 
.A1(n_486),
.A2(n_459),
.B1(n_394),
.B2(n_395),
.Y(n_614)
);

OAI22xp33_ASAP7_75t_L g615 ( 
.A1(n_529),
.A2(n_389),
.B1(n_398),
.B2(n_399),
.Y(n_615)
);

OAI22xp33_ASAP7_75t_SL g616 ( 
.A1(n_507),
.A2(n_422),
.B1(n_404),
.B2(n_423),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_491),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_501),
.Y(n_618)
);

OAI22xp33_ASAP7_75t_L g619 ( 
.A1(n_529),
.A2(n_424),
.B1(n_431),
.B2(n_432),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_556),
.B(n_447),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_SL g621 ( 
.A1(n_554),
.A2(n_449),
.B1(n_450),
.B2(n_457),
.Y(n_621)
);

OAI22xp33_ASAP7_75t_L g622 ( 
.A1(n_548),
.A2(n_458),
.B1(n_461),
.B2(n_463),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_557),
.B(n_328),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_548),
.B(n_331),
.Y(n_624)
);

AO22x2_ASAP7_75t_L g625 ( 
.A1(n_549),
.A2(n_466),
.B1(n_468),
.B2(n_469),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_501),
.Y(n_626)
);

OAI22xp33_ASAP7_75t_L g627 ( 
.A1(n_548),
.A2(n_551),
.B1(n_511),
.B2(n_516),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_523),
.B(n_29),
.Y(n_628)
);

OA22x2_ASAP7_75t_L g629 ( 
.A1(n_523),
.A2(n_471),
.B1(n_473),
.B2(n_477),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_509),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_509),
.Y(n_631)
);

BUFx10_ASAP7_75t_L g632 ( 
.A(n_568),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_551),
.B(n_337),
.Y(n_633)
);

INVx8_ASAP7_75t_L g634 ( 
.A(n_543),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_551),
.B(n_339),
.Y(n_635)
);

AO22x2_ASAP7_75t_L g636 ( 
.A1(n_552),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_584),
.B(n_340),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_517),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_SL g639 ( 
.A1(n_533),
.A2(n_481),
.B1(n_479),
.B2(n_455),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_584),
.B(n_342),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_497),
.A2(n_402),
.B1(n_451),
.B2(n_448),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_517),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_506),
.A2(n_452),
.B1(n_446),
.B2(n_445),
.Y(n_643)
);

BUFx10_ASAP7_75t_L g644 ( 
.A(n_512),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_538),
.A2(n_392),
.B1(n_442),
.B2(n_440),
.Y(n_645)
);

OAI22xp33_ASAP7_75t_L g646 ( 
.A1(n_515),
.A2(n_444),
.B1(n_439),
.B2(n_437),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_518),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_518),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_526),
.Y(n_649)
);

AND2x4_ASAP7_75t_SL g650 ( 
.A(n_579),
.B(n_344),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_520),
.B(n_30),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_521),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_550),
.Y(n_653)
);

NOR2x1p5_ASAP7_75t_L g654 ( 
.A(n_575),
.B(n_345),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_521),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_540),
.A2(n_430),
.B1(n_428),
.B2(n_427),
.Y(n_656)
);

AO22x2_ASAP7_75t_L g657 ( 
.A1(n_559),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_563),
.A2(n_425),
.B1(n_421),
.B2(n_420),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_567),
.A2(n_371),
.B1(n_411),
.B2(n_407),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_561),
.A2(n_534),
.B1(n_536),
.B2(n_541),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_521),
.Y(n_661)
);

NAND3x1_ASAP7_75t_L g662 ( 
.A(n_564),
.B(n_35),
.C(n_36),
.Y(n_662)
);

OR2x6_ASAP7_75t_L g663 ( 
.A(n_493),
.B(n_37),
.Y(n_663)
);

OAI22xp33_ASAP7_75t_L g664 ( 
.A1(n_566),
.A2(n_418),
.B1(n_405),
.B2(n_400),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_522),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_522),
.Y(n_666)
);

OAI22xp33_ASAP7_75t_SL g667 ( 
.A1(n_570),
.A2(n_396),
.B1(n_379),
.B2(n_377),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_644),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_600),
.B(n_558),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_652),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_666),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_588),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_590),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_591),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_620),
.B(n_520),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_597),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_598),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_587),
.B(n_572),
.Y(n_678)
);

XOR2xp5_ASAP7_75t_L g679 ( 
.A(n_603),
.B(n_578),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_632),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_601),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_655),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_665),
.Y(n_683)
);

INVxp67_ASAP7_75t_SL g684 ( 
.A(n_613),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_661),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_599),
.Y(n_686)
);

INVxp33_ASAP7_75t_L g687 ( 
.A(n_637),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_607),
.B(n_565),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_608),
.B(n_490),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_644),
.B(n_565),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_599),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_617),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_SL g693 ( 
.A(n_596),
.B(n_482),
.Y(n_693)
);

OR2x2_ASAP7_75t_SL g694 ( 
.A(n_628),
.B(n_651),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_617),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_620),
.B(n_530),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_631),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_631),
.Y(n_698)
);

XNOR2x1_ASAP7_75t_L g699 ( 
.A(n_657),
.B(n_37),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_618),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_605),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_626),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_594),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_630),
.Y(n_704)
);

NAND2x1p5_ASAP7_75t_L g705 ( 
.A(n_654),
.B(n_583),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_593),
.B(n_640),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_638),
.Y(n_707)
);

XNOR2x2_ASAP7_75t_L g708 ( 
.A(n_657),
.B(n_574),
.Y(n_708)
);

OAI21xp5_ASAP7_75t_L g709 ( 
.A1(n_660),
.A2(n_561),
.B(n_535),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_648),
.Y(n_710)
);

INVxp33_ASAP7_75t_L g711 ( 
.A(n_639),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_589),
.B(n_565),
.Y(n_712)
);

XOR2x2_ASAP7_75t_L g713 ( 
.A(n_621),
.B(n_610),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_604),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_642),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_647),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_608),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_625),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_632),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_614),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_594),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_625),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_614),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_623),
.Y(n_724)
);

AND2x2_ASAP7_75t_SL g725 ( 
.A(n_650),
.B(n_530),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_624),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_649),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_653),
.B(n_531),
.Y(n_728)
);

XNOR2xp5_ASAP7_75t_L g729 ( 
.A(n_609),
.B(n_645),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_633),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_635),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_663),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_634),
.Y(n_733)
);

XNOR2xp5_ASAP7_75t_L g734 ( 
.A(n_667),
.B(n_351),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_634),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_656),
.B(n_531),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_663),
.Y(n_737)
);

NOR2xp67_ASAP7_75t_L g738 ( 
.A(n_612),
.B(n_641),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_611),
.B(n_522),
.Y(n_739)
);

XNOR2x2_ASAP7_75t_L g740 ( 
.A(n_636),
.B(n_499),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_629),
.Y(n_741)
);

CKINVDCx16_ASAP7_75t_R g742 ( 
.A(n_606),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_658),
.B(n_525),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_616),
.Y(n_744)
);

INVxp67_ASAP7_75t_SL g745 ( 
.A(n_662),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_636),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_606),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_602),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_592),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_592),
.Y(n_750)
);

XOR2xp5_ASAP7_75t_L g751 ( 
.A(n_586),
.B(n_355),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_664),
.B(n_483),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_659),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_643),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_706),
.B(n_500),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_701),
.B(n_646),
.Y(n_756)
);

INVx3_ASAP7_75t_SL g757 ( 
.A(n_703),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_730),
.B(n_514),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_727),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_675),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_672),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_689),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_673),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_678),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_674),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_678),
.B(n_561),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_726),
.B(n_542),
.Y(n_767)
);

INVxp67_ASAP7_75t_SL g768 ( 
.A(n_684),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_676),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_669),
.B(n_595),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_687),
.B(n_754),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_677),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_681),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_724),
.B(n_627),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_689),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_721),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_753),
.B(n_488),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_717),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_675),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_682),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_696),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_744),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_683),
.Y(n_783)
);

NAND2x1p5_ASAP7_75t_L g784 ( 
.A(n_731),
.B(n_525),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_743),
.B(n_544),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_748),
.B(n_545),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_696),
.B(n_546),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_728),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_686),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_727),
.B(n_577),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_688),
.B(n_482),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_736),
.B(n_615),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_691),
.Y(n_793)
);

INVx4_ASAP7_75t_L g794 ( 
.A(n_739),
.Y(n_794)
);

AND2x4_ASAP7_75t_SL g795 ( 
.A(n_747),
.B(n_525),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_709),
.B(n_482),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_733),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_741),
.B(n_502),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_712),
.B(n_505),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_670),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_749),
.B(n_619),
.Y(n_801)
);

OAI21x1_ASAP7_75t_L g802 ( 
.A1(n_709),
.A2(n_508),
.B(n_360),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_692),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_739),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_695),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_752),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_693),
.B(n_357),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_718),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_712),
.B(n_569),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_697),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_705),
.B(n_569),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_738),
.B(n_684),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_752),
.B(n_569),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_671),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_722),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_698),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_705),
.B(n_573),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_690),
.B(n_573),
.Y(n_818)
);

NOR2xp67_ASAP7_75t_L g819 ( 
.A(n_685),
.B(n_483),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_690),
.B(n_573),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_750),
.B(n_576),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_702),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_720),
.B(n_576),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_723),
.B(n_576),
.Y(n_824)
);

INVx4_ASAP7_75t_L g825 ( 
.A(n_704),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_735),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_693),
.B(n_580),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_714),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_715),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_668),
.B(n_622),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_746),
.B(n_580),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_711),
.B(n_364),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_725),
.B(n_365),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_745),
.B(n_580),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_764),
.B(n_745),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_778),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_763),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_759),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_804),
.B(n_729),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_759),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_804),
.B(n_713),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_804),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_804),
.B(n_737),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_763),
.Y(n_844)
);

INVx8_ASAP7_75t_L g845 ( 
.A(n_804),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_794),
.B(n_700),
.Y(n_846)
);

OR2x6_ASAP7_75t_L g847 ( 
.A(n_797),
.B(n_747),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_768),
.B(n_734),
.Y(n_848)
);

OR2x6_ASAP7_75t_L g849 ( 
.A(n_797),
.B(n_747),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_790),
.B(n_732),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_806),
.B(n_694),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_806),
.B(n_708),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_794),
.B(n_716),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_808),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_778),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_763),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_794),
.B(n_707),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_815),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_773),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_789),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_762),
.B(n_771),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_762),
.B(n_770),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_789),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_762),
.B(n_710),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_790),
.B(n_732),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_762),
.B(n_732),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_778),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_773),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_773),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_775),
.B(n_762),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_755),
.B(n_751),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_775),
.B(n_47),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_755),
.B(n_680),
.Y(n_873)
);

INVx8_ASAP7_75t_L g874 ( 
.A(n_778),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_SL g875 ( 
.A(n_776),
.B(n_719),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_793),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_760),
.Y(n_877)
);

NOR2x1_ASAP7_75t_L g878 ( 
.A(n_812),
.B(n_833),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_795),
.Y(n_879)
);

BUFx4f_ASAP7_75t_L g880 ( 
.A(n_757),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_778),
.Y(n_881)
);

INVx4_ASAP7_75t_L g882 ( 
.A(n_760),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_779),
.B(n_48),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_770),
.B(n_740),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_785),
.B(n_367),
.Y(n_885)
);

CKINVDCx11_ASAP7_75t_R g886 ( 
.A(n_757),
.Y(n_886)
);

INVx5_ASAP7_75t_L g887 ( 
.A(n_847),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_866),
.B(n_779),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_874),
.Y(n_889)
);

INVx8_ASAP7_75t_L g890 ( 
.A(n_874),
.Y(n_890)
);

NAND2x1p5_ASAP7_75t_L g891 ( 
.A(n_866),
.B(n_842),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_838),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_876),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_838),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_862),
.A2(n_796),
.B(n_827),
.Y(n_895)
);

INVx3_ASAP7_75t_SL g896 ( 
.A(n_847),
.Y(n_896)
);

BUFx2_ASAP7_75t_L g897 ( 
.A(n_840),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_850),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_874),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_865),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_847),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_839),
.B(n_834),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_883),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_851),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_849),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_883),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_876),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_849),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_866),
.Y(n_909)
);

OR2x6_ASAP7_75t_L g910 ( 
.A(n_845),
.B(n_781),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_849),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_852),
.Y(n_912)
);

INVx6_ASAP7_75t_L g913 ( 
.A(n_873),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_880),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_835),
.Y(n_915)
);

INVxp33_ASAP7_75t_SL g916 ( 
.A(n_875),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_884),
.A2(n_792),
.B1(n_785),
.B2(n_782),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_880),
.Y(n_918)
);

BUFx2_ASAP7_75t_L g919 ( 
.A(n_877),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_886),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_893),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_907),
.Y(n_922)
);

INVx5_ASAP7_75t_L g923 ( 
.A(n_890),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_900),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_897),
.Y(n_925)
);

INVx4_ASAP7_75t_L g926 ( 
.A(n_890),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_900),
.Y(n_927)
);

BUFx2_ASAP7_75t_L g928 ( 
.A(n_892),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_917),
.A2(n_861),
.B1(n_884),
.B2(n_862),
.Y(n_929)
);

CKINVDCx20_ASAP7_75t_R g930 ( 
.A(n_920),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_909),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_913),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_898),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_917),
.A2(n_861),
.B1(n_870),
.B2(n_841),
.Y(n_934)
);

CKINVDCx6p67_ASAP7_75t_R g935 ( 
.A(n_896),
.Y(n_935)
);

INVx4_ASAP7_75t_SL g936 ( 
.A(n_903),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_902),
.B(n_832),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_903),
.A2(n_848),
.B1(n_863),
.B2(n_860),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_SL g939 ( 
.A1(n_916),
.A2(n_699),
.B1(n_871),
.B2(n_777),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_915),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_912),
.B(n_799),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_L g942 ( 
.A1(n_912),
.A2(n_799),
.B1(n_786),
.B2(n_807),
.Y(n_942)
);

INVx6_ASAP7_75t_L g943 ( 
.A(n_887),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_915),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_891),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_904),
.B(n_787),
.Y(n_946)
);

BUFx10_ASAP7_75t_L g947 ( 
.A(n_888),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_903),
.A2(n_842),
.B1(n_881),
.B2(n_867),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_906),
.A2(n_904),
.B1(n_836),
.B2(n_867),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_894),
.Y(n_950)
);

NOR2x1_ASAP7_75t_L g951 ( 
.A(n_926),
.B(n_914),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_SL g952 ( 
.A1(n_929),
.A2(n_913),
.B1(n_887),
.B2(n_742),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_939),
.A2(n_937),
.B1(n_942),
.B2(n_940),
.Y(n_953)
);

NAND3xp33_ASAP7_75t_L g954 ( 
.A(n_939),
.B(n_756),
.C(n_878),
.Y(n_954)
);

OAI222xp33_ASAP7_75t_L g955 ( 
.A1(n_934),
.A2(n_679),
.B1(n_894),
.B2(n_834),
.C1(n_843),
.C2(n_885),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_921),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_930),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_950),
.A2(n_817),
.B1(n_811),
.B2(n_872),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_SL g959 ( 
.A1(n_942),
.A2(n_830),
.B(n_795),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_941),
.A2(n_817),
.B1(n_811),
.B2(n_872),
.Y(n_960)
);

OAI222xp33_ASAP7_75t_L g961 ( 
.A1(n_938),
.A2(n_809),
.B1(n_872),
.B2(n_813),
.C1(n_910),
.C2(n_883),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_946),
.A2(n_786),
.B1(n_829),
.B2(n_906),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_933),
.A2(n_786),
.B1(n_829),
.B2(n_906),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_921),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_922),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_944),
.A2(n_887),
.B1(n_919),
.B2(n_882),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_SL g967 ( 
.A1(n_928),
.A2(n_776),
.B1(n_826),
.B2(n_918),
.Y(n_967)
);

OAI222xp33_ASAP7_75t_L g968 ( 
.A1(n_933),
.A2(n_809),
.B1(n_910),
.B2(n_901),
.C1(n_784),
.C2(n_882),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_925),
.A2(n_879),
.B1(n_908),
.B2(n_905),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_925),
.A2(n_786),
.B1(n_864),
.B2(n_758),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_932),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_924),
.A2(n_864),
.B1(n_758),
.B2(n_820),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_927),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_930),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_931),
.A2(n_864),
.B1(n_820),
.B2(n_767),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_L g976 ( 
.A1(n_935),
.A2(n_767),
.B1(n_888),
.B2(n_846),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_949),
.A2(n_846),
.B1(n_857),
.B2(n_853),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_L g978 ( 
.A1(n_943),
.A2(n_857),
.B1(n_846),
.B2(n_774),
.Y(n_978)
);

BUFx4f_ASAP7_75t_SL g979 ( 
.A(n_947),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_922),
.B(n_802),
.Y(n_980)
);

OAI21xp33_ASAP7_75t_L g981 ( 
.A1(n_945),
.A2(n_826),
.B(n_787),
.Y(n_981)
);

CKINVDCx11_ASAP7_75t_R g982 ( 
.A(n_947),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_943),
.A2(n_911),
.B1(n_766),
.B2(n_854),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_936),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_943),
.A2(n_858),
.B1(n_818),
.B2(n_910),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_973),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_L g987 ( 
.A1(n_954),
.A2(n_560),
.B1(n_793),
.B2(n_816),
.Y(n_987)
);

OAI21xp33_ASAP7_75t_L g988 ( 
.A1(n_981),
.A2(n_784),
.B(n_788),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_952),
.A2(n_857),
.B1(n_816),
.B2(n_803),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_976),
.A2(n_757),
.B1(n_784),
.B2(n_923),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_967),
.A2(n_923),
.B1(n_926),
.B2(n_891),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_953),
.A2(n_886),
.B1(n_781),
.B2(n_788),
.Y(n_992)
);

OAI211xp5_ASAP7_75t_SL g993 ( 
.A1(n_971),
.A2(n_801),
.B(n_765),
.C(n_769),
.Y(n_993)
);

OAI211xp5_ASAP7_75t_L g994 ( 
.A1(n_959),
.A2(n_801),
.B(n_821),
.C(n_831),
.Y(n_994)
);

NAND3xp33_ASAP7_75t_SL g995 ( 
.A(n_957),
.B(n_805),
.C(n_803),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_983),
.A2(n_810),
.B1(n_805),
.B2(n_783),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_SL g997 ( 
.A1(n_985),
.A2(n_802),
.B1(n_923),
.B2(n_560),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_958),
.A2(n_810),
.B1(n_772),
.B2(n_761),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_960),
.A2(n_821),
.B1(n_823),
.B2(n_824),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_962),
.A2(n_923),
.B1(n_836),
.B2(n_881),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_975),
.A2(n_772),
.B1(n_780),
.B2(n_761),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_SL g1002 ( 
.A1(n_966),
.A2(n_895),
.B1(n_947),
.B2(n_845),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_973),
.B(n_956),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_964),
.B(n_895),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_965),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_970),
.A2(n_824),
.B1(n_823),
.B2(n_831),
.Y(n_1006)
);

NAND2xp33_ASAP7_75t_SL g1007 ( 
.A(n_957),
.B(n_889),
.Y(n_1007)
);

AOI222xp33_ASAP7_75t_L g1008 ( 
.A1(n_955),
.A2(n_798),
.B1(n_765),
.B2(n_769),
.C1(n_814),
.C2(n_800),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_L g1009 ( 
.A1(n_972),
.A2(n_780),
.B1(n_783),
.B2(n_828),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_978),
.A2(n_828),
.B1(n_814),
.B2(n_800),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_963),
.A2(n_977),
.B1(n_979),
.B2(n_951),
.Y(n_1011)
);

NAND3xp33_ASAP7_75t_L g1012 ( 
.A(n_969),
.B(n_370),
.C(n_368),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_982),
.A2(n_825),
.B1(n_845),
.B2(n_822),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_982),
.A2(n_825),
.B1(n_822),
.B2(n_855),
.Y(n_1014)
);

AOI22xp33_ASAP7_75t_SL g1015 ( 
.A1(n_974),
.A2(n_890),
.B1(n_948),
.B2(n_855),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_974),
.A2(n_825),
.B1(n_791),
.B2(n_837),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_980),
.A2(n_984),
.B1(n_844),
.B2(n_837),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_980),
.B(n_936),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_984),
.B(n_936),
.Y(n_1019)
);

OAI222xp33_ASAP7_75t_L g1020 ( 
.A1(n_961),
.A2(n_373),
.B1(n_376),
.B2(n_869),
.C1(n_868),
.C2(n_859),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_968),
.A2(n_582),
.B1(n_581),
.B2(n_869),
.Y(n_1021)
);

NAND3xp33_ASAP7_75t_L g1022 ( 
.A(n_954),
.B(n_581),
.C(n_582),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_954),
.A2(n_581),
.B1(n_582),
.B2(n_868),
.Y(n_1023)
);

NAND4xp25_ASAP7_75t_L g1024 ( 
.A(n_987),
.B(n_798),
.C(n_504),
.D(n_38),
.Y(n_1024)
);

OAI221xp5_ASAP7_75t_SL g1025 ( 
.A1(n_992),
.A2(n_38),
.B1(n_39),
.B2(n_859),
.C(n_856),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1003),
.B(n_39),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_987),
.A2(n_988),
.B1(n_990),
.B2(n_1012),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_994),
.B(n_889),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_986),
.B(n_49),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_1005),
.B(n_51),
.Y(n_1030)
);

NAND3xp33_ASAP7_75t_L g1031 ( 
.A(n_1008),
.B(n_856),
.C(n_844),
.Y(n_1031)
);

AOI22xp33_ASAP7_75t_L g1032 ( 
.A1(n_1011),
.A2(n_899),
.B1(n_889),
.B2(n_819),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_1018),
.B(n_54),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1004),
.B(n_504),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_989),
.B(n_56),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_1021),
.A2(n_899),
.B1(n_819),
.B2(n_519),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1019),
.B(n_57),
.Y(n_1037)
);

NAND3xp33_ASAP7_75t_L g1038 ( 
.A(n_993),
.B(n_899),
.C(n_519),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_997),
.B(n_58),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1023),
.B(n_59),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1023),
.B(n_61),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1017),
.B(n_67),
.Y(n_1042)
);

NOR3xp33_ASAP7_75t_L g1043 ( 
.A(n_995),
.B(n_68),
.C(n_70),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_1022),
.B(n_519),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1021),
.B(n_1002),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_991),
.B(n_73),
.Y(n_1046)
);

NAND3xp33_ASAP7_75t_L g1047 ( 
.A(n_1016),
.B(n_77),
.C(n_80),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_1015),
.B(n_83),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_996),
.Y(n_1049)
);

OAI221xp5_ASAP7_75t_L g1050 ( 
.A1(n_1013),
.A2(n_1006),
.B1(n_999),
.B2(n_1014),
.C(n_1010),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1007),
.B(n_86),
.Y(n_1051)
);

AOI21xp33_ASAP7_75t_L g1052 ( 
.A1(n_1000),
.A2(n_87),
.B(n_88),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_998),
.B(n_89),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_1001),
.B(n_90),
.Y(n_1054)
);

AOI221xp5_ASAP7_75t_L g1055 ( 
.A1(n_1025),
.A2(n_1020),
.B1(n_1009),
.B2(n_99),
.C(n_100),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1026),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_1034),
.B(n_91),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_1033),
.B(n_95),
.Y(n_1058)
);

OAI211xp5_ASAP7_75t_SL g1059 ( 
.A1(n_1027),
.A2(n_105),
.B(n_106),
.C(n_107),
.Y(n_1059)
);

NOR2x1_ASAP7_75t_L g1060 ( 
.A(n_1038),
.B(n_115),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1049),
.B(n_116),
.Y(n_1061)
);

AOI22xp33_ASAP7_75t_L g1062 ( 
.A1(n_1024),
.A2(n_119),
.B1(n_123),
.B2(n_125),
.Y(n_1062)
);

NAND3xp33_ASAP7_75t_L g1063 ( 
.A(n_1039),
.B(n_126),
.C(n_131),
.Y(n_1063)
);

NAND3xp33_ASAP7_75t_L g1064 ( 
.A(n_1039),
.B(n_132),
.C(n_133),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1029),
.Y(n_1065)
);

NAND4xp75_ASAP7_75t_L g1066 ( 
.A(n_1028),
.B(n_1048),
.C(n_1046),
.D(n_1053),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1028),
.B(n_135),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1029),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1037),
.B(n_137),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_1030),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_1045),
.B(n_139),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_1030),
.B(n_1048),
.Y(n_1072)
);

NAND3xp33_ASAP7_75t_L g1073 ( 
.A(n_1043),
.B(n_1047),
.C(n_1053),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1032),
.B(n_143),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_1051),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1042),
.B(n_145),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1068),
.B(n_1042),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1065),
.Y(n_1078)
);

NAND4xp75_ASAP7_75t_SL g1079 ( 
.A(n_1066),
.B(n_1054),
.C(n_1058),
.D(n_1069),
.Y(n_1079)
);

XNOR2xp5_ASAP7_75t_L g1080 ( 
.A(n_1072),
.B(n_1050),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1056),
.B(n_1044),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1072),
.B(n_1054),
.Y(n_1082)
);

XNOR2xp5_ASAP7_75t_L g1083 ( 
.A(n_1063),
.B(n_1031),
.Y(n_1083)
);

INVx3_ASAP7_75t_SL g1084 ( 
.A(n_1071),
.Y(n_1084)
);

XNOR2xp5_ASAP7_75t_L g1085 ( 
.A(n_1063),
.B(n_1035),
.Y(n_1085)
);

NAND4xp75_ASAP7_75t_L g1086 ( 
.A(n_1055),
.B(n_1052),
.C(n_1041),
.D(n_1040),
.Y(n_1086)
);

NAND4xp75_ASAP7_75t_SL g1087 ( 
.A(n_1073),
.B(n_1036),
.C(n_1044),
.D(n_152),
.Y(n_1087)
);

OA22x2_ASAP7_75t_L g1088 ( 
.A1(n_1067),
.A2(n_146),
.B1(n_151),
.B2(n_153),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1070),
.B(n_166),
.Y(n_1089)
);

NAND3xp33_ASAP7_75t_L g1090 ( 
.A(n_1064),
.B(n_171),
.C(n_172),
.Y(n_1090)
);

CKINVDCx14_ASAP7_75t_R g1091 ( 
.A(n_1075),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1067),
.Y(n_1092)
);

NOR3xp33_ASAP7_75t_L g1093 ( 
.A(n_1073),
.B(n_176),
.C(n_177),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1064),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_1094)
);

NAND4xp75_ASAP7_75t_L g1095 ( 
.A(n_1060),
.B(n_183),
.C(n_188),
.D(n_192),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1057),
.B(n_193),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1078),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1092),
.B(n_1061),
.Y(n_1098)
);

INVxp67_ASAP7_75t_L g1099 ( 
.A(n_1081),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1081),
.B(n_1076),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1077),
.Y(n_1101)
);

BUFx12f_ASAP7_75t_L g1102 ( 
.A(n_1096),
.Y(n_1102)
);

XNOR2x2_ASAP7_75t_L g1103 ( 
.A(n_1083),
.B(n_1074),
.Y(n_1103)
);

OAI22x1_ASAP7_75t_L g1104 ( 
.A1(n_1080),
.A2(n_1062),
.B1(n_1059),
.B2(n_202),
.Y(n_1104)
);

XNOR2x2_ASAP7_75t_L g1105 ( 
.A(n_1090),
.B(n_194),
.Y(n_1105)
);

XNOR2xp5_ASAP7_75t_L g1106 ( 
.A(n_1079),
.B(n_288),
.Y(n_1106)
);

INVxp67_ASAP7_75t_L g1107 ( 
.A(n_1082),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1091),
.B(n_195),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1084),
.Y(n_1109)
);

INVx5_ASAP7_75t_L g1110 ( 
.A(n_1089),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1085),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_1088),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1088),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1090),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_1086),
.B(n_209),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1114),
.A2(n_1093),
.B1(n_1094),
.B2(n_1095),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1097),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1099),
.Y(n_1118)
);

XOR2xp5_ASAP7_75t_L g1119 ( 
.A(n_1103),
.B(n_1087),
.Y(n_1119)
);

AOI22x1_ASAP7_75t_L g1120 ( 
.A1(n_1112),
.A2(n_1113),
.B1(n_1104),
.B2(n_1106),
.Y(n_1120)
);

XOR2x2_ASAP7_75t_L g1121 ( 
.A(n_1111),
.B(n_1087),
.Y(n_1121)
);

XOR2x2_ASAP7_75t_L g1122 ( 
.A(n_1105),
.B(n_211),
.Y(n_1122)
);

INVx1_ASAP7_75t_SL g1123 ( 
.A(n_1108),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1098),
.Y(n_1124)
);

OAI22x1_ASAP7_75t_L g1125 ( 
.A1(n_1112),
.A2(n_214),
.B1(n_215),
.B2(n_217),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1098),
.Y(n_1126)
);

OA22x2_ASAP7_75t_L g1127 ( 
.A1(n_1109),
.A2(n_1107),
.B1(n_1100),
.B2(n_1101),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1115),
.A2(n_218),
.B1(n_219),
.B2(n_222),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1107),
.Y(n_1129)
);

OA22x2_ASAP7_75t_L g1130 ( 
.A1(n_1100),
.A2(n_223),
.B1(n_224),
.B2(n_226),
.Y(n_1130)
);

INVx5_ASAP7_75t_L g1131 ( 
.A(n_1110),
.Y(n_1131)
);

OA22x2_ASAP7_75t_SL g1132 ( 
.A1(n_1110),
.A2(n_227),
.B1(n_235),
.B2(n_243),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1110),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_1131),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1117),
.Y(n_1135)
);

INVxp67_ASAP7_75t_SL g1136 ( 
.A(n_1119),
.Y(n_1136)
);

BUFx2_ASAP7_75t_SL g1137 ( 
.A(n_1131),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_1131),
.Y(n_1138)
);

AO22x2_ASAP7_75t_L g1139 ( 
.A1(n_1136),
.A2(n_1119),
.B1(n_1133),
.B2(n_1129),
.Y(n_1139)
);

OAI22x1_ASAP7_75t_L g1140 ( 
.A1(n_1134),
.A2(n_1120),
.B1(n_1116),
.B2(n_1123),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1138),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1137),
.A2(n_1122),
.B1(n_1127),
.B2(n_1130),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1135),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1139),
.A2(n_1137),
.B1(n_1118),
.B2(n_1138),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1143),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1141),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_1140),
.Y(n_1147)
);

AO22x2_ASAP7_75t_L g1148 ( 
.A1(n_1146),
.A2(n_1138),
.B1(n_1135),
.B2(n_1126),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1147),
.A2(n_1142),
.B1(n_1121),
.B2(n_1124),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1145),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1144),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1149),
.A2(n_1125),
.B1(n_1128),
.B2(n_1102),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1148),
.Y(n_1153)
);

AND5x1_ASAP7_75t_L g1154 ( 
.A(n_1152),
.B(n_1151),
.C(n_1132),
.D(n_1150),
.E(n_248),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_1154),
.Y(n_1155)
);

OAI22x1_ASAP7_75t_L g1156 ( 
.A1(n_1155),
.A2(n_1153),
.B1(n_245),
.B2(n_247),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1156),
.Y(n_1157)
);

AO22x1_ASAP7_75t_L g1158 ( 
.A1(n_1157),
.A2(n_249),
.B1(n_251),
.B2(n_258),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1158),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1159),
.A2(n_259),
.B1(n_265),
.B2(n_266),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1160),
.Y(n_1161)
);

AOI221xp5_ASAP7_75t_L g1162 ( 
.A1(n_1161),
.A2(n_268),
.B1(n_270),
.B2(n_272),
.C(n_274),
.Y(n_1162)
);

AOI211xp5_ASAP7_75t_L g1163 ( 
.A1(n_1162),
.A2(n_278),
.B(n_280),
.C(n_284),
.Y(n_1163)
);


endmodule