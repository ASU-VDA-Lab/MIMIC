module real_jpeg_2832_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx2_ASAP7_75t_L g104 ( 
.A(n_0),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_1),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_2),
.B(n_26),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_2),
.B(n_38),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_2),
.B(n_31),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_2),
.B(n_49),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_2),
.B(n_61),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_3),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_3),
.B(n_38),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_3),
.B(n_31),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_3),
.B(n_49),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_4),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_4),
.B(n_38),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_4),
.B(n_31),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g80 ( 
.A(n_7),
.Y(n_80)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_9),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_9),
.B(n_26),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_9),
.B(n_61),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_10),
.B(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_10),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_10),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_10),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_10),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_10),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_10),
.B(n_26),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_26),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_12),
.B(n_31),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_12),
.B(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_12),
.B(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_12),
.B(n_61),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_12),
.B(n_102),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_12),
.B(n_124),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_13),
.B(n_26),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_13),
.B(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_13),
.B(n_31),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_13),
.B(n_61),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_13),
.B(n_49),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_13),
.B(n_102),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_13),
.B(n_80),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_13),
.B(n_124),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_14),
.B(n_26),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_14),
.B(n_38),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_14),
.B(n_31),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_14),
.B(n_49),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_14),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_14),
.B(n_102),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI31xp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_25),
.A3(n_162),
.B(n_322),
.Y(n_17)
);

OAI211xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_42),
.B(n_88),
.C(n_321),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_63),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_21),
.B(n_63),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_50),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_42),
.B2(n_43),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B1(n_29),
.B2(n_41),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_25),
.B(n_74),
.C(n_75),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_25),
.A2(n_41),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_26),
.Y(n_196)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_34),
.B(n_40),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_34),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_44),
.C(n_47),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_30),
.A2(n_47),
.B1(n_48),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_30),
.B(n_192),
.C(n_199),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_30),
.A2(n_54),
.B1(n_199),
.B2(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_31),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_34),
.A2(n_35),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_35),
.B(n_101),
.C(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_37),
.B(n_166),
.Y(n_165)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_40),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_45),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_44),
.A2(n_45),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_45),
.B(n_113),
.C(n_115),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_48),
.B1(n_59),
.B2(n_60),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_47),
.A2(n_48),
.B1(n_185),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_57),
.C(n_59),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_48),
.B(n_114),
.C(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_SL g219 ( 
.A(n_49),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_55),
.C(n_56),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_56),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_57),
.A2(n_58),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_59),
.A2(n_60),
.B1(n_78),
.B2(n_79),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_59),
.A2(n_60),
.B1(n_107),
.B2(n_147),
.Y(n_277)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_78),
.C(n_81),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_60),
.B(n_107),
.C(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_61),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_85),
.C(n_86),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_64),
.A2(n_65),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_77),
.C(n_82),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_66),
.A2(n_67),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_73),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_72),
.C(n_73),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_69),
.A2(n_70),
.B1(n_125),
.B2(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_69),
.A2(n_70),
.B1(n_170),
.B2(n_171),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_70),
.B(n_121),
.C(n_125),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_70),
.B(n_164),
.C(n_170),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_74),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_74),
.B(n_165),
.C(n_167),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_74),
.A2(n_118),
.B1(n_165),
.B2(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_77),
.B(n_82),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_79),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_SL g132 ( 
.A(n_78),
.B(n_96),
.C(n_100),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_78),
.A2(n_79),
.B1(n_256),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_79),
.B(n_256),
.C(n_257),
.Y(n_255)
);

INVx13_ASAP7_75t_L g227 ( 
.A(n_80),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_81),
.B(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_85),
.B(n_86),
.Y(n_318)
);

A2O1A1O1Ixp25_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_200),
.B(n_312),
.C(n_315),
.D(n_320),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_172),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_90),
.A2(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_138),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_91),
.B(n_138),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_126),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_92),
.B(n_127),
.C(n_137),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_116),
.C(n_120),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_93),
.B(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_105),
.C(n_109),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_94),
.A2(n_95),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_100),
.A2(n_101),
.B1(n_123),
.B2(n_153),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_105),
.B(n_109),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.C(n_108),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_106),
.B(n_108),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_113),
.A2(n_114),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_121),
.A2(n_122),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_152),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_123),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_183)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_124),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_125),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_126)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.C(n_132),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_128),
.A2(n_129),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_131),
.B(n_132),
.Y(n_142)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.C(n_144),
.Y(n_138)
);

FAx1_ASAP7_75t_SL g173 ( 
.A(n_139),
.B(n_141),
.CI(n_144),
.CON(n_173),
.SN(n_173)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_159),
.C(n_163),
.Y(n_144)
);

FAx1_ASAP7_75t_SL g175 ( 
.A(n_145),
.B(n_159),
.CI(n_163),
.CON(n_175),
.SN(n_175)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.C(n_156),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_146),
.B(n_150),
.Y(n_237)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_153),
.B(n_154),
.C(n_155),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_151),
.B(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_151),
.A2(n_152),
.B1(n_253),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_154),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_155),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_156),
.B(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_166),
.B(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_166),
.B(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_169),
.B(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_169),
.B(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_173),
.B(n_174),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_173),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.C(n_179),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_175),
.B(n_176),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_175),
.Y(n_327)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_177),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_179),
.B(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_189),
.C(n_191),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_180),
.A2(n_181),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.C(n_186),
.Y(n_181)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_182),
.B(n_184),
.CI(n_186),
.CON(n_266),
.SN(n_266)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_185),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_189),
.B(n_191),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_192),
.A2(n_193),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.C(n_198),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_197),
.A2(n_198),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_197),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_198),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_199),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_267),
.B(n_306),
.C(n_307),
.D(n_311),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_242),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_203),
.B(n_242),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_234),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_204),
.B(n_235),
.C(n_241),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_222),
.C(n_230),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_205),
.A2(n_206),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_211),
.C(n_215),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_207),
.B(n_298),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_211),
.A2(n_212),
.B1(n_215),
.B2(n_299),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_212),
.A2(n_213),
.B(n_214),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_215),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.C(n_220),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_216),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_250),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_222),
.B(n_230),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.C(n_228),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_224),
.B(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_228),
.Y(n_259)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_238),
.B2(n_241),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_239),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.C(n_265),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_243),
.A2(n_265),
.B1(n_266),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_243),
.Y(n_303)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_246),
.B(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_258),
.C(n_260),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_247),
.B(n_294),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_251),
.C(n_255),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_248),
.A2(n_249),
.B1(n_279),
.B2(n_281),
.Y(n_278)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_251),
.A2(n_252),
.B1(n_255),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_253),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_255),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_256),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_258),
.A2(n_260),
.B1(n_261),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_258),
.Y(n_295)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_266),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_300),
.B(n_305),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_292),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_278),
.C(n_282),
.Y(n_269)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_270),
.Y(n_328)
);

FAx1_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_275),
.CI(n_276),
.CON(n_270),
.SN(n_270)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_275),
.C(n_276),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.C(n_274),
.Y(n_271)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_279),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.C(n_290),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.C(n_289),
.Y(n_286)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_292),
.Y(n_325)
);

FAx1_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_296),
.CI(n_297),
.CON(n_292),
.SN(n_292)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_296),
.C(n_297),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_304),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_304),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_309),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_317),
.Y(n_320)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_318),
.Y(n_319)
);


endmodule