module real_jpeg_12465_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_216;
wire n_213;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g83 ( 
.A(n_2),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_3),
.A2(n_63),
.B1(n_65),
.B2(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_3),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_4),
.B(n_44),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_4),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_4),
.B(n_136),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_4),
.A2(n_36),
.B1(n_37),
.B2(n_100),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_4),
.B(n_65),
.C(n_83),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_4),
.B(n_35),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_4),
.A2(n_67),
.B(n_164),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_4),
.A2(n_27),
.B(n_34),
.C(n_191),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_100),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_5),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_62)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_66),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_7),
.A2(n_63),
.B1(n_65),
.B2(n_72),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_7),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_7),
.A2(n_36),
.B1(n_37),
.B2(n_72),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_46),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_46),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_9),
.A2(n_46),
.B1(n_63),
.B2(n_65),
.Y(n_170)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_11),
.A2(n_29),
.B1(n_44),
.B2(n_45),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_11),
.A2(n_29),
.B1(n_63),
.B2(n_65),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_11),
.A2(n_29),
.B1(n_36),
.B2(n_37),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_48),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_12),
.B(n_28),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_13),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_80),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_13),
.A2(n_63),
.B1(n_65),
.B2(n_80),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_14),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_14),
.A2(n_36),
.B1(n_37),
.B2(n_41),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_14),
.A2(n_41),
.B1(n_63),
.B2(n_65),
.Y(n_165)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_16),
.A2(n_63),
.B1(n_65),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_16),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_124),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_122),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_102),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_20),
.B(n_102),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.C(n_88),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_21),
.A2(n_22),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_56),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_42),
.B2(n_55),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_24),
.B(n_55),
.C(n_56),
.Y(n_121)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B(n_39),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_26),
.A2(n_30),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

AOI32xp33_ASAP7_75t_L g58 ( 
.A1(n_27),
.A2(n_45),
.A3(n_48),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_30),
.A2(n_39),
.B(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_31),
.B(n_40),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_35),
.Y(n_31)
);

AO22x1_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_33),
.A2(n_36),
.B(n_100),
.Y(n_191)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_36),
.A2(n_37),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_37),
.B(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_47),
.B(n_49),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_43),
.A2(n_47),
.B1(n_51),
.B2(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_45),
.A2(n_51),
.B(n_100),
.C(n_101),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_47),
.B(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_47),
.B(n_54),
.Y(n_98)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_47),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_61),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_57),
.A2(n_58),
.B1(n_61),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_67),
.B1(n_70),
.B2(n_73),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_62),
.A2(n_67),
.B1(n_73),
.B2(n_138),
.Y(n_137)
);

INVx5_ASAP7_75t_SL g65 ( 
.A(n_63),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_63),
.B(n_69),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_65),
.B1(n_83),
.B2(n_84),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_63),
.B(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_67),
.A2(n_73),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_67),
.A2(n_163),
.B(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_69),
.B1(n_71),
.B2(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_68),
.A2(n_69),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_68),
.B(n_165),
.Y(n_178)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_69),
.B(n_165),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_73),
.A2(n_170),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_73),
.B(n_100),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_73),
.A2(n_138),
.B(n_178),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_74),
.B(n_88),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_75),
.B(n_78),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_76),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_86),
.B1(n_87),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_81),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_81),
.A2(n_87),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_85),
.A2(n_90),
.B(n_91),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_85),
.A2(n_91),
.B(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_85),
.B(n_100),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_87),
.B(n_92),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.C(n_96),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_89),
.B(n_93),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_94),
.A2(n_95),
.B(n_119),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_95),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_97),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_121),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_113),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_120),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_142),
.B(n_222),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_139),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_126),
.B(n_139),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.C(n_132),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_127),
.B(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_130),
.B(n_132),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.C(n_137),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_133),
.B(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_134),
.A2(n_135),
.B1(n_137),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_137),
.Y(n_208)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_217),
.B(n_221),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_202),
.B(n_216),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_186),
.B(n_201),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_166),
.B(n_185),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_155),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_147),
.B(n_155),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_153),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_148),
.A2(n_149),
.B1(n_153),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_151),
.B(n_152),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_150),
.A2(n_152),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_162),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_160),
.C(n_162),
.Y(n_187)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_163),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_174),
.B(n_184),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_172),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_168),
.B(n_172),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_179),
.B(n_183),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_176),
.B(n_177),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_187),
.B(n_188),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_196),
.C(n_200),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_192),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_196),
.B1(n_199),
.B2(n_200),
.Y(n_193)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_194),
.Y(n_200)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_196),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_198),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_203),
.B(n_204),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_212),
.C(n_214),
.Y(n_218)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_218),
.B(n_219),
.Y(n_221)
);


endmodule