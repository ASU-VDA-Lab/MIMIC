module fake_jpeg_10941_n_178 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_178);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx11_ASAP7_75t_SL g74 ( 
.A(n_27),
.Y(n_74)
);

INVx5_ASAP7_75t_SL g75 ( 
.A(n_74),
.Y(n_75)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_79),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_58),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_79)
);

NAND2x1_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_58),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_51),
.B(n_5),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_83),
.Y(n_98)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_60),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_6),
.C(n_7),
.Y(n_117)
);

AO22x1_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_62),
.B1(n_70),
.B2(n_57),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_54),
.B1(n_71),
.B2(n_61),
.Y(n_105)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_92),
.B(n_5),
.Y(n_114)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g100 ( 
.A(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_77),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_107),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_80),
.B1(n_61),
.B2(n_59),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_105),
.B1(n_111),
.B2(n_47),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_83),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_63),
.C(n_53),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_49),
.B1(n_69),
.B2(n_52),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_74),
.B1(n_67),
.B2(n_65),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_120),
.B1(n_72),
.B2(n_68),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_72),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_113),
.B(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_6),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_25),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_7),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_121),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_89),
.A2(n_68),
.B1(n_56),
.B2(n_48),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_131),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_128),
.B(n_133),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_119),
.B(n_8),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_132),
.B(n_135),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_8),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_9),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_56),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_136),
.A2(n_144),
.B(n_30),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_9),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_137),
.B(n_143),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_106),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_141),
.B1(n_41),
.B2(n_34),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_103),
.A2(n_10),
.B1(n_11),
.B2(n_15),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_16),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_142),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_149),
.Y(n_161)
);

NAND4xp25_ASAP7_75t_SL g149 ( 
.A(n_130),
.B(n_17),
.C(n_18),
.D(n_19),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_129),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_158),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_21),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_152),
.C(n_123),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_24),
.C(n_28),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_159),
.B(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_165),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_125),
.B(n_138),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_164),
.A2(n_166),
.B(n_147),
.Y(n_168)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_131),
.C(n_139),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_168),
.B(n_169),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_161),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_163),
.C(n_160),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_173),
.B(n_172),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_154),
.A3(n_170),
.B1(n_153),
.B2(n_134),
.C1(n_145),
.C2(n_155),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_175),
.B(n_151),
.Y(n_176)
);

NOR4xp25_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_145),
.C(n_149),
.D(n_152),
.Y(n_177)
);

HAxp5_ASAP7_75t_SL g178 ( 
.A(n_177),
.B(n_32),
.CON(n_178),
.SN(n_178)
);


endmodule