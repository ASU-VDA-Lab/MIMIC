module fake_ibex_1358_n_981 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_182, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_981);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_182;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_981;

wire n_599;
wire n_822;
wire n_778;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_947;
wire n_972;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_375;
wire n_340;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_980;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_560;
wire n_429;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_392;
wire n_206;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_444;
wire n_564;
wire n_562;
wire n_506;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_615;
wire n_512;
wire n_950;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_499;
wire n_227;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_899;
wire n_843;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_379;
wire n_288;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_385;
wire n_233;
wire n_342;
wire n_414;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_912;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_298;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_72),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_22),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_33),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_88),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_45),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_13),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_34),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_9),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_39),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_96),
.Y(n_194)
);

INVxp67_ASAP7_75t_SL g195 ( 
.A(n_81),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_85),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_106),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_121),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_61),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_133),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_153),
.Y(n_202)
);

NOR2xp67_ASAP7_75t_L g203 ( 
.A(n_56),
.B(n_50),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_117),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_6),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_14),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_34),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_139),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_152),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_155),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_60),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_69),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_18),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_84),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_87),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_161),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_86),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_99),
.B(n_163),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_127),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_116),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_55),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_31),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_79),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_140),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_120),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_17),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_78),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_162),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_113),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_136),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_21),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_114),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_33),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_38),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_119),
.Y(n_238)
);

INVxp33_ASAP7_75t_L g239 ( 
.A(n_19),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_37),
.Y(n_240)
);

INVxp67_ASAP7_75t_SL g241 ( 
.A(n_16),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_145),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_47),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_46),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_40),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_101),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_66),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_135),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_16),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_174),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_122),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_115),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_143),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_52),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_105),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_130),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_57),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_83),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_75),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_107),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_22),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_181),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_76),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_98),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_2),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_20),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_36),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_74),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_144),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_146),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_173),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_148),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_150),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_137),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_7),
.Y(n_275)
);

INVxp67_ASAP7_75t_SL g276 ( 
.A(n_36),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_175),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_172),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_20),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_32),
.B(n_9),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_30),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_32),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_44),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_138),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_4),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_95),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_180),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_51),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_48),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_30),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_165),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_160),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_49),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_178),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_124),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_126),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_103),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_134),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_125),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_27),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_164),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_4),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_63),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_132),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_8),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_303),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_239),
.B(n_0),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_299),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_273),
.B(n_1),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

NAND2xp33_ASAP7_75t_L g311 ( 
.A(n_215),
.B(n_42),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_184),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_303),
.Y(n_313)
);

AND2x4_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_2),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_190),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_239),
.B(n_3),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_199),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_185),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_211),
.Y(n_319)
);

AND2x6_ASAP7_75t_L g320 ( 
.A(n_229),
.B(n_43),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_191),
.Y(n_321)
);

OA21x2_ASAP7_75t_L g322 ( 
.A1(n_199),
.A2(n_93),
.B(n_177),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_294),
.B(n_3),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_294),
.B(n_5),
.Y(n_324)
);

OA22x2_ASAP7_75t_SL g325 ( 
.A1(n_235),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_204),
.Y(n_326)
);

AND2x4_ASAP7_75t_L g327 ( 
.A(n_229),
.B(n_10),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_224),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_252),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_252),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_209),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_228),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_204),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_235),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_233),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_215),
.Y(n_336)
);

BUFx8_ASAP7_75t_L g337 ( 
.A(n_256),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_211),
.B(n_15),
.Y(n_338)
);

AND2x4_ASAP7_75t_SL g339 ( 
.A(n_219),
.B(n_53),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_230),
.B(n_15),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_256),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_257),
.B(n_17),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_185),
.B(n_18),
.Y(n_343)
);

BUFx8_ASAP7_75t_L g344 ( 
.A(n_257),
.Y(n_344)
);

BUFx8_ASAP7_75t_L g345 ( 
.A(n_259),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_234),
.B(n_19),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_230),
.B(n_21),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_204),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_236),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_267),
.B(n_23),
.Y(n_350)
);

AND2x4_ASAP7_75t_L g351 ( 
.A(n_234),
.B(n_23),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_267),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_259),
.Y(n_353)
);

OAI21x1_ASAP7_75t_L g354 ( 
.A1(n_296),
.A2(n_108),
.B(n_176),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_296),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_215),
.Y(n_356)
);

AND2x6_ASAP7_75t_L g357 ( 
.A(n_237),
.B(n_54),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_290),
.B(n_24),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_219),
.Y(n_359)
);

AND2x4_ASAP7_75t_L g360 ( 
.A(n_237),
.B(n_24),
.Y(n_360)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_263),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_232),
.B(n_58),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_249),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_261),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_215),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_204),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_279),
.Y(n_367)
);

INVx6_ASAP7_75t_L g368 ( 
.A(n_263),
.Y(n_368)
);

INVx5_ASAP7_75t_L g369 ( 
.A(n_268),
.Y(n_369)
);

OA21x2_ASAP7_75t_L g370 ( 
.A1(n_189),
.A2(n_109),
.B(n_171),
.Y(n_370)
);

NAND2x1_ASAP7_75t_L g371 ( 
.A(n_281),
.B(n_25),
.Y(n_371)
);

CKINVDCx6p67_ASAP7_75t_R g372 ( 
.A(n_268),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_290),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_282),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_285),
.B(n_25),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_192),
.Y(n_376)
);

OAI22x1_ASAP7_75t_L g377 ( 
.A1(n_241),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_302),
.Y(n_378)
);

AND2x6_ASAP7_75t_L g379 ( 
.A(n_193),
.B(n_59),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_226),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_206),
.B(n_26),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_196),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_232),
.B(n_28),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_197),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_200),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_272),
.B(n_274),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_314),
.A2(n_280),
.B1(n_277),
.B2(n_201),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_320),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_326),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_308),
.B(n_272),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_314),
.A2(n_254),
.B1(n_244),
.B2(n_202),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_339),
.A2(n_334),
.B1(n_358),
.B2(n_318),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_314),
.Y(n_393)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_320),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_324),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_324),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_327),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_306),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_327),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_327),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_346),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_313),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_313),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_346),
.Y(n_404)
);

AND2x6_ASAP7_75t_L g405 ( 
.A(n_346),
.B(n_213),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g406 ( 
.A(n_337),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_320),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_373),
.B(n_274),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_320),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_326),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_333),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_351),
.B(n_360),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_333),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_351),
.Y(n_414)
);

OR2x6_ASAP7_75t_L g415 ( 
.A(n_371),
.B(n_240),
.Y(n_415)
);

INVx8_ASAP7_75t_L g416 ( 
.A(n_319),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_351),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_360),
.Y(n_418)
);

BUFx4f_ASAP7_75t_L g419 ( 
.A(n_372),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_360),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_333),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_352),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_333),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_385),
.B(n_298),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_317),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_329),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_361),
.B(n_283),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_376),
.B(n_283),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_348),
.Y(n_429)
);

INVx5_ASAP7_75t_L g430 ( 
.A(n_357),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_329),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_307),
.B(n_284),
.Y(n_432)
);

AOI22x1_ASAP7_75t_L g433 ( 
.A1(n_382),
.A2(n_286),
.B1(n_216),
.B2(n_222),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_330),
.Y(n_434)
);

INVxp33_ASAP7_75t_L g435 ( 
.A(n_386),
.Y(n_435)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_357),
.Y(n_436)
);

NOR2x1p5_ASAP7_75t_L g437 ( 
.A(n_359),
.B(n_276),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_348),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_357),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_330),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_357),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_348),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_361),
.B(n_289),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_319),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_372),
.B(n_289),
.Y(n_445)
);

AND2x2_ASAP7_75t_SL g446 ( 
.A(n_339),
.B(n_223),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_382),
.B(n_225),
.Y(n_447)
);

BUFx8_ASAP7_75t_SL g448 ( 
.A(n_359),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_337),
.B(n_291),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_366),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_366),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_337),
.B(n_291),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_384),
.B(n_231),
.Y(n_453)
);

BUFx4f_ASAP7_75t_L g454 ( 
.A(n_338),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_341),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_341),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_344),
.B(n_243),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_353),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_312),
.B(n_248),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_366),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_344),
.B(n_250),
.Y(n_461)
);

NAND3xp33_ASAP7_75t_L g462 ( 
.A(n_316),
.B(n_300),
.C(n_265),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_353),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_355),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_366),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_355),
.Y(n_466)
);

NOR3xp33_ASAP7_75t_SL g467 ( 
.A(n_380),
.B(n_255),
.C(n_251),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_315),
.B(n_264),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_345),
.B(n_183),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_336),
.Y(n_470)
);

OAI22xp33_ASAP7_75t_L g471 ( 
.A1(n_331),
.A2(n_240),
.B1(n_266),
.B2(n_305),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_336),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_321),
.Y(n_473)
);

INVx3_ASAP7_75t_R g474 ( 
.A(n_375),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_368),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_336),
.Y(n_476)
);

BUFx10_ASAP7_75t_L g477 ( 
.A(n_328),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_345),
.B(n_269),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_332),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_335),
.B(n_270),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_349),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_356),
.Y(n_482)
);

INVx5_ASAP7_75t_L g483 ( 
.A(n_357),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_368),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_363),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_364),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_345),
.B(n_271),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_367),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_379),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_374),
.B(n_186),
.Y(n_490)
);

OR2x6_ASAP7_75t_L g491 ( 
.A(n_358),
.B(n_266),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_380),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_379),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_379),
.Y(n_494)
);

NAND2xp33_ASAP7_75t_L g495 ( 
.A(n_379),
.B(n_187),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_377),
.B(n_226),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_378),
.B(n_194),
.Y(n_497)
);

AND2x6_ASAP7_75t_L g498 ( 
.A(n_340),
.B(n_278),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_340),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_347),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_383),
.B(n_205),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_422),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_477),
.B(n_432),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_394),
.B(n_347),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_428),
.B(n_381),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_455),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_495),
.A2(n_412),
.B(n_457),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_395),
.A2(n_396),
.B1(n_405),
.B2(n_412),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_499),
.B(n_309),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_419),
.Y(n_510)
);

A2O1A1Ixp33_ASAP7_75t_SL g511 ( 
.A1(n_459),
.A2(n_311),
.B(n_301),
.C(n_287),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_416),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_454),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_393),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_495),
.A2(n_354),
.B(n_311),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_501),
.B(n_343),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_390),
.B(n_473),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_498),
.A2(n_323),
.B1(n_350),
.B2(n_304),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_387),
.A2(n_304),
.B1(n_247),
.B2(n_292),
.Y(n_519)
);

NAND2xp33_ASAP7_75t_L g520 ( 
.A(n_405),
.B(n_207),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_392),
.A2(n_377),
.B1(n_247),
.B2(n_292),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_498),
.A2(n_342),
.B1(n_362),
.B2(n_188),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_454),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_500),
.B(n_208),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_479),
.B(n_368),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_393),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_394),
.B(n_288),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_412),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_408),
.B(n_245),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_481),
.B(n_310),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_406),
.B(n_210),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_498),
.A2(n_342),
.B1(n_195),
.B2(n_293),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_462),
.B(n_203),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_485),
.B(n_212),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_398),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_455),
.Y(n_536)
);

O2A1O1Ixp33_ASAP7_75t_L g537 ( 
.A1(n_486),
.A2(n_297),
.B(n_198),
.C(n_227),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_458),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_405),
.A2(n_322),
.B1(n_370),
.B2(n_365),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_488),
.B(n_214),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_388),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_490),
.B(n_217),
.Y(n_542)
);

CKINVDCx11_ASAP7_75t_R g543 ( 
.A(n_491),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_458),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_497),
.B(n_218),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_437),
.B(n_369),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_492),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_491),
.B(n_369),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_498),
.A2(n_260),
.B1(n_238),
.B2(n_242),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_409),
.B(n_369),
.Y(n_550)
);

BUFx8_ASAP7_75t_L g551 ( 
.A(n_498),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_402),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_424),
.B(n_221),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_403),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_446),
.A2(n_295),
.B1(n_258),
.B2(n_262),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_424),
.B(n_246),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_391),
.B(n_253),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_391),
.B(n_322),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_436),
.B(n_220),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_449),
.B(n_322),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_475),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_425),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_452),
.B(n_356),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_405),
.A2(n_420),
.B1(n_418),
.B2(n_417),
.Y(n_564)
);

AND2x6_ASAP7_75t_SL g565 ( 
.A(n_491),
.B(n_325),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_427),
.B(n_356),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_426),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_415),
.B(n_29),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_461),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_443),
.B(n_370),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_431),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_397),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_387),
.B(n_370),
.Y(n_573)
);

A2O1A1Ixp33_ASAP7_75t_L g574 ( 
.A1(n_404),
.A2(n_29),
.B(n_31),
.C(n_35),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_445),
.B(n_35),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_475),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_434),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_416),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_469),
.B(n_38),
.Y(n_579)
);

OR2x6_ASAP7_75t_L g580 ( 
.A(n_416),
.B(n_39),
.Y(n_580)
);

OR2x6_ASAP7_75t_L g581 ( 
.A(n_415),
.B(n_40),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_446),
.A2(n_41),
.B1(n_62),
.B2(n_64),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_478),
.B(n_65),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_440),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_456),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_463),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_494),
.B(n_67),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_464),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_444),
.B(n_41),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_496),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_466),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_414),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_397),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_399),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_399),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_400),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_478),
.B(n_73),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_400),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_401),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_447),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_487),
.B(n_77),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_484),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_484),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_470),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_514),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_516),
.B(n_487),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_502),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_516),
.B(n_459),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_560),
.A2(n_494),
.B(n_483),
.Y(n_609)
);

A2O1A1Ixp33_ASAP7_75t_L g610 ( 
.A1(n_507),
.A2(n_468),
.B(n_480),
.C(n_435),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_503),
.B(n_474),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_526),
.Y(n_612)
);

A2O1A1Ixp33_ASAP7_75t_L g613 ( 
.A1(n_507),
.A2(n_468),
.B(n_480),
.C(n_435),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_555),
.B(n_444),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_527),
.A2(n_483),
.B(n_430),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_529),
.B(n_492),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_508),
.A2(n_467),
.B1(n_415),
.B2(n_433),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_580),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_572),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_578),
.B(n_407),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_519),
.A2(n_471),
.B1(n_453),
.B2(n_439),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_592),
.B(n_489),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_592),
.B(n_489),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_517),
.B(n_493),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_573),
.A2(n_441),
.B(n_493),
.Y(n_625)
);

NOR2xp67_ASAP7_75t_SL g626 ( 
.A(n_578),
.B(n_448),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_580),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_528),
.B(n_471),
.Y(n_628)
);

O2A1O1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_537),
.A2(n_482),
.B(n_476),
.C(n_472),
.Y(n_629)
);

NOR3xp33_ASAP7_75t_L g630 ( 
.A(n_521),
.B(n_547),
.C(n_543),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_505),
.B(n_524),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_509),
.B(n_482),
.Y(n_632)
);

O2A1O1Ixp33_ASAP7_75t_L g633 ( 
.A1(n_537),
.A2(n_476),
.B(n_472),
.C(n_470),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_580),
.Y(n_634)
);

A2O1A1Ixp33_ASAP7_75t_L g635 ( 
.A1(n_558),
.A2(n_465),
.B(n_460),
.C(n_451),
.Y(n_635)
);

O2A1O1Ixp33_ASAP7_75t_SL g636 ( 
.A1(n_511),
.A2(n_587),
.B(n_601),
.C(n_559),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_564),
.B(n_389),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_572),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_513),
.B(n_80),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_SL g640 ( 
.A1(n_581),
.A2(n_451),
.B1(n_450),
.B2(n_442),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_593),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_581),
.B(n_82),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_550),
.A2(n_438),
.B(n_429),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_564),
.B(n_389),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_581),
.A2(n_569),
.B1(n_551),
.B2(n_568),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_594),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_541),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_504),
.A2(n_423),
.B(n_421),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_598),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_523),
.B(n_89),
.Y(n_650)
);

O2A1O1Ixp33_ASAP7_75t_L g651 ( 
.A1(n_574),
.A2(n_413),
.B(n_411),
.C(n_410),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_510),
.B(n_90),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_546),
.B(n_91),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_551),
.B(n_92),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_546),
.B(n_94),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_518),
.A2(n_97),
.B1(n_100),
.B2(n_102),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_548),
.B(n_104),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_595),
.Y(n_658)
);

BUFx12f_ASAP7_75t_L g659 ( 
.A(n_565),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_582),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_530),
.B(n_118),
.Y(n_661)
);

NOR3xp33_ASAP7_75t_L g662 ( 
.A(n_590),
.B(n_123),
.C(n_128),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_566),
.A2(n_129),
.B(n_131),
.Y(n_663)
);

O2A1O1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_557),
.A2(n_182),
.B(n_141),
.C(n_142),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_596),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_589),
.B(n_170),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_553),
.B(n_556),
.Y(n_667)
);

OR2x6_ASAP7_75t_SL g668 ( 
.A(n_579),
.B(n_151),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_522),
.A2(n_154),
.B1(n_156),
.B2(n_157),
.Y(n_669)
);

BUFx12f_ASAP7_75t_L g670 ( 
.A(n_533),
.Y(n_670)
);

OR2x6_ASAP7_75t_SL g671 ( 
.A(n_575),
.B(n_159),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_539),
.A2(n_563),
.B(n_534),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_531),
.B(n_166),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_562),
.B(n_169),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_540),
.A2(n_599),
.B(n_542),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_535),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_545),
.B(n_576),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_SL g678 ( 
.A1(n_532),
.A2(n_597),
.B1(n_583),
.B2(n_549),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_520),
.A2(n_600),
.B(n_584),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_567),
.A2(n_586),
.B1(n_591),
.B2(n_554),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_597),
.B(n_533),
.Y(n_681)
);

NOR2x1_ASAP7_75t_L g682 ( 
.A(n_561),
.B(n_538),
.Y(n_682)
);

BUFx12f_ASAP7_75t_L g683 ( 
.A(n_602),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_607),
.Y(n_684)
);

AO221x1_ASAP7_75t_L g685 ( 
.A1(n_618),
.A2(n_538),
.B1(n_552),
.B2(n_585),
.C(n_571),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_647),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_627),
.B(n_603),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_676),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_631),
.B(n_577),
.Y(n_689)
);

INVx6_ASAP7_75t_L g690 ( 
.A(n_683),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_636),
.A2(n_588),
.B(n_525),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_616),
.B(n_506),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_614),
.B(n_536),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_608),
.B(n_544),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_634),
.B(n_657),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_659),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_632),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_L g698 ( 
.A1(n_672),
.A2(n_604),
.B(n_606),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_628),
.B(n_645),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_667),
.B(n_656),
.C(n_669),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_620),
.B(n_611),
.Y(n_701)
);

A2O1A1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_675),
.A2(n_651),
.B(n_679),
.C(n_633),
.Y(n_702)
);

BUFx12f_ASAP7_75t_L g703 ( 
.A(n_670),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_621),
.B(n_680),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_680),
.B(n_617),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_609),
.A2(n_625),
.B(n_624),
.Y(n_706)
);

AOI221xp5_ASAP7_75t_SL g707 ( 
.A1(n_617),
.A2(n_629),
.B1(n_681),
.B2(n_678),
.C(n_640),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_625),
.A2(n_622),
.B(n_623),
.Y(n_708)
);

OR2x6_ASAP7_75t_L g709 ( 
.A(n_642),
.B(n_626),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_677),
.B(n_605),
.Y(n_710)
);

BUFx10_ASAP7_75t_L g711 ( 
.A(n_653),
.Y(n_711)
);

NAND2x1p5_ASAP7_75t_L g712 ( 
.A(n_620),
.B(n_638),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_615),
.A2(n_644),
.B(n_637),
.Y(n_713)
);

O2A1O1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_660),
.A2(n_630),
.B(n_669),
.C(n_662),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_657),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_671),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_654),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_661),
.A2(n_648),
.B(n_674),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_612),
.B(n_665),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_641),
.Y(n_720)
);

NAND3x1_ASAP7_75t_L g721 ( 
.A(n_682),
.B(n_668),
.C(n_655),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_658),
.B(n_649),
.Y(n_722)
);

BUFx4f_ASAP7_75t_L g723 ( 
.A(n_652),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_646),
.B(n_666),
.Y(n_724)
);

A2O1A1Ixp33_ASAP7_75t_L g725 ( 
.A1(n_673),
.A2(n_664),
.B(n_650),
.C(n_639),
.Y(n_725)
);

A2O1A1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_663),
.A2(n_619),
.B(n_638),
.C(n_643),
.Y(n_726)
);

O2A1O1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_647),
.A2(n_613),
.B(n_610),
.C(n_617),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_647),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_636),
.A2(n_560),
.B(n_570),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_621),
.A2(n_454),
.B1(n_508),
.B2(n_518),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_616),
.A2(n_519),
.B1(n_502),
.B2(n_380),
.Y(n_731)
);

BUFx2_ASAP7_75t_L g732 ( 
.A(n_607),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_607),
.B(n_512),
.Y(n_733)
);

NAND3xp33_ASAP7_75t_L g734 ( 
.A(n_667),
.B(n_467),
.C(n_616),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_607),
.B(n_502),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_647),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_616),
.B(n_502),
.Y(n_737)
);

BUFx12f_ASAP7_75t_L g738 ( 
.A(n_659),
.Y(n_738)
);

INVx1_ASAP7_75t_SL g739 ( 
.A(n_607),
.Y(n_739)
);

CKINVDCx11_ASAP7_75t_R g740 ( 
.A(n_659),
.Y(n_740)
);

AO31x2_ASAP7_75t_L g741 ( 
.A1(n_635),
.A2(n_515),
.A3(n_573),
.B(n_672),
.Y(n_741)
);

BUFx12f_ASAP7_75t_L g742 ( 
.A(n_659),
.Y(n_742)
);

O2A1O1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_610),
.A2(n_613),
.B(n_617),
.C(n_608),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_616),
.A2(n_519),
.B1(n_502),
.B2(n_380),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_607),
.B(n_512),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_607),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_616),
.A2(n_519),
.B1(n_502),
.B2(n_380),
.Y(n_747)
);

AO31x2_ASAP7_75t_L g748 ( 
.A1(n_635),
.A2(n_515),
.A3(n_573),
.B(n_672),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_607),
.B(n_502),
.Y(n_749)
);

NOR2x1_ASAP7_75t_L g750 ( 
.A(n_642),
.B(n_512),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_607),
.B(n_512),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_676),
.Y(n_752)
);

OAI22x1_ASAP7_75t_L g753 ( 
.A1(n_618),
.A2(n_359),
.B1(n_380),
.B2(n_496),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_616),
.B(n_502),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_607),
.B(n_512),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_631),
.B(n_502),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_636),
.A2(n_560),
.B(n_570),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_636),
.A2(n_560),
.B(n_570),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_631),
.B(n_502),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_636),
.A2(n_560),
.B(n_570),
.Y(n_760)
);

BUFx12f_ASAP7_75t_L g761 ( 
.A(n_659),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_607),
.B(n_502),
.Y(n_762)
);

AO31x2_ASAP7_75t_L g763 ( 
.A1(n_635),
.A2(n_515),
.A3(n_573),
.B(n_672),
.Y(n_763)
);

AO31x2_ASAP7_75t_L g764 ( 
.A1(n_635),
.A2(n_515),
.A3(n_573),
.B(n_672),
.Y(n_764)
);

NAND2x1p5_ASAP7_75t_L g765 ( 
.A(n_626),
.B(n_512),
.Y(n_765)
);

OAI21xp5_ASAP7_75t_L g766 ( 
.A1(n_672),
.A2(n_573),
.B(n_558),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_616),
.B(n_502),
.Y(n_767)
);

OAI22x1_ASAP7_75t_L g768 ( 
.A1(n_618),
.A2(n_359),
.B1(n_380),
.B2(n_496),
.Y(n_768)
);

AO32x2_ASAP7_75t_L g769 ( 
.A1(n_640),
.A2(n_660),
.A3(n_617),
.B1(n_669),
.B2(n_680),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_636),
.A2(n_560),
.B(n_570),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_636),
.A2(n_560),
.B(n_570),
.Y(n_771)
);

OAI22x1_ASAP7_75t_L g772 ( 
.A1(n_618),
.A2(n_359),
.B1(n_380),
.B2(n_496),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_676),
.Y(n_773)
);

INVxp33_ASAP7_75t_L g774 ( 
.A(n_737),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_756),
.B(n_759),
.Y(n_775)
);

AO21x1_ASAP7_75t_L g776 ( 
.A1(n_714),
.A2(n_705),
.B(n_743),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_741),
.Y(n_777)
);

AO31x2_ASAP7_75t_L g778 ( 
.A1(n_702),
.A2(n_729),
.A3(n_771),
.B(n_770),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_723),
.A2(n_715),
.B1(n_704),
.B2(n_767),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_695),
.B(n_733),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_697),
.B(n_754),
.Y(n_781)
);

AO31x2_ASAP7_75t_L g782 ( 
.A1(n_757),
.A2(n_760),
.A3(n_758),
.B(n_706),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_699),
.A2(n_734),
.B1(n_730),
.B2(n_716),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_688),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_749),
.B(n_762),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_741),
.Y(n_786)
);

OA21x2_ASAP7_75t_L g787 ( 
.A1(n_766),
.A2(n_707),
.B(n_698),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_740),
.Y(n_788)
);

AO21x2_ASAP7_75t_L g789 ( 
.A1(n_691),
.A2(n_727),
.B(n_713),
.Y(n_789)
);

AO31x2_ASAP7_75t_L g790 ( 
.A1(n_708),
.A2(n_726),
.A3(n_718),
.B(n_725),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_752),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_700),
.A2(n_685),
.B1(n_693),
.B2(n_709),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_773),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_689),
.B(n_719),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_720),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_739),
.B(n_710),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_765),
.B(n_709),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_686),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_684),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_694),
.B(n_744),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_724),
.A2(n_722),
.B(n_701),
.Y(n_801)
);

AO21x2_ASAP7_75t_L g802 ( 
.A1(n_748),
.A2(n_764),
.B(n_763),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_731),
.B(n_747),
.Y(n_803)
);

CKINVDCx11_ASAP7_75t_R g804 ( 
.A(n_738),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_746),
.Y(n_805)
);

AO21x2_ASAP7_75t_L g806 ( 
.A1(n_748),
.A2(n_764),
.B(n_763),
.Y(n_806)
);

OAI21x1_ASAP7_75t_L g807 ( 
.A1(n_712),
.A2(n_721),
.B(n_750),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_L g808 ( 
.A1(n_692),
.A2(n_735),
.B(n_728),
.Y(n_808)
);

AO31x2_ASAP7_75t_L g809 ( 
.A1(n_748),
.A2(n_764),
.A3(n_763),
.B(n_769),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_732),
.Y(n_810)
);

AO21x2_ASAP7_75t_L g811 ( 
.A1(n_769),
.A2(n_687),
.B(n_686),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_L g812 ( 
.A1(n_687),
.A2(n_745),
.B(n_755),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_751),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_R g814 ( 
.A1(n_717),
.A2(n_742),
.B(n_761),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_753),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_711),
.B(n_768),
.Y(n_816)
);

OA21x2_ASAP7_75t_L g817 ( 
.A1(n_769),
.A2(n_736),
.B(n_772),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_696),
.A2(n_736),
.B(n_690),
.Y(n_818)
);

BUFx2_ASAP7_75t_L g819 ( 
.A(n_690),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_703),
.B(n_502),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_756),
.B(n_631),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_688),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_712),
.Y(n_823)
);

BUFx2_ASAP7_75t_R g824 ( 
.A(n_716),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_688),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_715),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_688),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_715),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_695),
.B(n_733),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_737),
.B(n_502),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_712),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_756),
.B(n_631),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_688),
.Y(n_833)
);

NAND2x1p5_ASAP7_75t_L g834 ( 
.A(n_723),
.B(n_512),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_686),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_688),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_777),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_776),
.B(n_784),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_774),
.B(n_820),
.Y(n_839)
);

INVx4_ASAP7_75t_SL g840 ( 
.A(n_797),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_791),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_793),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_822),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_825),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_L g845 ( 
.A1(n_774),
.A2(n_803),
.B(n_801),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_827),
.B(n_833),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_785),
.B(n_794),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_830),
.B(n_821),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_836),
.B(n_795),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_786),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_783),
.B(n_780),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_810),
.Y(n_852)
);

AO21x1_ASAP7_75t_SL g853 ( 
.A1(n_792),
.A2(n_812),
.B(n_783),
.Y(n_853)
);

OR2x2_ASAP7_75t_L g854 ( 
.A(n_775),
.B(n_796),
.Y(n_854)
);

OR2x2_ASAP7_75t_SL g855 ( 
.A(n_817),
.B(n_810),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_809),
.B(n_781),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_809),
.B(n_800),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_809),
.B(n_811),
.Y(n_858)
);

INVx5_ASAP7_75t_L g859 ( 
.A(n_798),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_832),
.B(n_815),
.Y(n_860)
);

NOR2xp67_ASAP7_75t_L g861 ( 
.A(n_792),
.B(n_815),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_809),
.B(n_806),
.Y(n_862)
);

BUFx4f_ASAP7_75t_SL g863 ( 
.A(n_819),
.Y(n_863)
);

INVx4_ASAP7_75t_L g864 ( 
.A(n_835),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_829),
.B(n_802),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_799),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_797),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_779),
.B(n_787),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_787),
.B(n_817),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_817),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_782),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_778),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_805),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_865),
.B(n_789),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_856),
.B(n_826),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_864),
.Y(n_876)
);

OR2x2_ASAP7_75t_SL g877 ( 
.A(n_856),
.B(n_814),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_850),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_837),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_838),
.B(n_789),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_860),
.A2(n_797),
.B1(n_813),
.B2(n_816),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_872),
.B(n_869),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_859),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_857),
.B(n_828),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_869),
.B(n_778),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_838),
.B(n_790),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_857),
.B(n_846),
.Y(n_887)
);

OR2x2_ASAP7_75t_L g888 ( 
.A(n_854),
.B(n_826),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_846),
.B(n_790),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_849),
.B(n_790),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_849),
.B(n_778),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_864),
.Y(n_892)
);

OR2x2_ASAP7_75t_L g893 ( 
.A(n_854),
.B(n_828),
.Y(n_893)
);

INVx5_ASAP7_75t_L g894 ( 
.A(n_864),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_874),
.B(n_870),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_879),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_878),
.Y(n_897)
);

INVx5_ASAP7_75t_L g898 ( 
.A(n_894),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_887),
.B(n_862),
.Y(n_899)
);

NOR2x1p5_ASAP7_75t_L g900 ( 
.A(n_876),
.B(n_868),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_874),
.B(n_870),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_887),
.B(n_862),
.Y(n_902)
);

OR2x2_ASAP7_75t_SL g903 ( 
.A(n_875),
.B(n_868),
.Y(n_903)
);

INVx5_ASAP7_75t_L g904 ( 
.A(n_894),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_874),
.B(n_871),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_888),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_891),
.B(n_889),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_890),
.B(n_858),
.Y(n_908)
);

OR2x2_ASAP7_75t_L g909 ( 
.A(n_875),
.B(n_855),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_893),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_907),
.B(n_885),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_907),
.B(n_885),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_908),
.B(n_885),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_897),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_896),
.Y(n_915)
);

INVxp67_ASAP7_75t_SL g916 ( 
.A(n_896),
.Y(n_916)
);

OR2x2_ASAP7_75t_L g917 ( 
.A(n_899),
.B(n_880),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_906),
.A2(n_881),
.B1(n_851),
.B2(n_861),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_908),
.B(n_882),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_899),
.B(n_880),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_910),
.B(n_886),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_905),
.B(n_882),
.Y(n_922)
);

OR2x6_ASAP7_75t_L g923 ( 
.A(n_900),
.B(n_892),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_902),
.B(n_884),
.Y(n_924)
);

NOR2x1_ASAP7_75t_L g925 ( 
.A(n_923),
.B(n_883),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_919),
.B(n_902),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_924),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_919),
.B(n_895),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_916),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_923),
.A2(n_904),
.B(n_898),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_911),
.B(n_895),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_917),
.B(n_920),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_915),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_911),
.B(n_901),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_924),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_917),
.B(n_901),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_914),
.Y(n_937)
);

NAND2x1p5_ASAP7_75t_L g938 ( 
.A(n_923),
.B(n_898),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_929),
.A2(n_866),
.B(n_839),
.C(n_873),
.Y(n_939)
);

NAND2x1p5_ASAP7_75t_L g940 ( 
.A(n_925),
.B(n_898),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_928),
.B(n_912),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_931),
.B(n_922),
.Y(n_942)
);

OAI221xp5_ASAP7_75t_L g943 ( 
.A1(n_938),
.A2(n_918),
.B1(n_881),
.B2(n_861),
.C(n_923),
.Y(n_943)
);

OAI22xp33_ASAP7_75t_L g944 ( 
.A1(n_938),
.A2(n_904),
.B1(n_898),
.B2(n_909),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_SL g945 ( 
.A1(n_930),
.A2(n_898),
.B1(n_904),
.B2(n_912),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_929),
.A2(n_904),
.B(n_898),
.Y(n_946)
);

OAI21xp33_ASAP7_75t_L g947 ( 
.A1(n_927),
.A2(n_921),
.B(n_909),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_935),
.A2(n_845),
.B(n_852),
.C(n_847),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_933),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_926),
.A2(n_904),
.B(n_807),
.Y(n_950)
);

OAI221xp5_ASAP7_75t_L g951 ( 
.A1(n_945),
.A2(n_932),
.B1(n_936),
.B2(n_937),
.C(n_920),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_939),
.A2(n_928),
.B(n_931),
.C(n_934),
.Y(n_952)
);

AOI21xp33_ASAP7_75t_L g953 ( 
.A1(n_948),
.A2(n_893),
.B(n_867),
.Y(n_953)
);

O2A1O1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_943),
.A2(n_867),
.B(n_847),
.C(n_848),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_947),
.B(n_934),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_940),
.A2(n_903),
.B1(n_877),
.B2(n_904),
.Y(n_956)
);

AOI221xp5_ASAP7_75t_SL g957 ( 
.A1(n_951),
.A2(n_947),
.B1(n_944),
.B2(n_950),
.C(n_877),
.Y(n_957)
);

NOR3xp33_ASAP7_75t_L g958 ( 
.A(n_954),
.B(n_804),
.C(n_788),
.Y(n_958)
);

NAND3xp33_ASAP7_75t_L g959 ( 
.A(n_952),
.B(n_946),
.C(n_949),
.Y(n_959)
);

OAI211xp5_ASAP7_75t_SL g960 ( 
.A1(n_958),
.A2(n_804),
.B(n_953),
.C(n_955),
.Y(n_960)
);

AOI221xp5_ASAP7_75t_L g961 ( 
.A1(n_957),
.A2(n_959),
.B1(n_956),
.B2(n_941),
.C(n_942),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_961),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_960),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_963),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_962),
.B(n_913),
.Y(n_965)
);

OR2x2_ASAP7_75t_L g966 ( 
.A(n_965),
.B(n_788),
.Y(n_966)
);

XOR2x2_ASAP7_75t_L g967 ( 
.A(n_965),
.B(n_824),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_966),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_967),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_968),
.Y(n_970)
);

AOI221xp5_ASAP7_75t_L g971 ( 
.A1(n_969),
.A2(n_964),
.B1(n_818),
.B2(n_841),
.C(n_843),
.Y(n_971)
);

XOR2xp5_ASAP7_75t_L g972 ( 
.A(n_968),
.B(n_834),
.Y(n_972)
);

XNOR2x1_ASAP7_75t_L g973 ( 
.A(n_969),
.B(n_834),
.Y(n_973)
);

XNOR2x1_ASAP7_75t_SL g974 ( 
.A(n_973),
.B(n_863),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_972),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_971),
.A2(n_808),
.B(n_831),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_970),
.A2(n_840),
.B1(n_851),
.B2(n_844),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_975),
.B(n_974),
.Y(n_978)
);

AOI21xp33_ASAP7_75t_L g979 ( 
.A1(n_977),
.A2(n_842),
.B(n_823),
.Y(n_979)
);

OR2x6_ASAP7_75t_L g980 ( 
.A(n_978),
.B(n_976),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_980),
.A2(n_979),
.B1(n_840),
.B2(n_853),
.Y(n_981)
);


endmodule