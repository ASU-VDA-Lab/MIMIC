module fake_jpeg_23281_n_233 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_233);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_37),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_0),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_18),
.B1(n_25),
.B2(n_16),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_39),
.A2(n_35),
.B1(n_31),
.B2(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_18),
.B1(n_25),
.B2(n_28),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_48),
.B(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_15),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_28),
.B1(n_21),
.B2(n_25),
.Y(n_48)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_50),
.B(n_53),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_32),
.A2(n_26),
.B1(n_23),
.B2(n_17),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_56),
.B(n_14),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_34),
.A2(n_26),
.B1(n_23),
.B2(n_16),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_23),
.B1(n_26),
.B2(n_34),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_59),
.A2(n_62),
.B1(n_72),
.B2(n_55),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_61),
.B(n_63),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_31),
.B1(n_27),
.B2(n_19),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_65),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_42),
.B(n_54),
.C(n_31),
.Y(n_92)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_71),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_69),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_56),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_36),
.B1(n_27),
.B2(n_24),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx8_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_30),
.Y(n_74)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_49),
.B(n_71),
.Y(n_80)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_49),
.C(n_41),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_93),
.C(n_74),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_58),
.A2(n_48),
.B1(n_44),
.B2(n_39),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_81),
.B1(n_92),
.B2(n_98),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_80),
.A2(n_90),
.B(n_46),
.Y(n_119)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_53),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_53),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_49),
.B(n_48),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_49),
.C(n_41),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

OA21x2_ASAP7_75t_SL g97 ( 
.A1(n_70),
.A2(n_53),
.B(n_69),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_97),
.A2(n_88),
.B1(n_84),
.B2(n_96),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_62),
.A2(n_42),
.B1(n_46),
.B2(n_43),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_102),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_109),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_79),
.A2(n_77),
.B1(n_75),
.B2(n_65),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_106),
.A2(n_111),
.B1(n_115),
.B2(n_120),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_89),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_116),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_97),
.B(n_63),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_110),
.B(n_112),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_78),
.A2(n_60),
.B1(n_67),
.B2(n_61),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_77),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_73),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_113),
.B(n_114),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_73),
.Y(n_114)
);

AOI22x1_ASAP7_75t_SL g115 ( 
.A1(n_80),
.A2(n_30),
.B1(n_54),
.B2(n_19),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_66),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_24),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_30),
.B1(n_66),
.B2(n_24),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_82),
.B1(n_83),
.B2(n_95),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_98),
.B(n_27),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_92),
.A2(n_68),
.B1(n_30),
.B2(n_27),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_22),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_87),
.Y(n_128)
);

INVxp67_ASAP7_75t_SL g122 ( 
.A(n_103),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_122),
.Y(n_153)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_136),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_130),
.B1(n_138),
.B2(n_140),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_105),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_128),
.B(n_133),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_82),
.B1(n_99),
.B2(n_94),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_134),
.B(n_135),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_94),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_107),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_24),
.B1(n_87),
.B2(n_15),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_87),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_121),
.Y(n_161)
);

AOI22x1_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_117),
.B1(n_120),
.B2(n_106),
.Y(n_142)
);

AOI322xp5_ASAP7_75t_L g145 ( 
.A1(n_142),
.A2(n_127),
.A3(n_129),
.B1(n_140),
.B2(n_116),
.C1(n_124),
.C2(n_110),
.Y(n_145)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_145),
.A2(n_22),
.B1(n_20),
.B2(n_8),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_101),
.Y(n_146)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_101),
.Y(n_148)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_119),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_109),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_160),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_115),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_155),
.B(n_157),
.Y(n_167)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_141),
.B(n_108),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

MAJx2_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_104),
.C(n_118),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_161),
.A2(n_133),
.B1(n_138),
.B2(n_126),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_142),
.B1(n_134),
.B2(n_124),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_162),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_123),
.B(n_87),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_158),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_15),
.C(n_22),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_171),
.C(n_175),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_15),
.C(n_22),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_156),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_22),
.C(n_20),
.Y(n_175)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_177),
.B(n_151),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_182),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_146),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_183),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_147),
.B1(n_144),
.B2(n_156),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_185),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_150),
.B1(n_153),
.B2(n_2),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_22),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_189),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_20),
.C(n_1),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_188),
.C(n_168),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_172),
.C(n_163),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_187),
.C(n_190),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_173),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_162),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_181),
.C(n_184),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_20),
.C(n_1),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_172),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_20),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_204),
.Y(n_217)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_163),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_203),
.A2(n_208),
.B(n_192),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_197),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_206),
.C(n_207),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_196),
.A2(n_8),
.B(n_12),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_8),
.C(n_12),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_210),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_20),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_198),
.Y(n_213)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_214),
.B(n_215),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_200),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_203),
.A2(n_191),
.B1(n_193),
.B2(n_192),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_216),
.A2(n_194),
.B1(n_191),
.B2(n_201),
.Y(n_218)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_218),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_217),
.A2(n_7),
.B1(n_11),
.B2(n_10),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_222),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_5),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_212),
.C(n_211),
.Y(n_223)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_223),
.Y(n_227)
);

AOI21x1_ASAP7_75t_L g228 ( 
.A1(n_224),
.A2(n_225),
.B(n_3),
.Y(n_228)
);

OAI321xp33_ASAP7_75t_L g225 ( 
.A1(n_220),
.A2(n_4),
.A3(n_5),
.B1(n_9),
.B2(n_10),
.C(n_12),
.Y(n_225)
);

NAND3xp33_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_10),
.C(n_4),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_219),
.B(n_226),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_218),
.C(n_227),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_9),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_5),
.C(n_3),
.Y(n_233)
);


endmodule