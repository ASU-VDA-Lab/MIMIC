module real_aes_6714_n_10 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_1, n_10);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_1;
output n_10;
wire n_17;
wire n_28;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_27;
wire n_23;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
NOR2xp33_ASAP7_75t_L g20 ( .A(n_0), .B(n_6), .Y(n_20) );
AOI322xp5_ASAP7_75t_L g10 ( .A1(n_1), .A2(n_2), .A3(n_8), .B1(n_11), .B2(n_25), .C1(n_29), .C2(n_30), .Y(n_10) );
CKINVDCx20_ASAP7_75t_R g24 ( .A(n_3), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_4), .B(n_23), .Y(n_22) );
INVx1_ASAP7_75t_L g19 ( .A(n_5), .Y(n_19) );
INVx1_ASAP7_75t_L g23 ( .A(n_7), .Y(n_23) );
INVx2_ASAP7_75t_L g16 ( .A(n_9), .Y(n_16) );
OR2x2_ASAP7_75t_L g28 ( .A(n_9), .B(n_17), .Y(n_28) );
INVx1_ASAP7_75t_SL g11 ( .A(n_12), .Y(n_11) );
HB1xp67_ASAP7_75t_L g29 ( .A(n_12), .Y(n_29) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_13), .Y(n_12) );
INVx1_ASAP7_75t_SL g32 ( .A(n_13), .Y(n_32) );
NAND2xp5_ASAP7_75t_SL g13 ( .A(n_14), .B(n_21), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_15), .Y(n_14) );
NOR2x2_ASAP7_75t_L g15 ( .A(n_16), .B(n_17), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g31 ( .A(n_17), .B(n_32), .Y(n_31) );
INVx2_ASAP7_75t_L g17 ( .A(n_18), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_19), .B(n_20), .Y(n_18) );
NOR2xp33_ASAP7_75t_SL g21 ( .A(n_22), .B(n_24), .Y(n_21) );
INVx1_ASAP7_75t_SL g25 ( .A(n_26), .Y(n_25) );
BUFx2_ASAP7_75t_L g26 ( .A(n_27), .Y(n_26) );
BUFx2_ASAP7_75t_L g27 ( .A(n_28), .Y(n_27) );
INVx1_ASAP7_75t_SL g30 ( .A(n_31), .Y(n_30) );
endmodule