module fake_jpeg_2531_n_70 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_70);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_70;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_4),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_18),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_21),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_9),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_14),
.A2(n_15),
.B1(n_12),
.B2(n_17),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_24),
.Y(n_32)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_19),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_9),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_20),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_36),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_32),
.A2(n_17),
.B1(n_13),
.B2(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_40),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_13),
.C(n_11),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_10),
.B(n_17),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_41),
.Y(n_46)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_20),
.B1(n_11),
.B2(n_10),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_30),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_39),
.B1(n_31),
.B2(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_30),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_36),
.B(n_35),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_37),
.B1(n_34),
.B2(n_40),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_55),
.B1(n_0),
.B2(n_2),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_49),
.B(n_6),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_31),
.C(n_21),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_49),
.B(n_16),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_16),
.B1(n_1),
.B2(n_2),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_50),
.A2(n_46),
.B1(n_45),
.B2(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_60),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_59),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_54),
.C(n_50),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_63),
.C(n_61),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_56),
.B(n_3),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_64),
.B(n_65),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_64),
.A2(n_4),
.B1(n_8),
.B2(n_0),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_8),
.B(n_3),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_67),
.C(n_66),
.Y(n_69)
);

BUFx24_ASAP7_75t_SL g70 ( 
.A(n_69),
.Y(n_70)
);


endmodule