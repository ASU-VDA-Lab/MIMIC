module real_jpeg_300_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_1),
.A2(n_44),
.B1(n_70),
.B2(n_72),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_1),
.A2(n_36),
.B1(n_38),
.B2(n_44),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_1),
.A2(n_44),
.B1(n_59),
.B2(n_65),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_2),
.B(n_29),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_2),
.B(n_39),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_2),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_2),
.A2(n_29),
.B(n_185),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_2),
.B(n_95),
.Y(n_247)
);

AOI21xp33_ASAP7_75t_L g254 ( 
.A1(n_2),
.A2(n_38),
.B(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_2),
.B(n_59),
.C(n_75),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_2),
.A2(n_70),
.B1(n_72),
.B2(n_221),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_2),
.B(n_62),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_2),
.B(n_79),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_3),
.A2(n_41),
.B1(n_59),
.B2(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_3),
.A2(n_41),
.B1(n_70),
.B2(n_72),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_3),
.A2(n_36),
.B1(n_38),
.B2(n_41),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_6),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_6),
.A2(n_36),
.B1(n_38),
.B2(n_176),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_6),
.A2(n_70),
.B1(n_72),
.B2(n_176),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_6),
.A2(n_59),
.B1(n_65),
.B2(n_176),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_7),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_7),
.A2(n_36),
.B1(n_38),
.B2(n_195),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_7),
.A2(n_70),
.B1(n_72),
.B2(n_195),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_7),
.A2(n_59),
.B1(n_65),
.B2(n_195),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_8),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_8),
.A2(n_36),
.B1(n_38),
.B2(n_142),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_8),
.A2(n_70),
.B1(n_72),
.B2(n_142),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_8),
.A2(n_59),
.B1(n_65),
.B2(n_142),
.Y(n_249)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_10),
.A2(n_36),
.B1(n_38),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_10),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_92),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_10),
.A2(n_70),
.B1(n_72),
.B2(n_92),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_10),
.A2(n_59),
.B1(n_65),
.B2(n_92),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_13),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_13),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_13),
.A2(n_36),
.B1(n_38),
.B2(n_69),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_69),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_13),
.A2(n_59),
.B1(n_65),
.B2(n_69),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_14),
.A2(n_15),
.B1(n_21),
.B2(n_22),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_14),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_16),
.A2(n_29),
.B1(n_30),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_16),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_16),
.A2(n_36),
.B1(n_38),
.B2(n_86),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_16),
.A2(n_70),
.B1(n_72),
.B2(n_86),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_L g212 ( 
.A1(n_16),
.A2(n_59),
.B1(n_65),
.B2(n_86),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_17),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_18),
.A2(n_29),
.B1(n_30),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_18),
.A2(n_36),
.B1(n_38),
.B2(n_84),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_18),
.A2(n_70),
.B1(n_72),
.B2(n_84),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_18),
.A2(n_59),
.B1(n_65),
.B2(n_84),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_47),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_45),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_42),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_39),
.B(n_40),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_27),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_27),
.A2(n_39),
.B1(n_141),
.B2(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_27),
.A2(n_39),
.B1(n_43),
.B2(n_323),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_35),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI32xp33_ASAP7_75t_L g184 ( 
.A1(n_30),
.A2(n_34),
.A3(n_38),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_35)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_32),
.B(n_36),
.Y(n_186)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_35),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_35),
.A2(n_82),
.B1(n_85),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_35),
.A2(n_82),
.B1(n_83),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_35),
.A2(n_82),
.B1(n_105),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_35),
.A2(n_82),
.B1(n_194),
.B2(n_196),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_35),
.A2(n_82),
.B1(n_194),
.B2(n_233),
.Y(n_232)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_36),
.A2(n_38),
.B1(n_96),
.B2(n_97),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_36),
.B(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI32xp33_ASAP7_75t_L g219 ( 
.A1(n_38),
.A2(n_70),
.A3(n_96),
.B1(n_220),
.B2(n_222),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_42),
.B(n_329),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_46),
.B(n_332),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_328),
.B(n_330),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_316),
.B(n_327),
.Y(n_48)
);

AO21x1_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_156),
.B(n_313),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_143),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_116),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_52),
.B(n_116),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_87),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_53),
.B(n_102),
.C(n_114),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_80),
.B(n_81),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_54),
.A2(n_55),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_66),
.Y(n_55)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_56),
.A2(n_80),
.B1(n_81),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_56),
.A2(n_66),
.B1(n_67),
.B2(n_80),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_61),
.B(n_63),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_57),
.A2(n_61),
.B1(n_130),
.B2(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_57),
.A2(n_61),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_57),
.A2(n_61),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_58),
.A2(n_62),
.B1(n_64),
.B2(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_58),
.A2(n_62),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_58),
.A2(n_62),
.B1(n_188),
.B2(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_58),
.A2(n_62),
.B1(n_225),
.B2(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_58),
.A2(n_62),
.B1(n_221),
.B2(n_275),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_58),
.A2(n_62),
.B1(n_275),
.B2(n_279),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_59),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_65),
.B1(n_75),
.B2(n_76),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_59),
.B(n_273),
.Y(n_272)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_73),
.B1(n_78),
.B2(n_79),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_68),
.A2(n_73),
.B1(n_79),
.B2(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_70),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_72),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

AO22x2_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_72),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_70),
.B(n_263),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_72),
.B(n_97),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_78),
.B1(n_79),
.B2(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_73),
.A2(n_79),
.B(n_101),
.Y(n_108)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_73),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_73),
.A2(n_79),
.B1(n_215),
.B2(n_217),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_73),
.A2(n_79),
.B1(n_217),
.B2(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_73),
.A2(n_79),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_73),
.A2(n_79),
.B1(n_245),
.B2(n_266),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_77),
.A2(n_134),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_77),
.A2(n_169),
.B1(n_216),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_102),
.B1(n_114),
.B2(n_115),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_88),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_88),
.A2(n_89),
.B(n_100),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_100),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_93),
.B1(n_95),
.B2(n_99),
.Y(n_89)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_91),
.A2(n_94),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_95),
.B1(n_99),
.B2(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_93),
.A2(n_95),
.B1(n_137),
.B2(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_93),
.A2(n_95),
.B(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_94),
.A2(n_112),
.B1(n_138),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_94),
.A2(n_138),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_94),
.A2(n_138),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_94),
.A2(n_138),
.B1(n_191),
.B2(n_207),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_94),
.A2(n_138),
.B1(n_206),
.B2(n_254),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_96),
.Y(n_97)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_103),
.A2(n_104),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_108),
.C(n_110),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_104),
.B(n_147),
.C(n_154),
.Y(n_317)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_113),
.Y(n_107)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_108),
.A2(n_113),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_108),
.B(n_150),
.C(n_152),
.Y(n_326)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_122),
.C(n_124),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_117),
.A2(n_118),
.B1(n_122),
.B2(n_123),
.Y(n_159)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_135),
.C(n_139),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_125),
.A2(n_126),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_127),
.A2(n_128),
.B1(n_131),
.B2(n_132),
.Y(n_197)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_139),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_143),
.A2(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_155),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_144),
.B(n_155),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_154),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_151),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_153),
.Y(n_323)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_177),
.B(n_312),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_158),
.B(n_160),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_165),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_164),
.Y(n_199)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_172),
.C(n_174),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_167),
.B(n_170),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_174),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_173),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_200),
.B(n_311),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_198),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_179),
.B(n_198),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.C(n_197),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_180),
.B(n_197),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_182),
.B(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_190),
.C(n_193),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_183),
.B(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_184),
.B(n_187),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_190),
.B(n_193),
.Y(n_301)
);

AOI31xp33_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_295),
.A3(n_304),
.B(n_308),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_240),
.B(n_294),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_227),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_203),
.B(n_227),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_214),
.C(n_218),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_204),
.B(n_291),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_209),
.C(n_213),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_213),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_211),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_214),
.B(n_218),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_223),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_223),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_229),
.B(n_230),
.C(n_231),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_232),
.B(n_235),
.C(n_239),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_238),
.B2(n_239),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_236),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_289),
.B(n_293),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_258),
.B(n_288),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_250),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_243),
.B(n_250),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_247),
.C(n_248),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_247),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_246),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_268),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_249),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_251),
.B(n_253),
.C(n_256),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_269),
.B(n_287),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_267),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_267),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_264),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_281),
.B(n_286),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_276),
.B(n_280),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_278),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_279),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_285),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_285),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_292),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_299),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.C(n_303),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_303),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_306),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_318),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_326),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_322),
.B1(n_324),
.B2(n_325),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_320),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_324),
.C(n_326),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_329),
.Y(n_332)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);


endmodule