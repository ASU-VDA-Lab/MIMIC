module fake_jpeg_3062_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_22),
.B(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_34),
.B1(n_32),
.B2(n_31),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_30),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_53),
.B(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

CKINVDCx6p67_ASAP7_75t_R g58 ( 
.A(n_54),
.Y(n_58)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_65),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_36),
.B(n_35),
.C(n_45),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_45),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_66),
.B(n_63),
.Y(n_86)
);

AND2x6_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_76),
.Y(n_82)
);

BUFx24_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_72),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_65),
.A2(n_52),
.B1(n_51),
.B2(n_46),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_59),
.B1(n_39),
.B2(n_36),
.Y(n_84)
);

AO22x1_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_54),
.B1(n_44),
.B2(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_54),
.C(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_48),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_40),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_47),
.Y(n_85)
);

OAI32xp33_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_58),
.A3(n_55),
.B1(n_48),
.B2(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_83),
.Y(n_95)
);

AO22x1_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_71),
.B1(n_55),
.B2(n_67),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_85),
.B(n_90),
.Y(n_93)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_41),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_89),
.Y(n_92)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_37),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_71),
.B1(n_59),
.B2(n_68),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_104),
.B1(n_18),
.B2(n_17),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_100),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_29),
.C(n_28),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_82),
.C(n_21),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_26),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_103),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_1),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_78),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_101),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_81),
.A2(n_4),
.B(n_5),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_102),
.Y(n_108)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

NOR2x1_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_83),
.Y(n_105)
);

OAI321xp33_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_95),
.A3(n_99),
.B1(n_93),
.B2(n_102),
.C(n_94),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_11),
.C(n_12),
.Y(n_120)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_111),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_80),
.B(n_84),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_114),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_8),
.Y(n_113)
);

OA21x2_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_115),
.B(n_116),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_9),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_11),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g117 ( 
.A(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_119),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_106),
.C(n_112),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_118),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_123),
.B(n_124),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_110),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_121),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_126),
.A3(n_108),
.B1(n_111),
.B2(n_105),
.C1(n_122),
.C2(n_15),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_12),
.B(n_13),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_130),
.A2(n_13),
.B(n_14),
.C(n_16),
.Y(n_131)
);

AOI21x1_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_14),
.B(n_16),
.Y(n_132)
);


endmodule