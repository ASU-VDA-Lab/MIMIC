module real_jpeg_6881_n_30 (n_17, n_8, n_0, n_21, n_2, n_29, n_180, n_10, n_175, n_9, n_178, n_12, n_24, n_176, n_6, n_28, n_171, n_177, n_179, n_23, n_11, n_14, n_172, n_25, n_7, n_22, n_18, n_3, n_174, n_5, n_4, n_173, n_1, n_26, n_27, n_20, n_19, n_16, n_15, n_13, n_30);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_29;
input n_180;
input n_10;
input n_175;
input n_9;
input n_178;
input n_12;
input n_24;
input n_176;
input n_6;
input n_28;
input n_171;
input n_177;
input n_179;
input n_23;
input n_11;
input n_14;
input n_172;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_174;
input n_5;
input n_4;
input n_173;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_30;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_150;
wire n_41;
wire n_74;
wire n_32;
wire n_80;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_0),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_1),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_2),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_2),
.B(n_149),
.Y(n_157)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_3),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_4),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_4),
.B(n_152),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_5),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_5),
.B(n_111),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_7),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_7),
.B(n_33),
.Y(n_159)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_7),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_8),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_10),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_10),
.B(n_60),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_11),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_12),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_13),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_14),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_14),
.B(n_70),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_15),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_16),
.Y(n_136)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_17),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_18),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_19),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_19),
.B(n_55),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_20),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_20),
.B(n_135),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_21),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_21),
.B(n_73),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_22),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_23),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_23),
.B(n_125),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_24),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_24),
.B(n_95),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_25),
.B(n_50),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_26),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_27),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_27),
.B(n_44),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_28),
.B(n_86),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_29),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_160),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_39),
.B(n_159),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_35),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_35),
.B(n_150),
.Y(n_149)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_71),
.Y(n_70)
);

BUFx8_ASAP7_75t_L g113 ( 
.A(n_37),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_147),
.B(n_156),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_127),
.B(n_141),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_65),
.B(n_115),
.C(n_124),
.Y(n_41)
);

NOR4xp25_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_49),
.C(n_54),
.D(n_59),
.Y(n_42)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_43),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_49),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_52),
.B(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_52),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_52),
.Y(n_167)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_53),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_54),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21x1_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_110),
.B(n_114),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_102),
.B(n_109),
.Y(n_66)
);

AO221x1_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_77),
.B1(n_99),
.B2(n_100),
.C(n_101),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_126),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_83),
.B(n_98),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_94),
.B(n_97),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_88),
.B(n_93),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_92),
.Y(n_93)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_108),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_136),
.Y(n_135)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B(n_121),
.C(n_122),
.D(n_123),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_133),
.C(n_137),
.Y(n_127)
);

A2O1A1O1Ixp25_ASAP7_75t_L g141 ( 
.A1(n_128),
.A2(n_137),
.B(n_142),
.C(n_145),
.D(n_146),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_130),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_134),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_140),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_157),
.B(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_169),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_168),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_168),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_171),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_172),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_173),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_174),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_175),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_176),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_177),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_178),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_179),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_180),
.Y(n_112)
);


endmodule