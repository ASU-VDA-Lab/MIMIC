module fake_jpeg_20952_n_107 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_107);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_48),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_51),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_45),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_55),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_39),
.B1(n_46),
.B2(n_42),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_57),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_15),
.C(n_27),
.Y(n_57)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_66),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_47),
.B1(n_44),
.B2(n_34),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_65),
.A2(n_62),
.B1(n_59),
.B2(n_3),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_41),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_68),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_70),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_37),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_74),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_77),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_76),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_1),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_1),
.B(n_2),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_13),
.Y(n_90)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_2),
.Y(n_81)
);

AO22x1_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_82),
.B1(n_10),
.B2(n_11),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_4),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_5),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_80),
.C(n_75),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_72),
.B1(n_16),
.B2(n_19),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_90),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_94),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_14),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_96),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_97),
.B(n_91),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_99),
.C(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_101),
.B(n_98),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_85),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_83),
.C(n_21),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_20),
.Y(n_107)
);


endmodule