module real_jpeg_11449_n_16 (n_5, n_4, n_8, n_0, n_12, n_400, n_1, n_11, n_14, n_2, n_13, n_15, n_401, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_400;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_401;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_0),
.Y(n_106)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_3),
.B(n_51),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_3),
.B(n_38),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_3),
.B(n_26),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_3),
.B(n_106),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_3),
.B(n_93),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_4),
.B(n_29),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_4),
.B(n_51),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_4),
.B(n_26),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_4),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_4),
.B(n_38),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_5),
.B(n_32),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_5),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_5),
.B(n_106),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_5),
.B(n_29),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_5),
.B(n_38),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_5),
.B(n_43),
.Y(n_305)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_7),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_7),
.B(n_93),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_7),
.B(n_32),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_7),
.B(n_29),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_7),
.B(n_51),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_7),
.B(n_38),
.Y(n_292)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_8),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_8),
.B(n_43),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_8),
.B(n_93),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_8),
.B(n_32),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_8),
.B(n_26),
.Y(n_324)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_11),
.B(n_26),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_11),
.B(n_29),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_11),
.B(n_93),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_11),
.B(n_32),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_11),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_11),
.B(n_51),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_11),
.B(n_38),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_11),
.B(n_43),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_13),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_13),
.B(n_29),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_13),
.B(n_51),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_13),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_13),
.B(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_13),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_13),
.B(n_38),
.Y(n_326)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_14),
.Y(n_95)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_15),
.B(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_15),
.B(n_106),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_15),
.B(n_93),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_15),
.B(n_26),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_15),
.B(n_29),
.Y(n_344)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_118),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_117),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_77),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_21),
.B(n_77),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_62),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_46),
.C(n_53),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_23),
.B(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_33),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_24),
.B(n_35),
.C(n_39),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.C(n_31),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_25),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_25),
.B(n_55),
.C(n_60),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_25),
.A2(n_31),
.B1(n_61),
.B2(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_25),
.A2(n_61),
.B1(n_107),
.B2(n_108),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_25),
.B(n_107),
.C(n_251),
.Y(n_271)
);

INVx5_ASAP7_75t_SL g147 ( 
.A(n_26),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_28),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_28),
.A2(n_81),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_28),
.B(n_289),
.C(n_292),
.Y(n_337)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_30),
.B(n_36),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_31),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_31),
.B(n_91),
.C(n_96),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_31),
.A2(n_84),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_31),
.B(n_199),
.C(n_201),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_31),
.A2(n_84),
.B1(n_91),
.B2(n_92),
.Y(n_371)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_32),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_36),
.B(n_135),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_41),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_41),
.B(n_109),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_42),
.B(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_42),
.B(n_178),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_42),
.B(n_136),
.Y(n_328)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_46),
.A2(n_53),
.B1(n_54),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.C(n_50),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_47),
.B(n_50),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_48),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_48),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_49),
.B(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_51),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_55),
.A2(n_56),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_105),
.C(n_107),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_60),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_59),
.A2(n_60),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_60),
.B(n_96),
.C(n_263),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_76),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_71),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_65),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_87),
.C(n_88),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_65),
.A2(n_69),
.B1(n_364),
.B2(n_365),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_66),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_67),
.A2(n_68),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_68),
.B(n_302),
.C(n_304),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_112),
.C(n_113),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_78),
.B(n_393),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_97),
.C(n_101),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_79),
.B(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_85),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_86),
.C(n_90),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_87),
.B(n_88),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_89),
.B(n_133),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_103),
.C(n_110),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_91),
.A2(n_92),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_91),
.A2(n_92),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_91),
.A2(n_92),
.B1(n_110),
.B2(n_359),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_92),
.B(n_159),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_92),
.B(n_342),
.C(n_344),
.Y(n_360)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_94),
.B(n_178),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_96),
.A2(n_260),
.B1(n_261),
.B2(n_264),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_96),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_96),
.A2(n_264),
.B1(n_370),
.B2(n_371),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_97),
.A2(n_101),
.B1(n_102),
.B2(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_97),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_99),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_103),
.A2(n_104),
.B1(n_357),
.B2(n_358),
.Y(n_356)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_105),
.B(n_138),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_105),
.A2(n_140),
.B1(n_206),
.B2(n_207),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_105),
.A2(n_107),
.B1(n_108),
.B2(n_140),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_105),
.B(n_207),
.C(n_305),
.Y(n_342)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_109),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_110),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_112),
.Y(n_394)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI321xp33_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_381),
.A3(n_390),
.B1(n_395),
.B2(n_396),
.C(n_400),
.Y(n_118)
);

AOI321xp33_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_313),
.A3(n_347),
.B1(n_375),
.B2(n_380),
.C(n_401),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_254),
.C(n_308),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_225),
.B(n_253),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_193),
.B(n_224),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_162),
.B(n_192),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_141),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_125),
.B(n_141),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.C(n_137),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_144),
.B1(n_145),
.B2(n_153),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_126),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_126),
.B(n_189),
.Y(n_188)
);

FAx1_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_128),
.CI(n_129),
.CON(n_126),
.SN(n_126)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_130),
.A2(n_131),
.B1(n_137),
.B2(n_190),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_132),
.B(n_134),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_135),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_136),
.B(n_147),
.Y(n_199)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_137),
.Y(n_190)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_154),
.B2(n_161),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_144),
.B(n_153),
.C(n_161),
.Y(n_194)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_146),
.B(n_149),
.C(n_152),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_151),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_155),
.B(n_157),
.C(n_158),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_159),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_159),
.A2(n_160),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_159),
.B(n_276),
.C(n_279),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_186),
.B(n_191),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_175),
.B(n_185),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_170),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_165),
.B(n_170),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_173),
.C(n_174),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_180),
.B(n_184),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_177),
.B(n_179),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_187),
.B(n_188),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_194),
.B(n_195),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_210),
.B2(n_211),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_212),
.C(n_223),
.Y(n_226)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_203),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_204),
.C(n_205),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_208),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_222),
.B2(n_223),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_221),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_218),
.C(n_220),
.Y(n_244)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_216),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_217),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_226),
.B(n_227),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_243),
.B2(n_252),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_242),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_230),
.B(n_242),
.C(n_252),
.Y(n_309)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_238),
.B2(n_239),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_233),
.B(n_240),
.C(n_241),
.Y(n_272)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g397 ( 
.A(n_234),
.Y(n_397)
);

FAx1_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_236),
.CI(n_237),
.CON(n_234),
.SN(n_234)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_235),
.B(n_236),
.C(n_237),
.Y(n_281)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_243),
.Y(n_252)
);

BUFx24_ASAP7_75t_SL g399 ( 
.A(n_243),
.Y(n_399)
);

FAx1_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_245),
.CI(n_249),
.CON(n_243),
.SN(n_243)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_244),
.B(n_245),
.C(n_249),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B(n_248),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_247),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_248),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_280)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_248),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI21xp33_ASAP7_75t_L g376 ( 
.A1(n_255),
.A2(n_377),
.B(n_378),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_285),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_256),
.B(n_285),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_273),
.C(n_284),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_257),
.B(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_272),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_265),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_259),
.B(n_265),
.C(n_272),
.Y(n_307)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_262),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_271),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_268),
.B(n_269),
.C(n_271),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_273),
.A2(n_274),
.B1(n_284),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_280),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_281),
.C(n_283),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_278),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_281),
.Y(n_282)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_284),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_307),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_296),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_287),
.B(n_296),
.C(n_307),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_293),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_288),
.B(n_294),
.C(n_295),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_297),
.B(n_299),
.C(n_300),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_304),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_302),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_309),
.B(n_310),
.Y(n_377)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_314),
.A2(n_376),
.B(n_379),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_315),
.B(n_316),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_346),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_318),
.B(n_319),
.C(n_346),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_338),
.B2(n_339),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_320),
.B(n_340),
.C(n_341),
.Y(n_374)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_330),
.B2(n_331),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_322),
.B(n_332),
.C(n_337),
.Y(n_353)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_324),
.B(n_326),
.C(n_328),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_326),
.A2(n_327),
.B1(n_328),
.B2(n_329),
.Y(n_325)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_326),
.Y(n_329)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_332),
.A2(n_333),
.B1(n_336),
.B2(n_337),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_344),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_348),
.B(n_349),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_374),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_361),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_351),
.B(n_361),
.C(n_374),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_352),
.B(n_356),
.C(n_360),
.Y(n_389)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_360),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_363),
.B1(n_366),
.B2(n_367),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_362),
.B(n_368),
.C(n_373),
.Y(n_385)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_369),
.B1(n_372),
.B2(n_373),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_373),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_382),
.B(n_383),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_389),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_385),
.B(n_386),
.C(n_389),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_391),
.B(n_392),
.Y(n_396)
);


endmodule