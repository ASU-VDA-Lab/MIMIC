module fake_jpeg_24662_n_343 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_44),
.Y(n_57)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_0),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_30),
.B1(n_23),
.B2(n_19),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_1),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_1),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_50),
.A2(n_55),
.B1(n_48),
.B2(n_42),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_49),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_67),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_30),
.B(n_19),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_35),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_59),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_66),
.B(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_35),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_23),
.B1(n_42),
.B2(n_48),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_100),
.B1(n_96),
.B2(n_54),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_75),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_83),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_59),
.B(n_41),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_41),
.C(n_43),
.Y(n_123)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_47),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_89),
.Y(n_101)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_48),
.B1(n_42),
.B2(n_38),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_87),
.A2(n_40),
.B1(n_62),
.B2(n_30),
.Y(n_125)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_47),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_60),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_19),
.B(n_38),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_57),
.B(n_22),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_92),
.B(n_58),
.Y(n_107)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_93),
.A2(n_96),
.B1(n_98),
.B2(n_100),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_64),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

BUFx2_ASAP7_75t_SL g95 ( 
.A(n_55),
.Y(n_95)
);

INVx6_ASAP7_75t_SL g114 ( 
.A(n_95),
.Y(n_114)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_22),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_97),
.B(n_17),
.Y(n_108)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_67),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_80),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_105),
.A2(n_129),
.B1(n_86),
.B2(n_46),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_108),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_119),
.A2(n_126),
.B(n_128),
.Y(n_148)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_120),
.Y(n_142)
);

INVx6_ASAP7_75t_SL g121 ( 
.A(n_84),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_121),
.A2(n_90),
.B1(n_43),
.B2(n_46),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_82),
.C(n_41),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_127),
.B1(n_90),
.B2(n_93),
.Y(n_135)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_78),
.A2(n_57),
.B(n_24),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_81),
.A2(n_40),
.B1(n_43),
.B2(n_41),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_41),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_80),
.A2(n_40),
.B1(n_19),
.B2(n_29),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_76),
.A2(n_62),
.B1(n_29),
.B2(n_19),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_131),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_135),
.A2(n_47),
.B1(n_45),
.B2(n_28),
.Y(n_190)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_132),
.Y(n_161)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_139),
.B(n_156),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_104),
.B(n_78),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_144),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_101),
.A2(n_87),
.B1(n_82),
.B2(n_79),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_147),
.B1(n_117),
.B2(n_102),
.Y(n_166)
);

NOR2x1_ASAP7_75t_R g145 ( 
.A(n_101),
.B(n_80),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_150),
.B(n_154),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_109),
.A2(n_118),
.B1(n_122),
.B2(n_132),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_45),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_21),
.B(n_20),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_114),
.A2(n_110),
.B1(n_127),
.B2(n_125),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_151),
.A2(n_155),
.B1(n_158),
.B2(n_124),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_152),
.A2(n_106),
.B1(n_116),
.B2(n_131),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_73),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_159),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_73),
.B(n_21),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_114),
.A2(n_21),
.B1(n_32),
.B2(n_29),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_157),
.B(n_18),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_21),
.B1(n_32),
.B2(n_33),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_109),
.B(n_18),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_105),
.B1(n_118),
.B2(n_122),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_160),
.A2(n_166),
.B1(n_183),
.B2(n_184),
.Y(n_207)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_128),
.B(n_107),
.C(n_102),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_162),
.A2(n_170),
.B(n_177),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_121),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_164),
.B(n_168),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_165),
.A2(n_187),
.B1(n_134),
.B2(n_137),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_140),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_167),
.Y(n_201)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_169),
.B(n_171),
.Y(n_220)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_108),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_177),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_142),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_176),
.Y(n_210)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_115),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_154),
.A2(n_21),
.B(n_32),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_178),
.A2(n_24),
.B(n_18),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_135),
.Y(n_179)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_45),
.Y(n_197)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_133),
.Y(n_203)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_117),
.B1(n_115),
.B2(n_120),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_106),
.Y(n_185)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_134),
.A2(n_99),
.B1(n_72),
.B2(n_33),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_140),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_188),
.Y(n_205)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_189),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_26),
.B1(n_34),
.B2(n_28),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_191),
.A2(n_215),
.B1(n_171),
.B2(n_187),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_149),
.C(n_148),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_206),
.C(n_208),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_145),
.B1(n_151),
.B2(n_157),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_194),
.A2(n_196),
.B1(n_211),
.B2(n_219),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_166),
.A2(n_158),
.B1(n_155),
.B2(n_139),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_197),
.B(n_186),
.Y(n_240)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_182),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_172),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_156),
.C(n_47),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_45),
.C(n_137),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_181),
.A2(n_36),
.B1(n_17),
.B2(n_31),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_18),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_178),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_1),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_213),
.A2(n_216),
.B(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_173),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_26),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_18),
.C(n_36),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_169),
.C(n_173),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_167),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_218),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_165),
.A2(n_31),
.B1(n_27),
.B2(n_28),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_162),
.A2(n_27),
.B1(n_28),
.B2(n_34),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_221),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_222),
.A2(n_24),
.B(n_34),
.Y(n_248)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_228),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_238),
.Y(n_260)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_168),
.Y(n_229)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_229),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_239),
.C(n_217),
.Y(n_252)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_234),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_L g233 ( 
.A1(n_220),
.A2(n_216),
.B(n_209),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_233),
.A2(n_236),
.B(n_241),
.Y(n_262)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_235),
.A2(n_247),
.B1(n_219),
.B2(n_192),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_SL g236 ( 
.A1(n_207),
.A2(n_201),
.B(n_205),
.C(n_191),
.Y(n_236)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_193),
.B(n_189),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_188),
.C(n_183),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_24),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_199),
.B(n_186),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_243),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_34),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_24),
.Y(n_261)
);

NAND3xp33_ASAP7_75t_L g245 ( 
.A(n_204),
.B(n_11),
.C(n_16),
.Y(n_245)
);

BUFx12f_ASAP7_75t_SL g269 ( 
.A(n_245),
.Y(n_269)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_200),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_229),
.B(n_223),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_251),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_230),
.C(n_260),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_225),
.B(n_194),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_254),
.B(n_240),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_241),
.A2(n_199),
.B1(n_196),
.B2(n_202),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_255),
.A2(n_256),
.B1(n_259),
.B2(n_236),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_246),
.A2(n_195),
.B1(n_212),
.B2(n_213),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_239),
.A2(n_211),
.B1(n_213),
.B2(n_222),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_263),
.B1(n_227),
.B2(n_231),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_246),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_268),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_236),
.A2(n_2),
.B(n_3),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_265),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_236),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_267)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_269),
.C(n_5),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_230),
.C(n_238),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_279),
.C(n_261),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_249),
.B(n_226),
.Y(n_272)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_233),
.Y(n_274)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_265),
.Y(n_275)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_275),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_268),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_254),
.C(n_264),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_282),
.Y(n_294)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_250),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_244),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_283),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_286),
.B(n_257),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_258),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_262),
.A2(n_248),
.B1(n_6),
.B2(n_8),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_281),
.B1(n_259),
.B2(n_269),
.Y(n_288)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

XOR2x2_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_262),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_289),
.B(n_280),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_274),
.A2(n_278),
.B1(n_285),
.B2(n_277),
.Y(n_291)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_291),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_299),
.C(n_302),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_298),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_255),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_256),
.C(n_263),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_311),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_286),
.B1(n_271),
.B2(n_276),
.Y(n_308)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_308),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_276),
.C(n_5),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_298),
.C(n_10),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_289),
.A2(n_300),
.B(n_294),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_6),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_312),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_8),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_314),
.Y(n_321)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_291),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_305),
.B(n_297),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_304),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_303),
.A2(n_301),
.B1(n_299),
.B2(n_302),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_322),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_320),
.B(n_323),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_306),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_10),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_316),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_317),
.B(n_309),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_325),
.B(n_12),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_309),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_327),
.A2(n_328),
.B(n_329),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_304),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_310),
.Y(n_329)
);

OAI21x1_ASAP7_75t_L g336 ( 
.A1(n_331),
.A2(n_324),
.B(n_13),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_320),
.C(n_319),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_332),
.A2(n_334),
.B(n_326),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_335),
.Y(n_337)
);

O2A1O1Ixp33_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_336),
.B(n_333),
.C(n_331),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_12),
.B(n_13),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_12),
.B(n_14),
.Y(n_340)
);

MAJx2_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_14),
.C(n_15),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_15),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_15),
.Y(n_343)
);


endmodule