module fake_jpeg_22505_n_222 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_222);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_7),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_38),
.B1(n_26),
.B2(n_28),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_7),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_24),
.B1(n_29),
.B2(n_20),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_41),
.Y(n_43)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_53),
.B1(n_40),
.B2(n_37),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_15),
.B1(n_18),
.B2(n_22),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_52),
.B1(n_30),
.B2(n_17),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

AO22x1_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_15),
.B1(n_18),
.B2(n_24),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_25),
.B1(n_17),
.B2(n_19),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_19),
.B1(n_17),
.B2(n_25),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_31),
.B1(n_23),
.B2(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_33),
.Y(n_70)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_36),
.C(n_34),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_72),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_67),
.B(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_71),
.A2(n_77),
.B1(n_80),
.B2(n_63),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_36),
.C(n_34),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_73),
.A2(n_79),
.B1(n_50),
.B2(n_45),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_40),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_83),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_10),
.B1(n_2),
.B2(n_3),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_40),
.B(n_37),
.C(n_36),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_8),
.B1(n_2),
.B2(n_4),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_64),
.B1(n_60),
.B2(n_47),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_50),
.B1(n_45),
.B2(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_37),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_44),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_85),
.B(n_89),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_62),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_65),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_43),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_91),
.B(n_95),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_92),
.A2(n_100),
.B1(n_71),
.B2(n_72),
.Y(n_108)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_43),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_76),
.B1(n_61),
.B2(n_69),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_68),
.B(n_53),
.Y(n_98)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_68),
.B(n_44),
.Y(n_99)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_1),
.Y(n_103)
);

NAND2x1_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_5),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_67),
.B(n_4),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_104),
.B(n_5),
.Y(n_115)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_101),
.B(n_73),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_103),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_108),
.A2(n_122),
.B1(n_125),
.B2(n_127),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_115),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_91),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_112),
.A2(n_98),
.B1(n_86),
.B2(n_87),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_47),
.A3(n_76),
.B1(n_69),
.B2(n_55),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_97),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_47),
.B1(n_84),
.B2(n_81),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_124),
.B(n_89),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_102),
.A2(n_81),
.B1(n_57),
.B2(n_12),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_95),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_86),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_100),
.A2(n_81),
.B1(n_11),
.B2(n_12),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_96),
.C(n_101),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_130),
.C(n_123),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_129),
.B(n_124),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_96),
.C(n_90),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVxp67_ASAP7_75t_SL g163 ( 
.A(n_131),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_85),
.B(n_93),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_134),
.B(n_117),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_94),
.B(n_99),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_87),
.Y(n_135)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_138),
.Y(n_150)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_146),
.Y(n_157)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_147),
.Y(n_161)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_121),
.A2(n_103),
.B1(n_104),
.B2(n_13),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_134),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_162),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_151),
.A2(n_6),
.B(n_11),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_138),
.A2(n_121),
.B1(n_118),
.B2(n_114),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_152),
.A2(n_13),
.B1(n_14),
.B2(n_149),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_159),
.C(n_130),
.Y(n_165)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_124),
.C(n_129),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_117),
.C(n_108),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_160),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_156),
.C(n_159),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_118),
.B1(n_127),
.B2(n_144),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_170),
.B1(n_176),
.B2(n_14),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_157),
.Y(n_185)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_139),
.A3(n_142),
.B1(n_146),
.B2(n_135),
.C1(n_140),
.C2(n_114),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_169),
.B(n_179),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_122),
.B1(n_131),
.B2(n_142),
.Y(n_170)
);

AOI321xp33_ASAP7_75t_L g171 ( 
.A1(n_158),
.A2(n_120),
.A3(n_133),
.B1(n_126),
.B2(n_137),
.C(n_147),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_171),
.A2(n_177),
.B(n_178),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_150),
.Y(n_172)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_161),
.B(n_136),
.Y(n_174)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_174),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_115),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_152),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_6),
.B1(n_11),
.B2(n_13),
.Y(n_176)
);

NAND2x1_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_6),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_SL g180 ( 
.A(n_168),
.B(n_161),
.C(n_157),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_180),
.B(n_174),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_183),
.B(n_189),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_171),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_178),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_178),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_188),
.C(n_190),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_153),
.C(n_154),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_166),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_197),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_183),
.A2(n_166),
.B(n_173),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_194),
.A2(n_188),
.B(n_184),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_185),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_182),
.A2(n_173),
.B1(n_167),
.B2(n_170),
.Y(n_197)
);

XOR2x2_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_187),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_181),
.B(n_179),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_180),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_175),
.B1(n_177),
.B2(n_176),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_200),
.A2(n_186),
.B1(n_190),
.B2(n_191),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_207),
.B1(n_195),
.B2(n_196),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_191),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_198),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_205),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_206),
.B(n_192),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_212),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_201),
.B(n_195),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_209),
.B(n_210),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_203),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_215),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_207),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_204),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_218),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_217),
.A2(n_216),
.B(n_205),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_216),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_219),
.Y(n_222)
);


endmodule