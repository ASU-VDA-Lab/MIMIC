module fake_ariane_2219_n_197 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_30, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_197);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_30;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_197;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_195;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_82;
wire n_178;
wire n_42;
wire n_31;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_144;
wire n_130;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_188;
wire n_185;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_41;
wire n_140;
wire n_55;
wire n_191;
wire n_151;
wire n_136;
wire n_192;
wire n_80;
wire n_146;
wire n_194;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_193;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVxp67_ASAP7_75t_SL g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

INVxp33_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_0),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

OA21x2_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_1),
.B(n_2),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_3),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_5),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_56),
.B(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_38),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_51),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_43),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_34),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

AND2x4_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_5),
.Y(n_88)
);

AO22x2_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_49),
.B1(n_40),
.B2(n_45),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g92 ( 
.A(n_75),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_62),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_85),
.B(n_68),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_60),
.Y(n_96)
);

AND3x1_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_72),
.C(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

AOI221xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_60),
.B1(n_37),
.B2(n_47),
.C(n_72),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_74),
.B1(n_92),
.B2(n_97),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_98),
.A2(n_82),
.B(n_84),
.C(n_80),
.Y(n_106)
);

O2A1O1Ixp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_83),
.B(n_84),
.C(n_88),
.Y(n_107)
);

AOI21x1_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_88),
.B(n_97),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_81),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_80),
.Y(n_110)
);

OA21x2_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_101),
.B(n_99),
.Y(n_111)
);

NOR3xp33_ASAP7_75t_SL g112 ( 
.A(n_108),
.B(n_100),
.C(n_95),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_74),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

OAI21x1_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_91),
.B(n_101),
.Y(n_116)
);

OA21x2_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_99),
.B(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

OA21x2_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_107),
.B(n_105),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_118),
.A2(n_113),
.B(n_109),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_102),
.C(n_114),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_122),
.Y(n_130)
);

NAND4xp25_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_110),
.C(n_109),
.D(n_71),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_96),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_133),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_125),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_96),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_127),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_125),
.Y(n_146)
);

NAND2x1_ASAP7_75t_SL g147 ( 
.A(n_140),
.B(n_129),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

AOI222xp33_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_113),
.B1(n_89),
.B2(n_116),
.C1(n_88),
.C2(n_80),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_128),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_128),
.Y(n_151)
);

NOR2xp67_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_130),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_138),
.Y(n_153)
);

NOR2x1_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_146),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

NAND2xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_112),
.Y(n_156)
);

NAND3xp33_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_112),
.C(n_63),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

NOR2x1_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_131),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_113),
.B(n_116),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_149),
.C(n_63),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_143),
.Y(n_165)
);

NOR2x1p5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_67),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_67),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_142),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_113),
.B1(n_89),
.B2(n_88),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_122),
.B(n_106),
.Y(n_170)
);

AOI221x1_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_89),
.B1(n_64),
.B2(n_70),
.C(n_66),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

NOR3x1_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_165),
.C(n_168),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_64),
.C(n_70),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_162),
.A2(n_122),
.B(n_117),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_170),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_66),
.Y(n_177)
);

NOR2x1_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_81),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

AOI221xp5_ASAP7_75t_L g180 ( 
.A1(n_175),
.A2(n_63),
.B1(n_58),
.B2(n_59),
.C(n_88),
.Y(n_180)
);

NAND4xp25_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_59),
.C(n_58),
.D(n_9),
.Y(n_181)
);

AOI221xp5_ASAP7_75t_L g182 ( 
.A1(n_175),
.A2(n_79),
.B1(n_87),
.B2(n_76),
.C(n_90),
.Y(n_182)
);

NAND4xp75_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_74),
.C(n_56),
.D(n_117),
.Y(n_183)
);

AOI221xp5_ASAP7_75t_SL g184 ( 
.A1(n_172),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.C(n_10),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_76),
.B1(n_56),
.B2(n_90),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_174),
.B(n_76),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_178),
.B1(n_56),
.B2(n_90),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_10),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_117),
.B1(n_111),
.B2(n_87),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_184),
.A2(n_117),
.B1(n_111),
.B2(n_79),
.Y(n_190)
);

AOI221xp5_ASAP7_75t_L g191 ( 
.A1(n_182),
.A2(n_11),
.B1(n_13),
.B2(n_16),
.C(n_17),
.Y(n_191)
);

OAI222xp33_ASAP7_75t_L g192 ( 
.A1(n_190),
.A2(n_185),
.B1(n_186),
.B2(n_183),
.C1(n_117),
.C2(n_111),
.Y(n_192)
);

AND4x1_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_18),
.C(n_21),
.D(n_23),
.Y(n_193)
);

O2A1O1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_191),
.A2(n_111),
.B(n_117),
.C(n_29),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_192),
.A2(n_188),
.B(n_189),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_194),
.A2(n_111),
.B(n_28),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_195),
.A2(n_196),
.B1(n_193),
.B2(n_30),
.Y(n_197)
);


endmodule