module fake_jpeg_22354_n_47 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_17),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_10),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_18),
.A2(n_19),
.B(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_21),
.B(n_9),
.Y(n_25)
);

OR2x4_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_2),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_2),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_23),
.B(n_5),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_25),
.B(n_18),
.Y(n_34)
);

OAI322xp33_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_27),
.A3(n_0),
.B1(n_1),
.B2(n_24),
.C1(n_25),
.C2(n_28),
.Y(n_38)
);

AND2x6_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_5),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_12),
.B1(n_7),
.B2(n_11),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_4),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_15),
.A2(n_7),
.B1(n_11),
.B2(n_12),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_19),
.A2(n_11),
.B1(n_2),
.B2(n_4),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_17),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_26),
.C(n_29),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_38),
.Y(n_40)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_36),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_0),
.B1(n_1),
.B2(n_16),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_40),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_35),
.B1(n_33),
.B2(n_36),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_39),
.B1(n_45),
.B2(n_44),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);


endmodule