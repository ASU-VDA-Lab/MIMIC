module fake_jpeg_17877_n_233 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_233);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx5_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_33),
.B(n_20),
.Y(n_64)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_41),
.A2(n_15),
.B1(n_30),
.B2(n_23),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_43),
.A2(n_51),
.B1(n_53),
.B2(n_57),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_30),
.B1(n_15),
.B2(n_31),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_47),
.B1(n_52),
.B2(n_58),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_31),
.B1(n_18),
.B2(n_26),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_18),
.B1(n_26),
.B2(n_24),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_29),
.B1(n_22),
.B2(n_27),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_39),
.B1(n_34),
.B2(n_29),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_35),
.B1(n_33),
.B2(n_20),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_19),
.B1(n_28),
.B2(n_16),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_27),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_60),
.B(n_17),
.Y(n_65)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_16),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_0),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_65),
.B(n_77),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_40),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_73),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_64),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_76),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_34),
.B1(n_42),
.B2(n_37),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_69),
.A2(n_79),
.B1(n_55),
.B2(n_50),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_36),
.B(n_17),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_72),
.A2(n_81),
.B(n_84),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_40),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

OR2x2_ASAP7_75t_SL g76 ( 
.A(n_63),
.B(n_32),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_40),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_48),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_SL g79 ( 
.A1(n_49),
.A2(n_32),
.B(n_40),
.C(n_37),
.Y(n_79)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_32),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_83),
.B(n_1),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_14),
.B(n_13),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_62),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_93),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_37),
.C(n_46),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_82),
.C(n_62),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_81),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_106),
.B1(n_55),
.B2(n_66),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_103),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_32),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_79),
.B(n_81),
.Y(n_112)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_1),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_99),
.A2(n_2),
.B(n_3),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_74),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_102),
.Y(n_113)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_44),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_44),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_71),
.A2(n_55),
.B1(n_50),
.B2(n_34),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_94),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_112),
.A2(n_117),
.B(n_118),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_122),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_71),
.B1(n_82),
.B2(n_79),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_121),
.B1(n_96),
.B2(n_92),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_72),
.B(n_76),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_66),
.B(n_70),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_87),
.A2(n_1),
.B(n_2),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_124),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_100),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_99),
.A2(n_80),
.B1(n_85),
.B2(n_4),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_80),
.Y(n_125)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_104),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_46),
.C(n_42),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_90),
.Y(n_136)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_4),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_96),
.B1(n_101),
.B2(n_86),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_88),
.B(n_42),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_130),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_120),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_135),
.Y(n_166)
);

AO22x1_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_99),
.B1(n_95),
.B2(n_98),
.Y(n_133)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_133),
.A2(n_149),
.B(n_126),
.Y(n_157)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_108),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_139),
.C(n_148),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_151),
.Y(n_168)
);

OAI32xp33_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_86),
.A3(n_106),
.B1(n_108),
.B2(n_98),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_124),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_118),
.B(n_109),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_115),
.B(n_129),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_150),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_117),
.Y(n_148)
);

OAI22x1_ASAP7_75t_SL g149 ( 
.A1(n_116),
.A2(n_97),
.B1(n_102),
.B2(n_42),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_97),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_152),
.B(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_164),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_132),
.B(n_144),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_156),
.A2(n_159),
.B(n_100),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_157),
.A2(n_107),
.B1(n_102),
.B2(n_46),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_110),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_139),
.C(n_113),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_129),
.B(n_111),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

NOR3xp33_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_134),
.C(n_132),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_114),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_140),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_113),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_127),
.Y(n_169)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_172),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_121),
.C(n_122),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_175),
.B(n_181),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_163),
.B(n_169),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_178),
.A2(n_164),
.B(n_154),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_161),
.B1(n_163),
.B2(n_166),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_5),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_6),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_183),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_12),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_12),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_13),
.Y(n_197)
);

AOI21x1_ASAP7_75t_L g186 ( 
.A1(n_178),
.A2(n_156),
.B(n_165),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_188),
.B(n_161),
.Y(n_201)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_176),
.Y(n_187)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_152),
.B(n_159),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_189),
.A2(n_193),
.B(n_185),
.Y(n_203)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

BUFx12_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_195),
.Y(n_204)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_182),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_199),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_205),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_201),
.A2(n_189),
.B(n_165),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_153),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_171),
.C(n_173),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_157),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_173),
.C(n_165),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_194),
.C(n_192),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

AOI21x1_ASAP7_75t_L g210 ( 
.A1(n_206),
.A2(n_165),
.B(n_157),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_211),
.C(n_214),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_155),
.B1(n_204),
.B2(n_198),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_199),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_192),
.C(n_194),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_214),
.B(n_196),
.Y(n_216)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_216),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_221),
.C(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_160),
.C(n_8),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_6),
.C(n_8),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_212),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_217),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_227),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_209),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_228),
.Y(n_230)
);

AOI321xp33_ASAP7_75t_L g231 ( 
.A1(n_229),
.A2(n_8),
.A3(n_10),
.B1(n_222),
.B2(n_219),
.C(n_176),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_230),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g233 ( 
.A(n_232),
.Y(n_233)
);


endmodule