module fake_jpeg_12846_n_98 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_98);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_98;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_2),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_30),
.B(n_2),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_37),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_3),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_34),
.B1(n_33),
.B2(n_31),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_36),
.B1(n_29),
.B2(n_20),
.Y(n_64)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_66),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_55),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_48),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_39),
.C(n_29),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_4),
.C(n_5),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_34),
.B1(n_33),
.B2(n_39),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_64),
.B1(n_65),
.B2(n_21),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_36),
.B1(n_4),
.B2(n_5),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_3),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_54),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_72),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_80),
.B(n_81),
.Y(n_84)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_6),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_79),
.A2(n_62),
.B1(n_6),
.B2(n_11),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_28),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_82),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_73),
.C(n_12),
.Y(n_91)
);

INVxp67_ASAP7_75t_SL g89 ( 
.A(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_90),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_92),
.B(n_86),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_84),
.Y(n_94)
);

AOI31xp33_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_82),
.A3(n_85),
.B(n_91),
.Y(n_95)
);

AOI322xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_88),
.A3(n_87),
.B1(n_14),
.B2(n_19),
.C1(n_22),
.C2(n_9),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_13),
.C(n_23),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_25),
.Y(n_98)
);


endmodule