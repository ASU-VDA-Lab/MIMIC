module fake_jpeg_2100_n_53 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_53);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_53;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_6),
.B(n_2),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx16_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_22),
.A2(n_23),
.B(n_10),
.Y(n_29)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_25),
.C(n_27),
.Y(n_31)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_10),
.B1(n_22),
.B2(n_20),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_0),
.Y(n_27)
);

INVxp67_ASAP7_75t_SL g38 ( 
.A(n_29),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_24),
.A2(n_12),
.B1(n_11),
.B2(n_17),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_34),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_18),
.A2(n_16),
.B1(n_17),
.B2(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_35),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_25),
.A2(n_16),
.B1(n_14),
.B2(n_7),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_18),
.A2(n_4),
.B1(n_6),
.B2(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_36),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_41),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_26),
.B(n_21),
.Y(n_41)
);

MAJx2_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_31),
.C(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_44),
.Y(n_48)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_32),
.B1(n_34),
.B2(n_30),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

AO21x1_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_50),
.B(n_47),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_39),
.B1(n_41),
.B2(n_40),
.Y(n_53)
);


endmodule