module fake_jpeg_30881_n_91 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_91);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_91;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_13),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_1),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_2),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_50),
.A2(n_51),
.B1(n_53),
.B2(n_36),
.Y(n_57)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

AO22x1_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_28),
.B1(n_38),
.B2(n_37),
.Y(n_56)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_42),
.B(n_3),
.Y(n_66)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_39),
.B1(n_40),
.B2(n_30),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_59),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_29),
.B1(n_31),
.B2(n_27),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_54),
.B(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_64),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_65),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_68),
.B1(n_60),
.B2(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_2),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_3),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_61),
.B1(n_44),
.B2(n_60),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_69),
.B1(n_5),
.B2(n_4),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_75),
.B(n_76),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_74),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_77),
.C(n_72),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_77),
.B(n_69),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_82),
.C(n_80),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_11),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_10),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_5),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_85),
.A2(n_7),
.B(n_8),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_SL g89 ( 
.A(n_86),
.B(n_12),
.C(n_15),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

BUFx24_ASAP7_75t_SL g90 ( 
.A(n_89),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_90),
.B(n_88),
.Y(n_91)
);


endmodule