module fake_aes_3619_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx6f_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
AND2x4_ASAP7_75t_L g12 ( .A(n_4), .B(n_6), .Y(n_12) );
BUFx6f_ASAP7_75t_L g13 ( .A(n_3), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_10), .B(n_1), .Y(n_14) );
AND2x4_ASAP7_75t_L g15 ( .A(n_8), .B(n_0), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_2), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_16), .B(n_0), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_12), .B(n_1), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_12), .B(n_2), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_14), .B(n_15), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_17), .Y(n_21) );
INVx1_ASAP7_75t_SL g22 ( .A(n_21), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_20), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_23), .B(n_21), .Y(n_25) );
NOR2x1_ASAP7_75t_L g26 ( .A(n_24), .B(n_19), .Y(n_26) );
NAND2xp5_ASAP7_75t_SL g27 ( .A(n_24), .B(n_20), .Y(n_27) );
NOR2x1_ASAP7_75t_L g28 ( .A(n_26), .B(n_25), .Y(n_28) );
OAI321xp33_ASAP7_75t_L g29 ( .A1(n_27), .A2(n_14), .A3(n_11), .B1(n_13), .B2(n_25), .C(n_3), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
O2A1O1Ixp33_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_15), .B(n_20), .C(n_13), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_28), .B(n_13), .Y(n_32) );
AO22x2_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_11), .B1(n_7), .B2(n_9), .Y(n_33) );
NOR2xp33_ASAP7_75t_R g34 ( .A(n_32), .B(n_5), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
AOI22xp33_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_34), .B1(n_11), .B2(n_31), .Y(n_36) );
endmodule