module fake_netlist_1_8032_n_744 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_744);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_744;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_721;
wire n_134;
wire n_438;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_33), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_31), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_74), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_64), .Y(n_85) );
BUFx3_ASAP7_75t_L g86 ( .A(n_79), .Y(n_86) );
HB1xp67_ASAP7_75t_L g87 ( .A(n_9), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_68), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_72), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_7), .Y(n_90) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_55), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_75), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_35), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_34), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_54), .Y(n_95) );
BUFx6f_ASAP7_75t_L g96 ( .A(n_45), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_66), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_29), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_71), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_76), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_47), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_27), .Y(n_102) );
CKINVDCx14_ASAP7_75t_R g103 ( .A(n_48), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_60), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_43), .Y(n_105) );
NOR2xp67_ASAP7_75t_L g106 ( .A(n_2), .B(n_67), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_38), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_3), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_65), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_14), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_69), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_5), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_77), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_46), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_5), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_22), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_52), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_12), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_73), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_1), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_18), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_12), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_21), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_14), .Y(n_125) );
BUFx2_ASAP7_75t_L g126 ( .A(n_62), .Y(n_126) );
BUFx2_ASAP7_75t_SL g127 ( .A(n_49), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_11), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_37), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_40), .Y(n_130) );
CKINVDCx16_ASAP7_75t_R g131 ( .A(n_58), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_126), .B(n_0), .Y(n_132) );
OAI22xp5_ASAP7_75t_SL g133 ( .A1(n_110), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_91), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_126), .B(n_4), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_91), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_91), .B(n_4), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_87), .B(n_6), .Y(n_138) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_110), .Y(n_139) );
OAI22xp33_ASAP7_75t_R g140 ( .A1(n_90), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_140) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_111), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_105), .B(n_8), .Y(n_142) );
INVx6_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
INVxp67_ASAP7_75t_L g144 ( .A(n_113), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_93), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_131), .B(n_9), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_86), .B(n_10), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_91), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_91), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_116), .B(n_10), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_88), .B(n_11), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_96), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_93), .Y(n_153) );
OAI22xp5_ASAP7_75t_SL g154 ( .A1(n_111), .A2(n_13), .B1(n_15), .B2(n_16), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_96), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_96), .Y(n_156) );
INVx2_ASAP7_75t_SL g157 ( .A(n_88), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_121), .B(n_13), .Y(n_158) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_94), .A2(n_41), .B(n_80), .Y(n_159) );
INVx4_ASAP7_75t_L g160 ( .A(n_96), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_94), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_96), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_115), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_122), .B(n_15), .Y(n_164) );
AOI22x1_ASAP7_75t_SL g165 ( .A1(n_128), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_95), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_115), .Y(n_167) );
AND2x6_ASAP7_75t_L g168 ( .A(n_95), .B(n_42), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_123), .B(n_17), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_125), .B(n_19), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_118), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_118), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_130), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_83), .B(n_19), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_130), .Y(n_175) );
BUFx2_ASAP7_75t_L g176 ( .A(n_128), .Y(n_176) );
NAND2xp33_ASAP7_75t_L g177 ( .A(n_168), .B(n_129), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_176), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_176), .B(n_104), .Y(n_179) );
INVx5_ASAP7_75t_L g180 ( .A(n_168), .Y(n_180) );
INVxp67_ASAP7_75t_SL g181 ( .A(n_135), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_143), .Y(n_182) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_151), .A2(n_103), .B1(n_127), .B2(n_108), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_151), .Y(n_184) );
INVx1_ASAP7_75t_SL g185 ( .A(n_139), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_132), .B(n_106), .Y(n_186) );
OR2x6_ASAP7_75t_L g187 ( .A(n_133), .B(n_127), .Y(n_187) );
INVxp33_ASAP7_75t_L g188 ( .A(n_141), .Y(n_188) );
INVx1_ASAP7_75t_SL g189 ( .A(n_142), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_151), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_132), .A2(n_84), .B1(n_100), .B2(n_102), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_147), .B(n_85), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_145), .B(n_89), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_151), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_143), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_145), .B(n_82), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_166), .B(n_107), .Y(n_197) );
INVx2_ASAP7_75t_SL g198 ( .A(n_142), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_144), .B(n_98), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_166), .B(n_109), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_153), .B(n_99), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_143), .Y(n_202) );
AND2x6_ASAP7_75t_L g203 ( .A(n_147), .B(n_112), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_153), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_144), .B(n_101), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_172), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_147), .B(n_114), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_147), .B(n_114), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_138), .A2(n_119), .B1(n_124), .B2(n_120), .Y(n_209) );
INVx1_ASAP7_75t_SL g210 ( .A(n_146), .Y(n_210) );
INVxp67_ASAP7_75t_L g211 ( .A(n_146), .Y(n_211) );
OR2x6_ASAP7_75t_L g212 ( .A(n_133), .B(n_117), .Y(n_212) );
NAND2xp33_ASAP7_75t_L g213 ( .A(n_168), .B(n_129), .Y(n_213) );
BUFx10_ASAP7_75t_L g214 ( .A(n_157), .Y(n_214) );
BUFx4f_ASAP7_75t_L g215 ( .A(n_168), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_153), .B(n_102), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_153), .B(n_104), .Y(n_217) );
AND2x6_ASAP7_75t_L g218 ( .A(n_161), .B(n_97), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_161), .B(n_92), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_143), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_175), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_161), .Y(n_222) );
INVx1_ASAP7_75t_SL g223 ( .A(n_135), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_161), .B(n_92), .Y(n_224) );
HB1xp67_ASAP7_75t_SL g225 ( .A(n_168), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_157), .B(n_97), .Y(n_226) );
AND2x6_ASAP7_75t_L g227 ( .A(n_138), .B(n_82), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_157), .B(n_20), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_173), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_173), .B(n_23), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_143), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_173), .Y(n_232) );
BUFx10_ASAP7_75t_L g233 ( .A(n_168), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_163), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_163), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_163), .Y(n_236) );
INVx4_ASAP7_75t_L g237 ( .A(n_168), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_167), .Y(n_238) );
AND2x2_ASAP7_75t_SL g239 ( .A(n_174), .B(n_24), .Y(n_239) );
OR2x2_ASAP7_75t_L g240 ( .A(n_150), .B(n_25), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_167), .B(n_26), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_167), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_175), .B(n_28), .Y(n_243) );
NOR2x2_ASAP7_75t_L g244 ( .A(n_187), .B(n_140), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_181), .B(n_174), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_233), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_233), .Y(n_247) );
AOI22xp33_ASAP7_75t_SL g248 ( .A1(n_212), .A2(n_165), .B1(n_154), .B2(n_169), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_223), .B(n_217), .Y(n_249) );
NOR2xp67_ASAP7_75t_L g250 ( .A(n_178), .B(n_171), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_184), .A2(n_168), .B1(n_171), .B2(n_175), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_223), .B(n_217), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_219), .B(n_158), .Y(n_253) );
INVx2_ASAP7_75t_SL g254 ( .A(n_214), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_237), .B(n_158), .Y(n_255) );
AOI221xp5_ASAP7_75t_L g256 ( .A1(n_189), .A2(n_154), .B1(n_170), .B2(n_169), .C(n_164), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_214), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_182), .Y(n_258) );
INVx2_ASAP7_75t_SL g259 ( .A(n_185), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_184), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_204), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_237), .B(n_164), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_202), .Y(n_263) );
NAND2x1p5_ASAP7_75t_L g264 ( .A(n_185), .B(n_137), .Y(n_264) );
NAND3xp33_ASAP7_75t_SL g265 ( .A(n_183), .B(n_170), .C(n_150), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_199), .B(n_171), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_179), .B(n_175), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_195), .Y(n_268) );
OR2x6_ASAP7_75t_L g269 ( .A(n_187), .B(n_140), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_215), .B(n_175), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_220), .Y(n_271) );
OAI22xp5_ASAP7_75t_SL g272 ( .A1(n_212), .A2(n_165), .B1(n_159), .B2(n_175), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_215), .B(n_172), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_188), .B(n_160), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_189), .Y(n_275) );
OAI22xp5_ASAP7_75t_SL g276 ( .A1(n_212), .A2(n_159), .B1(n_172), .B2(n_160), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_222), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_205), .B(n_160), .Y(n_278) );
INVx4_ASAP7_75t_L g279 ( .A(n_218), .Y(n_279) );
INVx2_ASAP7_75t_SL g280 ( .A(n_227), .Y(n_280) );
INVx8_ASAP7_75t_L g281 ( .A(n_203), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_186), .B(n_160), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_186), .B(n_172), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_190), .A2(n_172), .B1(n_159), .B2(n_162), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_211), .B(n_172), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_198), .B(n_162), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_207), .B(n_159), .Y(n_287) );
NAND3xp33_ASAP7_75t_SL g288 ( .A(n_210), .B(n_162), .C(n_155), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_227), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_191), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_196), .B(n_159), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_231), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_180), .B(n_156), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_194), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_180), .Y(n_295) );
INVx2_ASAP7_75t_SL g296 ( .A(n_227), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_226), .B(n_155), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_210), .A2(n_155), .B1(n_152), .B2(n_149), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_192), .B(n_152), .Y(n_299) );
NAND2x1p5_ASAP7_75t_L g300 ( .A(n_239), .B(n_152), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_208), .B(n_30), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_227), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_216), .B(n_32), .Y(n_303) );
INVxp67_ASAP7_75t_L g304 ( .A(n_218), .Y(n_304) );
INVxp67_ASAP7_75t_SL g305 ( .A(n_192), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_229), .Y(n_306) );
INVx4_ASAP7_75t_L g307 ( .A(n_218), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_218), .B(n_149), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_224), .B(n_149), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_234), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_203), .B(n_148), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_209), .B(n_148), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_193), .B(n_148), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_225), .A2(n_134), .B1(n_156), .B2(n_136), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_203), .A2(n_134), .B1(n_136), .B2(n_156), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_254), .B(n_228), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_287), .A2(n_291), .B(n_213), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_245), .B(n_203), .Y(n_318) );
OAI21xp5_ASAP7_75t_L g319 ( .A1(n_291), .A2(n_177), .B(n_180), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_259), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_249), .B(n_240), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_252), .B(n_200), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_275), .B(n_187), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_279), .B(n_180), .Y(n_324) );
BUFx2_ASAP7_75t_R g325 ( .A(n_290), .Y(n_325) );
NOR3xp33_ASAP7_75t_SL g326 ( .A(n_265), .B(n_193), .C(n_197), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_305), .A2(n_200), .B1(n_197), .B2(n_201), .Y(n_327) );
INVx3_ASAP7_75t_SL g328 ( .A(n_281), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_275), .B(n_201), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_257), .Y(n_330) );
AOI22xp5_ASAP7_75t_L g331 ( .A1(n_305), .A2(n_228), .B1(n_232), .B2(n_235), .Y(n_331) );
INVx4_ASAP7_75t_L g332 ( .A(n_281), .Y(n_332) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_279), .B(n_307), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_310), .Y(n_334) );
A2O1A1Ixp33_ASAP7_75t_SL g335 ( .A1(n_283), .A2(n_221), .B(n_242), .C(n_238), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_289), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_250), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_253), .B(n_236), .Y(n_338) );
NAND2xp5_ASAP7_75t_SL g339 ( .A(n_307), .B(n_230), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_276), .A2(n_230), .B(n_241), .Y(n_340) );
A2O1A1Ixp33_ASAP7_75t_L g341 ( .A1(n_294), .A2(n_241), .B(n_221), .C(n_134), .Y(n_341) );
NOR2xp33_ASAP7_75t_SL g342 ( .A(n_281), .B(n_206), .Y(n_342) );
NAND3xp33_ASAP7_75t_SL g343 ( .A(n_248), .B(n_243), .C(n_39), .Y(n_343) );
INVx4_ASAP7_75t_L g344 ( .A(n_295), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_269), .B(n_206), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_260), .Y(n_346) );
INVxp67_ASAP7_75t_L g347 ( .A(n_274), .Y(n_347) );
NOR2xp33_ASAP7_75t_R g348 ( .A(n_302), .B(n_36), .Y(n_348) );
CKINVDCx14_ASAP7_75t_R g349 ( .A(n_269), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_300), .A2(n_206), .B1(n_156), .B2(n_136), .Y(n_350) );
A2O1A1Ixp33_ASAP7_75t_SL g351 ( .A1(n_301), .A2(n_303), .B(n_285), .C(n_267), .Y(n_351) );
AOI21xp5_ASAP7_75t_L g352 ( .A1(n_255), .A2(n_156), .B(n_136), .Y(n_352) );
OAI22xp5_ASAP7_75t_SL g353 ( .A1(n_248), .A2(n_156), .B1(n_136), .B2(n_51), .Y(n_353) );
OAI21xp5_ASAP7_75t_L g354 ( .A1(n_284), .A2(n_136), .B(n_50), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_295), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_265), .B(n_44), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_262), .A2(n_81), .B(n_56), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_269), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_312), .B(n_78), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_264), .B(n_53), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_256), .B(n_70), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_295), .Y(n_362) );
NOR2xp33_ASAP7_75t_R g363 ( .A(n_288), .B(n_57), .Y(n_363) );
NAND2x1p5_ASAP7_75t_L g364 ( .A(n_280), .B(n_63), .Y(n_364) );
AND2x2_ASAP7_75t_SL g365 ( .A(n_244), .B(n_59), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_286), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_268), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_264), .B(n_61), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_300), .B(n_306), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_271), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g371 ( .A1(n_308), .A2(n_284), .B(n_278), .Y(n_371) );
AO21x2_ASAP7_75t_L g372 ( .A1(n_340), .A2(n_288), .B(n_297), .Y(n_372) );
AOI221x1_ASAP7_75t_L g373 ( .A1(n_340), .A2(n_272), .B1(n_314), .B2(n_266), .C(n_286), .Y(n_373) );
BUFx2_ASAP7_75t_L g374 ( .A(n_320), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_321), .A2(n_251), .B1(n_299), .B2(n_296), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_334), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_355), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_329), .B(n_282), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_338), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_322), .B(n_313), .Y(n_380) );
AO31x2_ASAP7_75t_L g381 ( .A1(n_317), .A2(n_277), .A3(n_261), .B(n_292), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_346), .Y(n_382) );
OAI221xp5_ASAP7_75t_L g383 ( .A1(n_323), .A2(n_298), .B1(n_251), .B2(n_309), .C(n_304), .Y(n_383) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_355), .Y(n_384) );
A2O1A1Ixp33_ASAP7_75t_L g385 ( .A1(n_326), .A2(n_304), .B(n_311), .C(n_270), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_327), .B(n_263), .Y(n_386) );
O2A1O1Ixp33_ASAP7_75t_L g387 ( .A1(n_326), .A2(n_273), .B(n_258), .C(n_293), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_317), .A2(n_295), .B(n_247), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_361), .A2(n_315), .B1(n_246), .B2(n_247), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_365), .A2(n_315), .B1(n_246), .B2(n_247), .Y(n_390) );
O2A1O1Ixp33_ASAP7_75t_SL g391 ( .A1(n_356), .A2(n_246), .B(n_247), .C(n_341), .Y(n_391) );
OAI21xp5_ASAP7_75t_L g392 ( .A1(n_371), .A2(n_246), .B(n_319), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_366), .Y(n_393) );
BUFx10_ASAP7_75t_L g394 ( .A(n_330), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_358), .B(n_345), .Y(n_395) );
INVxp67_ASAP7_75t_L g396 ( .A(n_325), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_367), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_353), .A2(n_343), .B1(n_316), .B2(n_369), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_370), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_349), .B(n_328), .Y(n_400) );
A2O1A1Ixp33_ASAP7_75t_SL g401 ( .A1(n_354), .A2(n_347), .B(n_371), .C(n_357), .Y(n_401) );
BUFx8_ASAP7_75t_L g402 ( .A(n_336), .Y(n_402) );
OAI21x1_ASAP7_75t_L g403 ( .A1(n_352), .A2(n_364), .B(n_350), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_337), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_316), .Y(n_405) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_331), .A2(n_343), .B1(n_347), .B2(n_328), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_401), .A2(n_359), .B(n_351), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_379), .A2(n_318), .B1(n_364), .B2(n_368), .Y(n_408) );
O2A1O1Ixp33_ASAP7_75t_L g409 ( .A1(n_379), .A2(n_335), .B(n_360), .C(n_339), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_376), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_376), .B(n_332), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_382), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_397), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_380), .B(n_344), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_401), .A2(n_352), .B(n_357), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_381), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_399), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_378), .B(n_332), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_398), .A2(n_344), .B1(n_362), .B2(n_355), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_398), .A2(n_362), .B1(n_333), .B2(n_363), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_381), .Y(n_421) );
A2O1A1Ixp33_ASAP7_75t_L g422 ( .A1(n_386), .A2(n_387), .B(n_390), .C(n_405), .Y(n_422) );
OAI22xp33_ASAP7_75t_L g423 ( .A1(n_396), .A2(n_342), .B1(n_362), .B2(n_348), .Y(n_423) );
OA21x2_ASAP7_75t_L g424 ( .A1(n_392), .A2(n_324), .B(n_373), .Y(n_424) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_395), .A2(n_404), .B1(n_374), .B2(n_393), .C(n_385), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_381), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_381), .Y(n_427) );
BUFx2_ASAP7_75t_SL g428 ( .A(n_394), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_406), .A2(n_402), .B1(n_394), .B2(n_383), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_400), .B(n_372), .Y(n_430) );
INVx2_ASAP7_75t_SL g431 ( .A(n_402), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_377), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_406), .B(n_384), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_377), .B(n_384), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_372), .B(n_384), .Y(n_435) );
CKINVDCx11_ASAP7_75t_R g436 ( .A(n_384), .Y(n_436) );
OAI211xp5_ASAP7_75t_L g437 ( .A1(n_429), .A2(n_385), .B(n_389), .C(n_391), .Y(n_437) );
AO21x2_ASAP7_75t_L g438 ( .A1(n_407), .A2(n_391), .B(n_388), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_412), .A2(n_375), .B1(n_403), .B2(n_425), .C(n_420), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_410), .B(n_430), .Y(n_440) );
OA21x2_ASAP7_75t_L g441 ( .A1(n_415), .A2(n_427), .B(n_421), .Y(n_441) );
OA21x2_ASAP7_75t_L g442 ( .A1(n_416), .A2(n_427), .B(n_426), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_412), .B(n_430), .Y(n_443) );
OA21x2_ASAP7_75t_L g444 ( .A1(n_416), .A2(n_427), .B(n_426), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_416), .Y(n_445) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_422), .A2(n_420), .B(n_408), .Y(n_446) );
INVx3_ASAP7_75t_L g447 ( .A(n_436), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_421), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_410), .B(n_426), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_421), .Y(n_450) );
AO21x2_ASAP7_75t_L g451 ( .A1(n_433), .A2(n_435), .B(n_408), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_435), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_432), .Y(n_453) );
OA21x2_ASAP7_75t_L g454 ( .A1(n_432), .A2(n_419), .B(n_417), .Y(n_454) );
OR2x6_ASAP7_75t_L g455 ( .A(n_424), .B(n_434), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_424), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_413), .B(n_417), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_413), .B(n_414), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_409), .B(n_424), .C(n_414), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_424), .Y(n_460) );
AO21x2_ASAP7_75t_L g461 ( .A1(n_434), .A2(n_423), .B(n_418), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_428), .A2(n_431), .B1(n_411), .B2(n_434), .Y(n_462) );
INVx2_ASAP7_75t_SL g463 ( .A(n_434), .Y(n_463) );
OAI21xp33_ASAP7_75t_SL g464 ( .A1(n_431), .A2(n_411), .B(n_428), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_411), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_411), .B(n_430), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_416), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_416), .Y(n_468) );
AO21x2_ASAP7_75t_L g469 ( .A1(n_407), .A2(n_415), .B(n_340), .Y(n_469) );
INVxp67_ASAP7_75t_SL g470 ( .A(n_416), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_416), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_412), .B(n_430), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_430), .B(n_379), .Y(n_473) );
BUFx2_ASAP7_75t_L g474 ( .A(n_464), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_473), .B(n_440), .Y(n_475) );
OAI21xp33_ASAP7_75t_SL g476 ( .A1(n_470), .A2(n_450), .B(n_468), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_442), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_450), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_450), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_473), .B(n_440), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_440), .B(n_452), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_452), .B(n_455), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_445), .Y(n_483) );
NOR2xp33_ASAP7_75t_SL g484 ( .A(n_464), .B(n_446), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_440), .B(n_452), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_467), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_452), .B(n_449), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_449), .B(n_466), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_458), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_449), .B(n_466), .Y(n_490) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_446), .A2(n_459), .B(n_469), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_466), .B(n_458), .Y(n_492) );
NOR2x1_ASAP7_75t_R g493 ( .A(n_447), .B(n_464), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_445), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_458), .B(n_472), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_455), .B(n_468), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_445), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_443), .B(n_472), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_443), .B(n_473), .Y(n_499) );
INVxp67_ASAP7_75t_L g500 ( .A(n_470), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_447), .B(n_457), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_467), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_467), .B(n_468), .Y(n_503) );
OAI321xp33_ASAP7_75t_L g504 ( .A1(n_462), .A2(n_437), .A3(n_439), .B1(n_459), .B2(n_465), .C(n_457), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_445), .B(n_471), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_455), .B(n_471), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_448), .B(n_471), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_442), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_442), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_448), .B(n_442), .Y(n_510) );
INVxp67_ASAP7_75t_L g511 ( .A(n_442), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_448), .B(n_453), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_448), .Y(n_513) );
AOI31xp33_ASAP7_75t_L g514 ( .A1(n_462), .A2(n_439), .A3(n_465), .B(n_437), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_453), .B(n_465), .Y(n_515) );
INVxp33_ASAP7_75t_L g516 ( .A(n_453), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_442), .B(n_444), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_444), .B(n_463), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_444), .B(n_463), .Y(n_519) );
OAI33xp33_ASAP7_75t_L g520 ( .A1(n_459), .A2(n_460), .A3(n_456), .B1(n_469), .B2(n_461), .B3(n_447), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_444), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_444), .B(n_463), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_444), .B(n_463), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_451), .B(n_455), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_483), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_474), .B(n_455), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_478), .Y(n_527) );
INVx1_ASAP7_75t_SL g528 ( .A(n_503), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_500), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_481), .B(n_455), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_478), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_481), .B(n_455), .Y(n_532) );
NAND2xp33_ASAP7_75t_L g533 ( .A(n_503), .B(n_447), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_479), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_485), .B(n_487), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_479), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_486), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_485), .B(n_455), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_486), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_487), .B(n_451), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_488), .B(n_451), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_483), .Y(n_542) );
NOR3xp33_ASAP7_75t_SL g543 ( .A(n_504), .B(n_520), .C(n_501), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_484), .A2(n_469), .B(n_461), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_488), .B(n_451), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_500), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_475), .B(n_451), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_495), .B(n_447), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_490), .B(n_441), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_490), .B(n_441), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_502), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_483), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_495), .B(n_447), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_494), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_492), .B(n_441), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_502), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_498), .B(n_461), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_475), .B(n_441), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_494), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_480), .B(n_441), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_492), .B(n_441), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_498), .B(n_461), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_508), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_480), .B(n_456), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_489), .B(n_456), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_518), .B(n_456), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_518), .B(n_460), .Y(n_567) );
AND2x4_ASAP7_75t_SL g568 ( .A(n_496), .B(n_506), .Y(n_568) );
AND2x4_ASAP7_75t_L g569 ( .A(n_474), .B(n_460), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_499), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_508), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_522), .B(n_460), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_509), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_499), .B(n_515), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_496), .B(n_469), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_522), .B(n_523), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_509), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_515), .B(n_461), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_521), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_494), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_523), .B(n_469), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_521), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_497), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_510), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_497), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_535), .B(n_482), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_527), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_584), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_533), .A2(n_484), .B1(n_496), .B2(n_476), .Y(n_589) );
OR2x6_ASAP7_75t_L g590 ( .A(n_526), .B(n_496), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_527), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_581), .B(n_477), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_535), .B(n_482), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_576), .B(n_482), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_576), .B(n_482), .Y(n_595) );
INVx3_ASAP7_75t_SL g596 ( .A(n_570), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_528), .B(n_510), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_531), .Y(n_598) );
INVx3_ASAP7_75t_L g599 ( .A(n_568), .Y(n_599) );
OR2x6_ASAP7_75t_L g600 ( .A(n_526), .B(n_493), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_529), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_531), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_534), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_548), .B(n_517), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_581), .B(n_477), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_574), .B(n_519), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_530), .B(n_517), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_530), .B(n_506), .Y(n_608) );
INVxp67_ASAP7_75t_L g609 ( .A(n_546), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_553), .B(n_493), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_563), .B(n_512), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_558), .B(n_519), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_534), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_558), .B(n_511), .Y(n_614) );
AO21x1_ASAP7_75t_L g615 ( .A1(n_544), .A2(n_514), .B(n_516), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_560), .B(n_511), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_560), .B(n_561), .Y(n_617) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_543), .A2(n_476), .B(n_514), .Y(n_618) );
INVx1_ASAP7_75t_SL g619 ( .A(n_565), .Y(n_619) );
INVx1_ASAP7_75t_SL g620 ( .A(n_565), .Y(n_620) );
INVxp67_ASAP7_75t_L g621 ( .A(n_555), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_563), .B(n_512), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_532), .B(n_506), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_575), .A2(n_506), .B1(n_524), .B2(n_491), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_575), .A2(n_524), .B1(n_491), .B2(n_520), .Y(n_625) );
INVx3_ASAP7_75t_L g626 ( .A(n_568), .Y(n_626) );
NOR2xp67_ASAP7_75t_L g627 ( .A(n_526), .B(n_504), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_566), .Y(n_628) );
INVxp67_ASAP7_75t_SL g629 ( .A(n_525), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_532), .B(n_505), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_536), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_571), .B(n_491), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_555), .B(n_513), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_536), .Y(n_634) );
AND2x4_ASAP7_75t_L g635 ( .A(n_568), .B(n_505), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_537), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_537), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_561), .B(n_497), .Y(n_638) );
INVx1_ASAP7_75t_SL g639 ( .A(n_566), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_539), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_615), .B(n_526), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_617), .B(n_547), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_614), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_616), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_587), .Y(n_645) );
INVx1_ASAP7_75t_SL g646 ( .A(n_596), .Y(n_646) );
OR2x2_ASAP7_75t_L g647 ( .A(n_612), .B(n_547), .Y(n_647) );
AND2x4_ASAP7_75t_L g648 ( .A(n_590), .B(n_575), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_601), .B(n_545), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_609), .B(n_562), .Y(n_650) );
AOI222xp33_ASAP7_75t_L g651 ( .A1(n_618), .A2(n_545), .B1(n_541), .B2(n_557), .C1(n_540), .C2(n_575), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_601), .B(n_541), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_591), .Y(n_653) );
AND2x4_ASAP7_75t_L g654 ( .A(n_590), .B(n_569), .Y(n_654) );
INVxp67_ASAP7_75t_L g655 ( .A(n_588), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_609), .B(n_540), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_639), .B(n_549), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_639), .B(n_549), .Y(n_658) );
NOR2xp33_ASAP7_75t_SL g659 ( .A(n_599), .B(n_550), .Y(n_659) );
AND2x4_ASAP7_75t_SL g660 ( .A(n_599), .B(n_550), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_607), .B(n_538), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_592), .B(n_582), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_592), .B(n_582), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_605), .B(n_573), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_633), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_638), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_605), .B(n_573), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_598), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_600), .A2(n_578), .B(n_491), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_619), .B(n_571), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_602), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_600), .A2(n_564), .B1(n_538), .B2(n_579), .Y(n_672) );
INVxp33_ASAP7_75t_L g673 ( .A(n_627), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_619), .B(n_579), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_586), .B(n_572), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_603), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_613), .Y(n_677) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_620), .Y(n_678) );
INVx2_ASAP7_75t_SL g679 ( .A(n_626), .Y(n_679) );
NAND2x1p5_ASAP7_75t_L g680 ( .A(n_654), .B(n_626), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_650), .B(n_621), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_671), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_673), .A2(n_600), .B1(n_589), .B2(n_590), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_671), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_650), .B(n_620), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_662), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_663), .Y(n_687) );
OAI21xp33_ASAP7_75t_L g688 ( .A1(n_673), .A2(n_625), .B(n_624), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_661), .B(n_593), .Y(n_689) );
AOI22xp33_ASAP7_75t_SL g690 ( .A1(n_659), .A2(n_635), .B1(n_610), .B2(n_604), .Y(n_690) );
OR2x2_ASAP7_75t_L g691 ( .A(n_642), .B(n_597), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_641), .A2(n_632), .B1(n_622), .B2(n_611), .C(n_636), .Y(n_692) );
OAI21xp5_ASAP7_75t_L g693 ( .A1(n_641), .A2(n_635), .B(n_632), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_657), .Y(n_694) );
OAI21xp5_ASAP7_75t_L g695 ( .A1(n_646), .A2(n_629), .B(n_577), .Y(n_695) );
AOI22xp5_ASAP7_75t_SL g696 ( .A1(n_672), .A2(n_594), .B1(n_595), .B2(n_628), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_664), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_667), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_643), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_660), .B(n_608), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_644), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_645), .Y(n_702) );
AOI211xp5_ASAP7_75t_L g703 ( .A1(n_669), .A2(n_606), .B(n_623), .C(n_634), .Y(n_703) );
OAI211xp5_ASAP7_75t_SL g704 ( .A1(n_688), .A2(n_651), .B(n_655), .C(n_656), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g705 ( .A1(n_692), .A2(n_655), .B1(n_678), .B2(n_652), .C(n_649), .Y(n_705) );
OAI21xp33_ASAP7_75t_SL g706 ( .A1(n_692), .A2(n_679), .B(n_678), .Y(n_706) );
OAI21xp5_ASAP7_75t_L g707 ( .A1(n_693), .A2(n_654), .B(n_658), .Y(n_707) );
AOI21xp5_ASAP7_75t_SL g708 ( .A1(n_683), .A2(n_654), .B(n_648), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_690), .A2(n_660), .B1(n_648), .B2(n_647), .Y(n_709) );
AOI222xp33_ASAP7_75t_L g710 ( .A1(n_699), .A2(n_677), .B1(n_676), .B2(n_653), .C1(n_668), .C2(n_670), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g711 ( .A1(n_690), .A2(n_674), .B(n_666), .Y(n_711) );
AOI322xp5_ASAP7_75t_L g712 ( .A1(n_681), .A2(n_675), .A3(n_666), .B1(n_665), .B2(n_630), .C1(n_622), .C2(n_611), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_696), .B(n_665), .Y(n_713) );
NAND3xp33_ASAP7_75t_SL g714 ( .A(n_703), .B(n_564), .C(n_577), .Y(n_714) );
O2A1O1Ixp33_ASAP7_75t_L g715 ( .A1(n_695), .A2(n_640), .B(n_637), .C(n_631), .Y(n_715) );
NOR2x1_ASAP7_75t_L g716 ( .A(n_700), .B(n_556), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_680), .A2(n_569), .B(n_572), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_680), .A2(n_569), .B(n_567), .Y(n_718) );
OAI321xp33_ASAP7_75t_L g719 ( .A1(n_704), .A2(n_685), .A3(n_701), .B1(n_698), .B2(n_697), .C(n_686), .Y(n_719) );
NAND3xp33_ASAP7_75t_L g720 ( .A(n_706), .B(n_702), .C(n_687), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_708), .A2(n_694), .B1(n_684), .B2(n_682), .C(n_689), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_715), .Y(n_722) );
INVxp67_ASAP7_75t_L g723 ( .A(n_710), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_709), .B(n_691), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_708), .A2(n_694), .B1(n_689), .B2(n_569), .C(n_556), .Y(n_725) );
OAI221xp5_ASAP7_75t_L g726 ( .A1(n_705), .A2(n_551), .B1(n_539), .B2(n_567), .C(n_585), .Y(n_726) );
OAI22xp33_ASAP7_75t_L g727 ( .A1(n_714), .A2(n_551), .B1(n_585), .B2(n_552), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_722), .Y(n_728) );
AOI221xp5_ASAP7_75t_L g729 ( .A1(n_723), .A2(n_711), .B1(n_713), .B2(n_707), .C(n_717), .Y(n_729) );
NAND5xp2_ASAP7_75t_L g730 ( .A(n_719), .B(n_712), .C(n_718), .D(n_716), .E(n_507), .Y(n_730) );
OAI221xp5_ASAP7_75t_L g731 ( .A1(n_721), .A2(n_542), .B1(n_583), .B2(n_580), .C(n_559), .Y(n_731) );
NAND5xp2_ASAP7_75t_L g732 ( .A(n_725), .B(n_507), .C(n_454), .D(n_438), .E(n_542), .Y(n_732) );
AOI211xp5_ASAP7_75t_L g733 ( .A1(n_730), .A2(n_724), .B(n_727), .C(n_720), .Y(n_733) );
NAND3xp33_ASAP7_75t_SL g734 ( .A(n_729), .B(n_726), .C(n_552), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_728), .B(n_552), .Y(n_735) );
INVx1_ASAP7_75t_SL g736 ( .A(n_735), .Y(n_736) );
XNOR2xp5_ASAP7_75t_L g737 ( .A(n_733), .B(n_731), .Y(n_737) );
OAI22xp5_ASAP7_75t_SL g738 ( .A1(n_737), .A2(n_734), .B1(n_732), .B2(n_454), .Y(n_738) );
OAI21xp5_ASAP7_75t_L g739 ( .A1(n_736), .A2(n_454), .B(n_542), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_738), .A2(n_554), .B1(n_583), .B2(n_580), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_740), .A2(n_739), .B1(n_554), .B2(n_559), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_741), .B(n_438), .Y(n_742) );
AOI22x1_ASAP7_75t_L g743 ( .A1(n_742), .A2(n_554), .B1(n_583), .B2(n_580), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_743), .A2(n_525), .B1(n_559), .B2(n_585), .Y(n_744) );
endmodule