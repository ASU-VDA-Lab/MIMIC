module real_jpeg_25860_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_11;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_3),
.A2(n_24),
.B1(n_27),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_3),
.A2(n_33),
.B1(n_40),
.B2(n_42),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_3),
.A2(n_18),
.B(n_27),
.C(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_3),
.B(n_16),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_3),
.A2(n_19),
.B1(n_20),
.B2(n_33),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_3),
.B(n_39),
.C(n_40),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_3),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_3),
.B(n_37),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_4),
.A2(n_19),
.B1(n_20),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_4),
.A2(n_40),
.B1(n_42),
.B2(n_47),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_6),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_23)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_6),
.A2(n_19),
.B1(n_20),
.B2(n_26),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_6),
.A2(n_26),
.B1(n_40),
.B2(n_42),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_8),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_8),
.B(n_71),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_74),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_72),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_58),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_12),
.B(n_58),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_48),
.Y(n_12)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_34),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_28),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_23),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_17)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_18),
.A2(n_22),
.B1(n_24),
.B2(n_27),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_19),
.A2(n_20),
.B1(n_38),
.B2(n_39),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g56 ( 
.A1(n_19),
.A2(n_22),
.B(n_33),
.Y(n_56)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_20),
.B(n_82),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_43),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_35),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_46),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_40),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_40),
.B(n_98),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_44),
.B(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_55),
.B2(n_57),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_53),
.B(n_54),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_70),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_51),
.B(n_54),
.Y(n_102)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_55),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.C(n_64),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_63),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_65),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_106),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_87),
.B(n_110),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_83),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_76),
.B(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_80),
.B1(n_81),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_95),
.B(n_109),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_103),
.B(n_108),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_104),
.B(n_105),
.Y(n_108)
);


endmodule