module fake_aes_2783_n_16 (n_1, n_2, n_0, n_16);
input n_1;
input n_2;
input n_0;
output n_16;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
NAND2xp5_ASAP7_75t_L g5 ( .A(n_4), .B(n_0), .Y(n_5) );
OAI22xp5_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_6) );
INVx2_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_6), .B(n_3), .Y(n_8) );
AND2x2_ASAP7_75t_L g9 ( .A(n_7), .B(n_0), .Y(n_9) );
INVx1_ASAP7_75t_SL g10 ( .A(n_8), .Y(n_10) );
AOI21xp5_ASAP7_75t_L g11 ( .A1(n_9), .A2(n_0), .B(n_1), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_9), .B(n_1), .Y(n_12) );
NOR2x1p5_ASAP7_75t_L g13 ( .A(n_12), .B(n_10), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_11), .Y(n_14) );
OR2x2_ASAP7_75t_L g15 ( .A(n_13), .B(n_10), .Y(n_15) );
OAI22xp5_ASAP7_75t_SL g16 ( .A1(n_15), .A2(n_2), .B1(n_14), .B2(n_12), .Y(n_16) );
endmodule