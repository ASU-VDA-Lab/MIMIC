module fake_jpeg_4455_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_34),
.B(n_37),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_43),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_41),
.B(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_46),
.Y(n_86)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_52),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_33),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_39),
.B1(n_16),
.B2(n_43),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_56),
.B1(n_68),
.B2(n_70),
.Y(n_75)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_16),
.B1(n_26),
.B2(n_28),
.Y(n_56)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_31),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_66),
.Y(n_97)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_16),
.B1(n_18),
.B2(n_26),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_18),
.B1(n_26),
.B2(n_28),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_20),
.B(n_24),
.C(n_30),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_40),
.A2(n_18),
.B1(n_26),
.B2(n_28),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_42),
.A2(n_28),
.B1(n_24),
.B2(n_30),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_27),
.B(n_19),
.Y(n_80)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_90),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_48),
.B(n_42),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_91),
.C(n_56),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_80),
.A2(n_88),
.B(n_66),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_27),
.B1(n_19),
.B2(n_23),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_83),
.A2(n_64),
.B1(n_62),
.B2(n_17),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_42),
.C(n_25),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_25),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_42),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_44),
.B(n_40),
.C(n_29),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_60),
.A2(n_17),
.B1(n_32),
.B2(n_20),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_61),
.B(n_54),
.C(n_49),
.Y(n_111)
);

MAJx2_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_69),
.C(n_50),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_99),
.C(n_118),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_45),
.B(n_52),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_105),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_72),
.B(n_50),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_114),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_92),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_107),
.A2(n_111),
.B1(n_32),
.B2(n_19),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_91),
.A2(n_70),
.B1(n_71),
.B2(n_57),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_100),
.B1(n_99),
.B2(n_118),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_20),
.Y(n_110)
);

NOR2x1_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_119),
.Y(n_137)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_115),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_86),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_122),
.B1(n_74),
.B2(n_88),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_121),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_79),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_79),
.A2(n_51),
.B(n_59),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_124),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_92),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_123),
.B(n_93),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_84),
.A2(n_67),
.B(n_63),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_54),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_127),
.A2(n_148),
.B1(n_125),
.B2(n_124),
.Y(n_167)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_143),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_107),
.Y(n_131)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_86),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_135),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_75),
.B1(n_88),
.B2(n_84),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_136),
.B1(n_145),
.B2(n_117),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_74),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_96),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_150),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_140),
.B(n_146),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_141),
.B(n_151),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_75),
.B1(n_93),
.B2(n_57),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_144),
.B1(n_149),
.B2(n_101),
.Y(n_173)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_65),
.B1(n_58),
.B2(n_90),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_65),
.B1(n_58),
.B2(n_78),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_100),
.A2(n_55),
.B1(n_77),
.B2(n_65),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_98),
.A2(n_76),
.B1(n_73),
.B2(n_44),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_105),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_87),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_118),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_116),
.B(n_120),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_155),
.A2(n_163),
.B(n_178),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_156),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_118),
.C(n_98),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_166),
.C(n_168),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_144),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_161),
.Y(n_184)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_137),
.A2(n_115),
.B1(n_111),
.B2(n_119),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_148),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_110),
.B1(n_102),
.B2(n_119),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_165),
.A2(n_170),
.B1(n_149),
.B2(n_141),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_127),
.B(n_111),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_173),
.B1(n_145),
.B2(n_142),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_126),
.C(n_152),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_171),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_110),
.B1(n_121),
.B2(n_76),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

XNOR2x1_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_87),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_172),
.B(n_179),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_139),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_175),
.Y(n_208)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_126),
.A2(n_104),
.B(n_101),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_SL g179 ( 
.A1(n_138),
.A2(n_104),
.B(n_32),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_128),
.A2(n_131),
.B(n_140),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_151),
.B(n_150),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_172),
.A2(n_143),
.B1(n_130),
.B2(n_129),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_183),
.A2(n_187),
.B1(n_197),
.B2(n_203),
.Y(n_231)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_189),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_186),
.A2(n_29),
.B1(n_25),
.B2(n_81),
.Y(n_222)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_163),
.B(n_129),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_198),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_204),
.C(n_157),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_180),
.Y(n_211)
);

OAI32xp33_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_23),
.A3(n_27),
.B1(n_31),
.B2(n_44),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_195),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_73),
.Y(n_196)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_173),
.A2(n_108),
.B1(n_24),
.B2(n_30),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_199),
.A2(n_200),
.B(n_201),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_167),
.A2(n_108),
.B1(n_23),
.B2(n_40),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_87),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_156),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_206),
.B(n_203),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_213),
.C(n_219),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_187),
.A2(n_165),
.B1(n_154),
.B2(n_174),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_210),
.A2(n_212),
.B1(n_214),
.B2(n_221),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_211),
.B(n_217),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_154),
.B1(n_171),
.B2(n_155),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_166),
.C(n_164),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_201),
.A2(n_169),
.B1(n_176),
.B2(n_161),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_158),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_158),
.C(n_176),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_158),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_224),
.C(n_225),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_81),
.B1(n_89),
.B2(n_87),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_222),
.A2(n_208),
.B1(n_205),
.B2(n_184),
.Y(n_240)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_191),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_82),
.C(n_89),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_185),
.C(n_194),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_229),
.C(n_233),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_82),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_190),
.A2(n_197),
.B1(n_200),
.B2(n_189),
.Y(n_232)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_182),
.B(n_89),
.C(n_78),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_230),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_253),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_186),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_236),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_227),
.B(n_196),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_199),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_237),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_222),
.B1(n_227),
.B2(n_207),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_238),
.B(n_251),
.Y(n_258)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_207),
.Y(n_242)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_224),
.B(n_183),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_247),
.C(n_0),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_216),
.A2(n_207),
.B1(n_195),
.B2(n_78),
.Y(n_246)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_209),
.B(n_25),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_215),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_249),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_226),
.A2(n_14),
.B1(n_13),
.B2(n_29),
.Y(n_250)
);

AO21x1_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_0),
.B(n_1),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_215),
.A2(n_13),
.B1(n_1),
.B2(n_2),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_218),
.B(n_0),
.Y(n_254)
);

AOI221xp5_ASAP7_75t_L g259 ( 
.A1(n_254),
.A2(n_231),
.B1(n_229),
.B2(n_225),
.C(n_3),
.Y(n_259)
);

FAx1_ASAP7_75t_SL g256 ( 
.A(n_236),
.B(n_211),
.CI(n_220),
.CON(n_256),
.SN(n_256)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_266),
.Y(n_278)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_245),
.A2(n_226),
.B1(n_219),
.B2(n_231),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_263),
.B1(n_4),
.B2(n_5),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_245),
.A2(n_217),
.B1(n_1),
.B2(n_2),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_8),
.Y(n_285)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_234),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_9),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_248),
.A2(n_3),
.B(n_4),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_269),
.A2(n_6),
.B(n_7),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_255),
.C(n_252),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_273),
.C(n_12),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_3),
.C(n_4),
.Y(n_273)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_239),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_274),
.B(n_250),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_271),
.A2(n_243),
.B(n_246),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_275),
.A2(n_277),
.B(n_281),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_261),
.A2(n_244),
.B1(n_235),
.B2(n_255),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_276),
.A2(n_282),
.B1(n_284),
.B2(n_287),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_244),
.B(n_252),
.Y(n_277)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_247),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_272),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_271),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_283),
.A2(n_286),
.B(n_290),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_260),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_288),
.C(n_273),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_10),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_10),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_299),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_270),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_292),
.A2(n_297),
.B(n_303),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_264),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_295),
.B(n_301),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_289),
.B(n_265),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_298),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_274),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_257),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_277),
.A2(n_258),
.B(n_262),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_267),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_302),
.B(n_10),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_268),
.C(n_262),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_294),
.A2(n_265),
.B1(n_287),
.B2(n_281),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_307),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_294),
.A2(n_275),
.B1(n_256),
.B2(n_285),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_266),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_291),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_303),
.A2(n_269),
.B(n_256),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_11),
.B(n_12),
.Y(n_323)
);

A2O1A1Ixp33_ASAP7_75t_SL g312 ( 
.A1(n_304),
.A2(n_266),
.B(n_11),
.C(n_12),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_312),
.A2(n_314),
.B(n_11),
.Y(n_321)
);

INVx11_ASAP7_75t_L g313 ( 
.A(n_297),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_292),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_300),
.Y(n_316)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_316),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_320),
.C(n_322),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_321),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_305),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_293),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_314),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_317),
.Y(n_324)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_324),
.Y(n_330)
);

MAJx2_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_309),
.C(n_312),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_329),
.B(n_328),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_331),
.A2(n_318),
.B(n_326),
.Y(n_332)
);

O2A1O1Ixp33_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_330),
.B(n_325),
.C(n_312),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_11),
.Y(n_334)
);


endmodule