module fake_jpeg_24043_n_333 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_4),
.B(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_30),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_43),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_51),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_1),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_48),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx2_ASAP7_75t_R g48 ( 
.A(n_25),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_1),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_36),
.B1(n_18),
.B2(n_31),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_54),
.A2(n_61),
.B1(n_83),
.B2(n_38),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_36),
.B1(n_31),
.B2(n_29),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_62),
.A2(n_65),
.B1(n_67),
.B2(n_73),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_48),
.A2(n_36),
.B1(n_31),
.B2(n_18),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_68),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_36),
.B1(n_18),
.B2(n_20),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_70),
.B(n_74),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_33),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_71),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_17),
.B1(n_26),
.B2(n_20),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_72),
.A2(n_28),
.B1(n_22),
.B2(n_21),
.Y(n_103)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_34),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_75),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_34),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_76),
.Y(n_115)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_78),
.Y(n_86)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_29),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_29),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_46),
.A2(n_17),
.B1(n_38),
.B2(n_35),
.Y(n_83)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_27),
.Y(n_102)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_56),
.B(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_101),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_46),
.B1(n_17),
.B2(n_20),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_90),
.A2(n_95),
.B1(n_97),
.B2(n_112),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_92),
.A2(n_120),
.B1(n_66),
.B2(n_53),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_64),
.A2(n_26),
.B1(n_35),
.B2(n_38),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_64),
.A2(n_26),
.B1(n_35),
.B2(n_47),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_45),
.C(n_50),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_108),
.C(n_110),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_32),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_102),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g154 ( 
.A1(n_103),
.A2(n_37),
.B1(n_23),
.B2(n_21),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_52),
.B(n_42),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_107),
.Y(n_135)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_113),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_32),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_50),
.C(n_40),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_32),
.C(n_27),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_69),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_28),
.B1(n_22),
.B2(n_23),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_28),
.Y(n_114)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_82),
.B(n_22),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_116),
.B(n_2),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

OR2x2_ASAP7_75t_SL g118 ( 
.A(n_82),
.B(n_27),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_118),
.A2(n_21),
.B(n_19),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_58),
.A2(n_37),
.B1(n_23),
.B2(n_21),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_60),
.B(n_27),
.Y(n_121)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_124),
.A2(n_146),
.B1(n_106),
.B2(n_153),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_77),
.C(n_68),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_126),
.B(n_119),
.C(n_99),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_1),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_132),
.B(n_147),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_85),
.CI(n_70),
.CON(n_133),
.SN(n_133)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_133),
.B(n_143),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_89),
.B(n_32),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_140),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_96),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_138),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_96),
.B(n_80),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_59),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_95),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_148),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_80),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_145),
.Y(n_163)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_92),
.A2(n_78),
.B1(n_74),
.B2(n_73),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_2),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_37),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_151),
.Y(n_164)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_155),
.Y(n_168)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_153),
.B(n_11),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_154),
.A2(n_93),
.B1(n_62),
.B2(n_122),
.Y(n_160)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

FAx1_ASAP7_75t_SL g156 ( 
.A(n_110),
.B(n_37),
.CI(n_23),
.CON(n_156),
.SN(n_156)
);

XOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_156),
.B(n_157),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_19),
.Y(n_158)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_160),
.A2(n_152),
.B1(n_151),
.B2(n_155),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_121),
.B(n_118),
.C(n_91),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_161),
.A2(n_12),
.B(n_5),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_144),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_162),
.Y(n_206)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_180),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_148),
.A2(n_124),
.B1(n_146),
.B2(n_125),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_176),
.B1(n_186),
.B2(n_187),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_130),
.A2(n_122),
.B1(n_88),
.B2(n_104),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_171),
.A2(n_154),
.B(n_19),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_88),
.B1(n_102),
.B2(n_87),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_172),
.A2(n_177),
.B1(n_139),
.B2(n_156),
.Y(n_193)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_174),
.B(n_178),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_125),
.B1(n_126),
.B2(n_141),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_179),
.B(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_138),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_147),
.C(n_123),
.Y(n_200)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_135),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_184),
.B(n_185),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_131),
.B(n_109),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_134),
.A2(n_122),
.B1(n_116),
.B2(n_109),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_134),
.A2(n_94),
.B1(n_115),
.B2(n_19),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_137),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_188),
.Y(n_219)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_190),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_193),
.A2(n_195),
.B1(n_212),
.B2(n_161),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_173),
.A2(n_156),
.B1(n_133),
.B2(n_139),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_133),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_200),
.Y(n_236)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_221),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_184),
.Y(n_202)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_203),
.A2(n_207),
.B1(n_209),
.B2(n_211),
.Y(n_247)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_204),
.B(n_217),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_170),
.A2(n_154),
.B1(n_123),
.B2(n_147),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_132),
.C(n_98),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_183),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_173),
.A2(n_154),
.B1(n_132),
.B2(n_131),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_190),
.A2(n_98),
.B1(n_3),
.B2(n_4),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_2),
.B(n_3),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_216),
.B(n_159),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_176),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_214),
.A2(n_166),
.B1(n_167),
.B2(n_178),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_183),
.B(n_166),
.C(n_12),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_180),
.A2(n_4),
.B(n_6),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_169),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_222),
.B(n_162),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_219),
.B(n_188),
.Y(n_224)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_224),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_226),
.B(n_195),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_221),
.A2(n_169),
.B1(n_192),
.B2(n_189),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_227),
.A2(n_214),
.B1(n_218),
.B2(n_183),
.Y(n_267)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_234),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_216),
.B(n_215),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_200),
.C(n_207),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_205),
.A2(n_192),
.B1(n_172),
.B2(n_160),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_232),
.A2(n_243),
.B1(n_212),
.B2(n_187),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_167),
.Y(n_233)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_206),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_238),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_240),
.A2(n_242),
.B1(n_244),
.B2(n_246),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_206),
.Y(n_241)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_241),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_223),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_199),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_213),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_210),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_248),
.A2(n_217),
.B1(n_204),
.B2(n_179),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_251),
.Y(n_283)
);

XNOR2x1_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_196),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_250),
.B(n_253),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_193),
.Y(n_251)
);

XNOR2x1_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_208),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_258),
.C(n_259),
.Y(n_276)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_257),
.B(n_267),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_228),
.C(n_225),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_247),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_264),
.A2(n_266),
.B1(n_239),
.B2(n_227),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_232),
.A2(n_205),
.B1(n_211),
.B2(n_222),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_265),
.B(n_198),
.Y(n_269)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_279),
.B1(n_273),
.B2(n_274),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_260),
.B(n_268),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_271),
.A2(n_277),
.B(n_229),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_225),
.B1(n_243),
.B2(n_245),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_272),
.A2(n_285),
.B1(n_264),
.B2(n_240),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g275 ( 
.A(n_262),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_275),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_260),
.A2(n_234),
.B(n_241),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_252),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_279),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_233),
.C(n_248),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_282),
.C(n_249),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_244),
.C(n_235),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_231),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_286),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_267),
.A2(n_245),
.B1(n_237),
.B2(n_224),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_242),
.Y(n_286)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_290),
.B(n_271),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_272),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_293),
.C(n_296),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_250),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_257),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_294),
.A2(n_295),
.B(n_289),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_259),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_251),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_194),
.C(n_197),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_297),
.A2(n_6),
.B(n_14),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_285),
.A2(n_194),
.B1(n_198),
.B2(n_13),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_282),
.B1(n_276),
.B2(n_14),
.Y(n_304)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_301),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_307),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_304),
.A2(n_291),
.B1(n_288),
.B2(n_302),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_298),
.B(n_276),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_307),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_283),
.B(n_7),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_306),
.A2(n_287),
.B(n_300),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_283),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_308),
.A2(n_287),
.B(n_294),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_310),
.A2(n_288),
.B(n_290),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_311),
.A2(n_315),
.B(n_316),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_304),
.B(n_297),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_317),
.B(n_318),
.Y(n_323)
);

NAND3xp33_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_314),
.C(n_306),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_319),
.A2(n_311),
.B(n_300),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_309),
.C(n_303),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_296),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_309),
.B(n_318),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_325),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_326),
.Y(n_327)
);

OAI21x1_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_320),
.B(n_321),
.Y(n_329)
);

O2A1O1Ixp33_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_328),
.B(n_293),
.C(n_16),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_15),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_15),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_15),
.B(n_16),
.Y(n_333)
);


endmodule