module fake_netlist_6_2012_n_1724 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1724);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1724;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g156 ( 
.A(n_68),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_34),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_106),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_25),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_38),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_35),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_0),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_127),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_77),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_7),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_90),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_43),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_85),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_11),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_104),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_145),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_11),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_46),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_110),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_38),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_89),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_50),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_84),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_131),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_57),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_17),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_91),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_142),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_54),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_56),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_75),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_88),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_155),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_116),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_54),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_4),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_32),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_71),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_78),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_50),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_136),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_14),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_69),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_20),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_64),
.Y(n_209)
);

BUFx2_ASAP7_75t_SL g210 ( 
.A(n_67),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_31),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_39),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_108),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_95),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_105),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_72),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_129),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_5),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_1),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_6),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_134),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_97),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_152),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_94),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_39),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_34),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_22),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_119),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_30),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_125),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_17),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_93),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_126),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_62),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_74),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_28),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_121),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_35),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_9),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_137),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_16),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_10),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_12),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_41),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_132),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_23),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_47),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_55),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_128),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_102),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_22),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_2),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_49),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_70),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_41),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_79),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_57),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_49),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_15),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_14),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_5),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_139),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_151),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_56),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_31),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_13),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_26),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_47),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_59),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_33),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_122),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_138),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_81),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_1),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_23),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_120),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_0),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_92),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_52),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_63),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_135),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_103),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_141),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_12),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_4),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_148),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_98),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_6),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_33),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_111),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_118),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_55),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_80),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_133),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_28),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_76),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_20),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_40),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_7),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_48),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_10),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_29),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_140),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_18),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_43),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_9),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_2),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_150),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_44),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_163),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_299),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_159),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_215),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_241),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_241),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_241),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_196),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_241),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_168),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_169),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_272),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_R g322 ( 
.A(n_308),
.B(n_147),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_193),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_241),
.Y(n_324)
);

BUFx2_ASAP7_75t_SL g325 ( 
.A(n_162),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_172),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_156),
.B(n_3),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_176),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_299),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_241),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_160),
.B(n_3),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_177),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_218),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_181),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_218),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_193),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_156),
.B(n_8),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_202),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_183),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_202),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_295),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_162),
.B(n_8),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_228),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_236),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_162),
.B(n_13),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_186),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_190),
.Y(n_348)
);

INVxp33_ASAP7_75t_SL g349 ( 
.A(n_158),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_204),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_228),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_195),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_236),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_236),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_242),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_242),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_204),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_242),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_160),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_196),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_170),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_157),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_170),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_276),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_179),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_200),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_213),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_214),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_269),
.Y(n_369)
);

NOR2xp67_ASAP7_75t_L g370 ( 
.A(n_179),
.B(n_15),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_197),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_157),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_204),
.B(n_16),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_273),
.B(n_18),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_R g375 ( 
.A(n_276),
.B(n_58),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_216),
.Y(n_376)
);

INVxp33_ASAP7_75t_SL g377 ( 
.A(n_161),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_197),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_222),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_273),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_223),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_230),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_211),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_211),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_165),
.B(n_19),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_370),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_314),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_314),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_315),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_315),
.B(n_273),
.Y(n_390)
);

CKINVDCx8_ASAP7_75t_R g391 ( 
.A(n_341),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_362),
.B(n_189),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_316),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_316),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_318),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_318),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_317),
.B(n_269),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_324),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_324),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_317),
.B(n_165),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_330),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_375),
.B(n_263),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_370),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_330),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_317),
.B(n_171),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_362),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_376),
.Y(n_407)
);

BUFx8_ASAP7_75t_L g408 ( 
.A(n_350),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_372),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_372),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_350),
.B(n_189),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_350),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_345),
.B(n_353),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_357),
.B(n_201),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_357),
.B(n_201),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_333),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_345),
.B(n_171),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_333),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_335),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_335),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_353),
.B(n_174),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_340),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_340),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_357),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_380),
.Y(n_425)
);

OA21x2_ASAP7_75t_L g426 ( 
.A1(n_342),
.A2(n_219),
.B(n_212),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_380),
.Y(n_427)
);

INVx6_ASAP7_75t_L g428 ( 
.A(n_331),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_341),
.B(n_263),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_354),
.B(n_174),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_380),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_327),
.B(n_245),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_354),
.B(n_180),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_342),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_323),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_359),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_355),
.B(n_180),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_355),
.B(n_245),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_337),
.B(n_194),
.Y(n_439)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_331),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_311),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_359),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_356),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_363),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_363),
.Y(n_445)
);

OAI21x1_ASAP7_75t_L g446 ( 
.A1(n_343),
.A2(n_206),
.B(n_194),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_SL g447 ( 
.A1(n_385),
.A2(n_307),
.B1(n_203),
.B2(n_226),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_365),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_365),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_371),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_371),
.Y(n_451)
);

AND3x1_ASAP7_75t_L g452 ( 
.A(n_346),
.B(n_374),
.C(n_373),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_378),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_378),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_349),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_440),
.B(n_312),
.Y(n_456)
);

OR2x6_ASAP7_75t_L g457 ( 
.A(n_429),
.B(n_325),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_408),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_412),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_425),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_425),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_452),
.A2(n_382),
.B1(n_379),
.B2(n_344),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_440),
.B(n_319),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_440),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_425),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_428),
.A2(n_344),
.B1(n_310),
.B2(n_329),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_425),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_402),
.B(n_320),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_402),
.B(n_326),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_407),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_443),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_425),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_426),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_426),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_L g475 ( 
.A1(n_440),
.A2(n_360),
.B1(n_369),
.B2(n_325),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_425),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_440),
.B(n_328),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_407),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_440),
.B(n_332),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_435),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_426),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_426),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_391),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_439),
.A2(n_275),
.B1(n_247),
.B2(n_246),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_441),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_425),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_428),
.B(n_377),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_426),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_431),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_412),
.Y(n_490)
);

NAND2xp33_ASAP7_75t_L g491 ( 
.A(n_439),
.B(n_185),
.Y(n_491)
);

INVx4_ASAP7_75t_SL g492 ( 
.A(n_428),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_431),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_426),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_429),
.B(n_334),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_428),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_412),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_431),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_428),
.B(n_339),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_400),
.B(n_356),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_391),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_428),
.B(n_347),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_431),
.Y(n_503)
);

NAND3xp33_ASAP7_75t_L g504 ( 
.A(n_447),
.B(n_352),
.C(n_348),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_428),
.B(n_366),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_428),
.B(n_367),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_386),
.B(n_368),
.Y(n_507)
);

CKINVDCx6p67_ASAP7_75t_R g508 ( 
.A(n_435),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_386),
.B(n_381),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_400),
.B(n_358),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_412),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_441),
.B(n_358),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_386),
.B(n_361),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_431),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_403),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_426),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_431),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_403),
.B(n_278),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_426),
.Y(n_519)
);

NAND3xp33_ASAP7_75t_SL g520 ( 
.A(n_447),
.B(n_338),
.C(n_336),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_431),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_400),
.B(n_206),
.Y(n_522)
);

OR2x6_ASAP7_75t_L g523 ( 
.A(n_439),
.B(n_210),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_403),
.B(n_322),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_412),
.Y(n_525)
);

BUFx10_ASAP7_75t_L g526 ( 
.A(n_390),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_443),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_400),
.B(n_232),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_412),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_405),
.B(n_233),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_405),
.B(n_234),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_412),
.Y(n_532)
);

INVx1_ASAP7_75t_SL g533 ( 
.A(n_435),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_387),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_387),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_432),
.B(n_351),
.Y(n_536)
);

NAND3xp33_ASAP7_75t_L g537 ( 
.A(n_447),
.B(n_166),
.C(n_164),
.Y(n_537)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_432),
.B(n_210),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_432),
.A2(n_212),
.B1(n_264),
.B2(n_265),
.Y(n_539)
);

OR2x6_ASAP7_75t_L g540 ( 
.A(n_446),
.B(n_219),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_412),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_387),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_405),
.A2(n_298),
.B1(n_264),
.B2(n_265),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_391),
.B(n_364),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_443),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_405),
.B(n_235),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_412),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_412),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_413),
.B(n_383),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_443),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_452),
.A2(n_321),
.B1(n_313),
.B2(n_274),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_389),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_397),
.B(n_237),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_443),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_413),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_391),
.B(n_263),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_413),
.Y(n_557)
);

OR2x6_ASAP7_75t_L g558 ( 
.A(n_446),
.B(n_238),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_397),
.B(n_208),
.Y(n_559)
);

INVx1_ASAP7_75t_SL g560 ( 
.A(n_435),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_413),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_436),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_389),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_397),
.B(n_167),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_389),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_393),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_397),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_436),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_393),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_424),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_390),
.B(n_249),
.Y(n_571)
);

NAND3xp33_ASAP7_75t_L g572 ( 
.A(n_452),
.B(n_227),
.C(n_309),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_436),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_417),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_393),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_417),
.B(n_383),
.Y(n_576)
);

OAI22xp33_ASAP7_75t_L g577 ( 
.A1(n_442),
.A2(n_270),
.B1(n_279),
.B2(n_259),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g578 ( 
.A(n_442),
.B(n_263),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_390),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_399),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_399),
.Y(n_581)
);

AND2x6_ASAP7_75t_L g582 ( 
.A(n_417),
.B(n_185),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_417),
.B(n_384),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_399),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_SL g585 ( 
.A1(n_421),
.A2(n_248),
.B1(n_184),
.B2(n_243),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_401),
.Y(n_586)
);

INVx6_ASAP7_75t_L g587 ( 
.A(n_408),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_390),
.B(n_250),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_421),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_421),
.B(n_384),
.Y(n_590)
);

INVx1_ASAP7_75t_SL g591 ( 
.A(n_421),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_438),
.A2(n_257),
.B1(n_238),
.B2(n_298),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_390),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_438),
.A2(n_257),
.B1(n_246),
.B2(n_247),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_430),
.B(n_433),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_424),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_442),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_430),
.A2(n_296),
.B1(n_294),
.B2(n_293),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_430),
.B(n_208),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_430),
.Y(n_600)
);

INVx5_ASAP7_75t_L g601 ( 
.A(n_424),
.Y(n_601)
);

NAND3xp33_ASAP7_75t_L g602 ( 
.A(n_433),
.B(n_199),
.C(n_305),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_579),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_593),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_455),
.B(n_433),
.Y(n_605)
);

OR2x6_ASAP7_75t_L g606 ( 
.A(n_457),
.B(n_446),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_534),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_487),
.A2(n_433),
.B1(n_437),
.B2(n_438),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_589),
.B(n_437),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_536),
.B(n_437),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_534),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_555),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_535),
.Y(n_613)
);

O2A1O1Ixp33_ASAP7_75t_L g614 ( 
.A1(n_473),
.A2(n_411),
.B(n_414),
.C(n_415),
.Y(n_614)
);

O2A1O1Ixp5_ASAP7_75t_L g615 ( 
.A1(n_473),
.A2(n_415),
.B(n_414),
.C(n_411),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_535),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_600),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_591),
.B(n_437),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_555),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_557),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_600),
.B(n_438),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_557),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_464),
.A2(n_209),
.B1(n_217),
.B2(n_221),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_512),
.Y(n_624)
);

O2A1O1Ixp33_ASAP7_75t_L g625 ( 
.A1(n_474),
.A2(n_411),
.B(n_414),
.C(n_415),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_474),
.A2(n_446),
.B1(n_438),
.B2(n_284),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_595),
.B(n_438),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_464),
.B(n_408),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_515),
.B(n_173),
.Y(n_629)
);

INVxp67_ASAP7_75t_SL g630 ( 
.A(n_471),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_595),
.B(n_438),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_542),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_561),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_507),
.B(n_175),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_561),
.B(n_445),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_549),
.Y(n_636)
);

INVxp67_ASAP7_75t_SL g637 ( 
.A(n_471),
.Y(n_637)
);

NOR3xp33_ASAP7_75t_L g638 ( 
.A(n_520),
.B(n_253),
.C(n_251),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_509),
.B(n_178),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_574),
.B(n_408),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_513),
.B(n_182),
.Y(n_641)
);

AND2x6_ASAP7_75t_L g642 ( 
.A(n_481),
.B(n_209),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_513),
.B(n_187),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_574),
.B(n_408),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_549),
.Y(n_645)
);

NAND3xp33_ASAP7_75t_L g646 ( 
.A(n_537),
.B(n_572),
.C(n_564),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_456),
.B(n_408),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_481),
.A2(n_275),
.B1(n_268),
.B2(n_288),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_463),
.B(n_408),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_512),
.B(n_485),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_477),
.B(n_185),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_567),
.B(n_254),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_567),
.B(n_188),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g654 ( 
.A(n_518),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_479),
.B(n_444),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_496),
.B(n_185),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_576),
.B(n_444),
.Y(n_657)
);

O2A1O1Ixp33_ASAP7_75t_L g658 ( 
.A1(n_482),
.A2(n_392),
.B(n_445),
.C(n_451),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_480),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_576),
.B(n_590),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_499),
.A2(n_392),
.B(n_409),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_527),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_590),
.B(n_444),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_524),
.B(n_191),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_562),
.B(n_444),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_562),
.B(n_444),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_496),
.B(n_185),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_482),
.A2(n_284),
.B1(n_267),
.B2(n_288),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_542),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_504),
.A2(n_282),
.B1(n_283),
.B2(n_262),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_545),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_L g672 ( 
.A1(n_475),
.A2(n_240),
.B1(n_290),
.B2(n_303),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_502),
.B(n_185),
.Y(n_673)
);

INVxp33_ASAP7_75t_L g674 ( 
.A(n_585),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_568),
.B(n_444),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_533),
.B(n_445),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_560),
.B(n_450),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_545),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_568),
.B(n_444),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_505),
.B(n_291),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_523),
.A2(n_271),
.B1(n_287),
.B2(n_286),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_500),
.B(n_450),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_573),
.B(n_444),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_573),
.B(n_500),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_510),
.B(n_444),
.Y(n_685)
);

INVx8_ASAP7_75t_L g686 ( 
.A(n_457),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_L g687 ( 
.A1(n_488),
.A2(n_516),
.B(n_494),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_466),
.B(n_192),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_523),
.B(n_198),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_552),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_550),
.Y(n_691)
);

AO22x2_ASAP7_75t_L g692 ( 
.A1(n_556),
.A2(n_217),
.B1(n_221),
.B2(n_224),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_583),
.B(n_450),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_510),
.B(n_444),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_523),
.B(n_205),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_597),
.B(n_392),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_470),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_550),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_506),
.B(n_291),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_488),
.B(n_291),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_523),
.B(n_538),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_552),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_554),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_599),
.B(n_494),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_516),
.B(n_291),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_563),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_599),
.B(n_401),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_583),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_563),
.Y(n_709)
);

A2O1A1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_519),
.A2(n_224),
.B(n_240),
.C(n_290),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_519),
.B(n_291),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_522),
.B(n_404),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_526),
.B(n_291),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_538),
.A2(n_457),
.B1(n_530),
.B2(n_546),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_538),
.B(n_207),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_559),
.B(n_404),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_565),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_565),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_566),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_526),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_478),
.Y(n_721)
);

NAND2xp33_ASAP7_75t_L g722 ( 
.A(n_582),
.B(n_256),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_559),
.B(n_404),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_483),
.B(n_231),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_538),
.A2(n_303),
.B1(n_280),
.B2(n_281),
.Y(n_725)
);

NOR3xp33_ASAP7_75t_L g726 ( 
.A(n_495),
.B(n_302),
.C(n_225),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_483),
.B(n_231),
.Y(n_727)
);

BUFx12f_ASAP7_75t_L g728 ( 
.A(n_457),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_528),
.B(n_448),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_553),
.Y(n_730)
);

A2O1A1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_602),
.A2(n_571),
.B(n_588),
.C(n_491),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_SL g732 ( 
.A(n_578),
.B(n_231),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_492),
.B(n_451),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_531),
.B(n_448),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_566),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_468),
.B(n_220),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_469),
.A2(n_451),
.B1(n_454),
.B2(n_453),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_492),
.B(n_424),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_569),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_598),
.B(n_229),
.Y(n_740)
);

NOR2xp67_ASAP7_75t_L g741 ( 
.A(n_462),
.B(n_416),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_551),
.A2(n_454),
.B1(n_453),
.B2(n_449),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_544),
.B(n_231),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_569),
.B(n_448),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_575),
.Y(n_745)
);

O2A1O1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_540),
.A2(n_267),
.B(n_268),
.C(n_449),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_492),
.B(n_424),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_575),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_580),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_540),
.A2(n_454),
.B1(n_453),
.B2(n_449),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_580),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_581),
.Y(n_752)
);

INVx8_ASAP7_75t_L g753 ( 
.A(n_501),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_540),
.A2(n_454),
.B1(n_453),
.B2(n_449),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_581),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_584),
.B(n_448),
.Y(n_756)
);

BUFx8_ASAP7_75t_L g757 ( 
.A(n_508),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_577),
.B(n_239),
.Y(n_758)
);

AND2x4_ASAP7_75t_SL g759 ( 
.A(n_501),
.B(n_416),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_584),
.B(n_449),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_539),
.B(n_416),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_540),
.B(n_244),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_586),
.Y(n_763)
);

NAND2x1_ASAP7_75t_L g764 ( 
.A(n_587),
.B(n_424),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_492),
.B(n_424),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_558),
.B(n_252),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_558),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_586),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_610),
.B(n_558),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_654),
.B(n_508),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_687),
.A2(n_458),
.B(n_596),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_617),
.Y(n_772)
);

BUFx8_ASAP7_75t_L g773 ( 
.A(n_728),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_617),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_735),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_733),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_610),
.B(n_558),
.Y(n_777)
);

BUFx12f_ASAP7_75t_L g778 ( 
.A(n_757),
.Y(n_778)
);

BUFx10_ASAP7_75t_L g779 ( 
.A(n_653),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_L g780 ( 
.A1(n_704),
.A2(n_497),
.B(n_511),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_729),
.A2(n_570),
.B(n_596),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_648),
.A2(n_484),
.B1(n_594),
.B2(n_592),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_624),
.B(n_641),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_734),
.A2(n_490),
.B(n_570),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_635),
.Y(n_785)
);

A2O1A1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_688),
.A2(n_543),
.B(n_511),
.C(n_525),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_635),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_714),
.B(n_646),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_735),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_650),
.B(n_255),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_605),
.B(n_497),
.Y(n_791)
);

AOI21x1_ASAP7_75t_L g792 ( 
.A1(n_700),
.A2(n_476),
.B(n_472),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_674),
.B(n_258),
.Y(n_793)
);

OAI21xp33_ASAP7_75t_L g794 ( 
.A1(n_758),
.A2(n_300),
.B(n_306),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_745),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_730),
.B(n_497),
.Y(n_796)
);

AOI21xp33_ASAP7_75t_L g797 ( 
.A1(n_688),
.A2(n_292),
.B(n_261),
.Y(n_797)
);

CKINVDCx6p67_ASAP7_75t_R g798 ( 
.A(n_753),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_612),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_697),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_660),
.B(n_459),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_627),
.A2(n_547),
.B(n_541),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_767),
.B(n_529),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_608),
.A2(n_587),
.B1(n_511),
.B2(n_525),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_653),
.B(n_260),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_631),
.A2(n_529),
.B(n_548),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_701),
.A2(n_582),
.B1(n_521),
.B2(n_465),
.Y(n_807)
);

AOI21x1_ASAP7_75t_L g808 ( 
.A1(n_700),
.A2(n_486),
.B(n_461),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_619),
.B(n_525),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_621),
.A2(n_655),
.B(n_696),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_672),
.A2(n_453),
.B(n_454),
.C(n_410),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_708),
.B(n_266),
.Y(n_812)
);

NOR2x2_ASAP7_75t_L g813 ( 
.A(n_606),
.B(n_277),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_661),
.A2(n_529),
.B(n_548),
.Y(n_814)
);

NOR2x1_ASAP7_75t_L g815 ( 
.A(n_676),
.B(n_532),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_620),
.B(n_532),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_622),
.B(n_532),
.Y(n_817)
);

O2A1O1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_623),
.A2(n_410),
.B(n_422),
.C(n_423),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_641),
.B(n_419),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_701),
.A2(n_582),
.B1(n_465),
.B2(n_460),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_762),
.A2(n_489),
.B(n_460),
.C(n_461),
.Y(n_821)
);

OR2x6_ASAP7_75t_L g822 ( 
.A(n_753),
.B(n_686),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_685),
.A2(n_529),
.B(n_541),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_694),
.A2(n_541),
.B(n_547),
.Y(n_824)
);

NOR2x1_ASAP7_75t_L g825 ( 
.A(n_677),
.B(n_467),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_615),
.A2(n_486),
.B(n_472),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_633),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_657),
.A2(n_547),
.B(n_548),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_609),
.B(n_582),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_745),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_751),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_618),
.B(n_582),
.Y(n_832)
);

AOI21x1_ASAP7_75t_L g833 ( 
.A1(n_705),
.A2(n_489),
.B(n_493),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_721),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_663),
.A2(n_547),
.B(n_548),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_682),
.B(n_582),
.Y(n_836)
);

OAI21xp5_ASAP7_75t_L g837 ( 
.A1(n_705),
.A2(n_498),
.B(n_467),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_682),
.B(n_476),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_603),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_643),
.B(n_419),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_643),
.B(n_634),
.Y(n_841)
);

AOI21x1_ASAP7_75t_L g842 ( 
.A1(n_711),
.A2(n_498),
.B(n_493),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_732),
.B(n_548),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_604),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_733),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_724),
.B(n_419),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_753),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_711),
.A2(n_601),
.B(n_503),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_713),
.A2(n_601),
.B(n_503),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_684),
.B(n_514),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_713),
.A2(n_601),
.B(n_514),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_636),
.B(n_517),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_645),
.B(n_517),
.Y(n_853)
);

INVxp67_ASAP7_75t_L g854 ( 
.A(n_659),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_634),
.B(n_521),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_762),
.A2(n_587),
.B1(n_410),
.B2(n_420),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_639),
.B(n_285),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_614),
.A2(n_625),
.B(n_731),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_639),
.B(n_289),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_766),
.A2(n_587),
.B1(n_420),
.B2(n_423),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_766),
.A2(n_420),
.B1(n_422),
.B2(n_423),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_761),
.B(n_693),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_664),
.A2(n_740),
.B1(n_741),
.B2(n_736),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_630),
.A2(n_601),
.B(n_409),
.Y(n_864)
);

AOI21x1_ASAP7_75t_L g865 ( 
.A1(n_651),
.A2(n_409),
.B(n_434),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_751),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_626),
.A2(n_297),
.B1(n_301),
.B2(n_304),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_727),
.B(n_19),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_637),
.A2(n_601),
.B(n_409),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_626),
.A2(n_394),
.B(n_395),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_664),
.B(n_422),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_629),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_648),
.B(n_395),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_740),
.A2(n_434),
.B(n_418),
.C(n_395),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_662),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_712),
.A2(n_406),
.B(n_427),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_658),
.A2(n_395),
.B(n_396),
.Y(n_877)
);

OAI21xp5_ASAP7_75t_L g878 ( 
.A1(n_651),
.A2(n_395),
.B(n_396),
.Y(n_878)
);

OAI21x1_ASAP7_75t_L g879 ( 
.A1(n_764),
.A2(n_394),
.B(n_395),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_671),
.Y(n_880)
);

NAND2xp33_ASAP7_75t_L g881 ( 
.A(n_642),
.B(n_424),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_678),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_668),
.B(n_394),
.Y(n_883)
);

NOR2xp67_ASAP7_75t_L g884 ( 
.A(n_670),
.B(n_82),
.Y(n_884)
);

INVx4_ASAP7_75t_L g885 ( 
.A(n_720),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_716),
.A2(n_406),
.B(n_427),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_723),
.A2(n_406),
.B(n_427),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_668),
.B(n_394),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_759),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_629),
.B(n_21),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_640),
.B(n_427),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_707),
.A2(n_406),
.B(n_427),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_647),
.A2(n_406),
.B(n_427),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_691),
.B(n_394),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_649),
.A2(n_699),
.B(n_680),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_644),
.B(n_427),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_673),
.A2(n_406),
.B(n_427),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_673),
.A2(n_427),
.B(n_396),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_680),
.A2(n_427),
.B(n_396),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_698),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_703),
.B(n_396),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_715),
.B(n_21),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_715),
.B(n_24),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_699),
.A2(n_396),
.B(n_395),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_742),
.B(n_396),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_738),
.A2(n_394),
.B(n_418),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_743),
.B(n_434),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_758),
.B(n_434),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_710),
.A2(n_394),
.B(n_434),
.C(n_418),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_718),
.B(n_418),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_689),
.B(n_695),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_738),
.A2(n_418),
.B(n_398),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_754),
.B(n_398),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_719),
.B(n_398),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_746),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_915)
);

NAND2x1p5_ASAP7_75t_L g916 ( 
.A(n_720),
.B(n_398),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_736),
.B(n_398),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_689),
.B(n_695),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_681),
.A2(n_398),
.B(n_388),
.C(n_30),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_748),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_652),
.B(n_27),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_725),
.B(n_27),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_686),
.B(n_29),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_755),
.B(n_398),
.Y(n_924)
);

NOR2xp67_ASAP7_75t_SL g925 ( 
.A(n_628),
.B(n_747),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_686),
.B(n_32),
.Y(n_926)
);

AOI21x1_ASAP7_75t_L g927 ( 
.A1(n_765),
.A2(n_398),
.B(n_388),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_763),
.B(n_398),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_754),
.B(n_398),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_SL g930 ( 
.A(n_757),
.B(n_388),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_638),
.B(n_36),
.Y(n_931)
);

BUFx12f_ASAP7_75t_L g932 ( 
.A(n_606),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_750),
.A2(n_388),
.B(n_73),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_642),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_607),
.B(n_388),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_642),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_606),
.B(n_36),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_611),
.B(n_613),
.Y(n_938)
);

NOR2xp67_ASAP7_75t_L g939 ( 
.A(n_737),
.B(n_83),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_616),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_628),
.A2(n_388),
.B(n_86),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_632),
.B(n_37),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_692),
.Y(n_943)
);

A2O1A1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_726),
.A2(n_388),
.B(n_40),
.C(n_42),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_669),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_656),
.A2(n_388),
.B(n_87),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_656),
.A2(n_388),
.B(n_66),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_690),
.B(n_768),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_667),
.A2(n_388),
.B(n_99),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_841),
.A2(n_890),
.B1(n_903),
.B2(n_902),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_810),
.A2(n_760),
.B(n_756),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_841),
.B(n_752),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_845),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_819),
.B(n_692),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_857),
.A2(n_749),
.B(n_702),
.C(n_739),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_771),
.A2(n_744),
.B(n_683),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_840),
.B(n_857),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_863),
.A2(n_692),
.B1(n_717),
.B2(n_709),
.Y(n_958)
);

NOR2xp67_ASAP7_75t_L g959 ( 
.A(n_854),
.B(n_667),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_872),
.B(n_706),
.Y(n_960)
);

O2A1O1Ixp5_ASAP7_75t_L g961 ( 
.A1(n_788),
.A2(n_858),
.B(n_890),
.C(n_859),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_800),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_839),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_859),
.B(n_642),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_834),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_L g966 ( 
.A1(n_911),
.A2(n_642),
.B1(n_722),
.B2(n_675),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_875),
.Y(n_967)
);

NAND2x1p5_ASAP7_75t_L g968 ( 
.A(n_845),
.B(n_666),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_862),
.B(n_679),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_882),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_805),
.B(n_665),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_932),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_769),
.A2(n_65),
.B(n_130),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_844),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_845),
.Y(n_975)
);

INVxp67_ASAP7_75t_L g976 ( 
.A(n_846),
.Y(n_976)
);

BUFx12f_ASAP7_75t_L g977 ( 
.A(n_773),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_911),
.A2(n_37),
.B(n_42),
.C(n_44),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_845),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_805),
.B(n_45),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_777),
.A2(n_100),
.B(n_123),
.Y(n_981)
);

OR2x6_ASAP7_75t_L g982 ( 
.A(n_822),
.B(n_61),
.Y(n_982)
);

OAI22x1_ASAP7_75t_L g983 ( 
.A1(n_902),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_778),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_798),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_918),
.A2(n_107),
.B1(n_117),
.B2(n_114),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_903),
.A2(n_101),
.B1(n_113),
.B2(n_109),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_921),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_921),
.A2(n_51),
.B(n_53),
.C(n_60),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_799),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_827),
.Y(n_991)
);

BUFx2_ASAP7_75t_L g992 ( 
.A(n_847),
.Y(n_992)
);

NOR2x1_ASAP7_75t_R g993 ( 
.A(n_889),
.B(n_144),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_788),
.A2(n_895),
.B(n_855),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_931),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_SL g996 ( 
.A(n_770),
.B(n_779),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_793),
.B(n_783),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_779),
.B(n_868),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_793),
.B(n_770),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_908),
.B(n_907),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_775),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_785),
.B(n_787),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_789),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_773),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_868),
.B(n_776),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_933),
.A2(n_797),
.B(n_922),
.C(n_794),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_822),
.Y(n_1007)
);

NOR2xp67_ASAP7_75t_SL g1008 ( 
.A(n_934),
.B(n_936),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_822),
.Y(n_1009)
);

AO32x1_ASAP7_75t_L g1010 ( 
.A1(n_920),
.A2(n_867),
.A3(n_900),
.B1(n_880),
.B2(n_945),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_782),
.B(n_825),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_944),
.A2(n_919),
.B(n_943),
.C(n_922),
.Y(n_1012)
);

INVx1_ASAP7_75t_SL g1013 ( 
.A(n_813),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_791),
.A2(n_780),
.B(n_806),
.Y(n_1014)
);

AND2x2_ASAP7_75t_SL g1015 ( 
.A(n_930),
.B(n_937),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_782),
.A2(n_937),
.B(n_941),
.C(n_790),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_790),
.B(n_774),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_923),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_923),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_943),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_SL g1021 ( 
.A(n_885),
.B(n_926),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_815),
.B(n_772),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_838),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_776),
.Y(n_1024)
);

AOI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_871),
.A2(n_843),
.B1(n_926),
.B2(n_884),
.Y(n_1025)
);

CKINVDCx11_ASAP7_75t_R g1026 ( 
.A(n_934),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_885),
.B(n_812),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_795),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_850),
.B(n_812),
.Y(n_1029)
);

NOR3xp33_ASAP7_75t_SL g1030 ( 
.A(n_915),
.B(n_803),
.C(n_942),
.Y(n_1030)
);

O2A1O1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_786),
.A2(n_818),
.B(n_874),
.C(n_942),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_852),
.B(n_853),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_934),
.B(n_936),
.Y(n_1033)
);

INVxp67_ASAP7_75t_L g1034 ( 
.A(n_852),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_SL g1035 ( 
.A1(n_925),
.A2(n_877),
.B(n_826),
.C(n_860),
.Y(n_1035)
);

INVx3_ASAP7_75t_SL g1036 ( 
.A(n_934),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_830),
.Y(n_1037)
);

NOR3xp33_ASAP7_75t_SL g1038 ( 
.A(n_803),
.B(n_853),
.C(n_836),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_940),
.B(n_861),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_831),
.Y(n_1040)
);

BUFx12f_ASAP7_75t_L g1041 ( 
.A(n_936),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_802),
.A2(n_784),
.B(n_781),
.Y(n_1042)
);

NAND3xp33_ASAP7_75t_SL g1043 ( 
.A(n_856),
.B(n_832),
.C(n_829),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_929),
.A2(n_796),
.B1(n_905),
.B2(n_936),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_940),
.B(n_866),
.Y(n_1045)
);

INVxp67_ASAP7_75t_L g1046 ( 
.A(n_948),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_938),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_916),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_939),
.B(n_807),
.Y(n_1049)
);

AND2x6_ASAP7_75t_L g1050 ( 
.A(n_820),
.B(n_873),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_801),
.A2(n_917),
.B1(n_913),
.B2(n_948),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_801),
.B(n_817),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_809),
.B(n_816),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_SL g1054 ( 
.A1(n_893),
.A2(n_814),
.B(n_909),
.C(n_811),
.Y(n_1054)
);

INVx1_ASAP7_75t_SL g1055 ( 
.A(n_910),
.Y(n_1055)
);

INVx4_ASAP7_75t_L g1056 ( 
.A(n_916),
.Y(n_1056)
);

O2A1O1Ixp5_ASAP7_75t_L g1057 ( 
.A1(n_891),
.A2(n_896),
.B(n_821),
.C(n_804),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_894),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_913),
.B(n_883),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_901),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_878),
.Y(n_1061)
);

CKINVDCx8_ASAP7_75t_R g1062 ( 
.A(n_946),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_914),
.Y(n_1063)
);

AND2x2_ASAP7_75t_SL g1064 ( 
.A(n_881),
.B(n_888),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_891),
.A2(n_896),
.B(n_835),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_870),
.B(n_824),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_924),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_876),
.A2(n_886),
.B(n_887),
.C(n_892),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_928),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_935),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_879),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_837),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_823),
.B(n_828),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_792),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_808),
.B(n_833),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_906),
.A2(n_949),
.B(n_947),
.C(n_904),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_865),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_864),
.B(n_869),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_848),
.A2(n_849),
.B(n_851),
.Y(n_1079)
);

BUFx4f_ASAP7_75t_L g1080 ( 
.A(n_927),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_SL g1081 ( 
.A1(n_898),
.A2(n_899),
.B1(n_897),
.B2(n_912),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_842),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_841),
.A2(n_890),
.B(n_903),
.C(n_902),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_841),
.A2(n_890),
.B1(n_903),
.B2(n_902),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_841),
.A2(n_857),
.B(n_859),
.C(n_863),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_783),
.B(n_536),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_841),
.A2(n_857),
.B(n_859),
.C(n_863),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_810),
.A2(n_771),
.B(n_858),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_841),
.A2(n_890),
.B(n_903),
.C(n_902),
.Y(n_1089)
);

INVx4_ASAP7_75t_L g1090 ( 
.A(n_845),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_841),
.B(n_610),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_SL g1092 ( 
.A1(n_841),
.A2(n_447),
.B1(n_585),
.B2(n_674),
.Y(n_1092)
);

NOR3xp33_ASAP7_75t_SL g1093 ( 
.A(n_841),
.B(n_520),
.C(n_537),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_841),
.A2(n_863),
.B1(n_769),
.B2(n_777),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_841),
.B(n_610),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_841),
.B(n_863),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_841),
.B(n_863),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_875),
.Y(n_1098)
);

AO21x1_ASAP7_75t_L g1099 ( 
.A1(n_1083),
.A2(n_1089),
.B(n_1096),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_950),
.A2(n_1084),
.B1(n_1087),
.B2(n_1085),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_977),
.Y(n_1101)
);

OR2x6_ASAP7_75t_L g1102 ( 
.A(n_982),
.B(n_962),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_965),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_1024),
.Y(n_1104)
);

AOI221xp5_ASAP7_75t_L g1105 ( 
.A1(n_1092),
.A2(n_1083),
.B1(n_1089),
.B2(n_980),
.C(n_999),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1042),
.A2(n_1079),
.B(n_1065),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_997),
.A2(n_1097),
.B1(n_957),
.B2(n_995),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_992),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1088),
.A2(n_994),
.B(n_1000),
.Y(n_1109)
);

INVx4_ASAP7_75t_L g1110 ( 
.A(n_953),
.Y(n_1110)
);

OAI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1091),
.A2(n_1095),
.B1(n_1019),
.B2(n_1018),
.Y(n_1111)
);

AOI31xp67_ASAP7_75t_L g1112 ( 
.A1(n_1078),
.A2(n_966),
.A3(n_1073),
.B(n_964),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_974),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1006),
.A2(n_952),
.B1(n_1029),
.B2(n_1016),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_961),
.A2(n_1094),
.B(n_1011),
.Y(n_1115)
);

NOR4xp25_ASAP7_75t_L g1116 ( 
.A(n_988),
.B(n_978),
.C(n_989),
.D(n_1012),
.Y(n_1116)
);

AND2x6_ASAP7_75t_L g1117 ( 
.A(n_1032),
.B(n_953),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1035),
.A2(n_1066),
.B(n_1014),
.Y(n_1118)
);

AO31x2_ASAP7_75t_L g1119 ( 
.A1(n_1014),
.A2(n_1042),
.A3(n_1068),
.B(n_1075),
.Y(n_1119)
);

AOI31xp67_ASAP7_75t_L g1120 ( 
.A1(n_1049),
.A2(n_1051),
.A3(n_1025),
.B(n_971),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_951),
.A2(n_956),
.B(n_1031),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_961),
.A2(n_1093),
.B(n_1012),
.C(n_1031),
.Y(n_1122)
);

NOR2xp67_ASAP7_75t_L g1123 ( 
.A(n_967),
.B(n_970),
.Y(n_1123)
);

NAND3x1_ASAP7_75t_L g1124 ( 
.A(n_1086),
.B(n_987),
.C(n_991),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_951),
.A2(n_956),
.B(n_1065),
.Y(n_1125)
);

AO31x2_ASAP7_75t_L g1126 ( 
.A1(n_958),
.A2(n_1044),
.A3(n_1079),
.B(n_955),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_SL g1127 ( 
.A1(n_1033),
.A2(n_954),
.B(n_1027),
.C(n_1034),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1053),
.A2(n_1043),
.B(n_969),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_976),
.B(n_1023),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_1077),
.A2(n_1072),
.A3(n_1052),
.B(n_1010),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_1007),
.B(n_1009),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_1026),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1043),
.A2(n_1054),
.B(n_1057),
.Y(n_1133)
);

NAND3xp33_ASAP7_75t_SL g1134 ( 
.A(n_1093),
.B(n_996),
.C(n_998),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1024),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_976),
.B(n_1017),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1005),
.A2(n_960),
.B(n_1030),
.C(n_1020),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1057),
.A2(n_1059),
.B(n_1080),
.Y(n_1138)
);

AOI221xp5_ASAP7_75t_L g1139 ( 
.A1(n_983),
.A2(n_1013),
.B1(n_1030),
.B2(n_981),
.C(n_973),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1080),
.A2(n_1076),
.B(n_1064),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_984),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1076),
.A2(n_968),
.B(n_1048),
.Y(n_1142)
);

NAND2xp33_ASAP7_75t_L g1143 ( 
.A(n_953),
.B(n_1024),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_1009),
.B(n_1002),
.Y(n_1144)
);

AO31x2_ASAP7_75t_L g1145 ( 
.A1(n_1010),
.A2(n_973),
.A3(n_981),
.B(n_1067),
.Y(n_1145)
);

AND2x6_ASAP7_75t_L g1146 ( 
.A(n_1048),
.B(n_1039),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1046),
.A2(n_1034),
.B(n_1038),
.Y(n_1147)
);

INVxp67_ASAP7_75t_L g1148 ( 
.A(n_972),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1015),
.B(n_1047),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_SL g1150 ( 
.A(n_985),
.B(n_993),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1098),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1063),
.A2(n_1060),
.B(n_1058),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1055),
.B(n_1021),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1046),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1009),
.B(n_1002),
.Y(n_1155)
);

AO31x2_ASAP7_75t_L g1156 ( 
.A1(n_1010),
.A2(n_1061),
.A3(n_1070),
.B(n_1022),
.Y(n_1156)
);

INVx1_ASAP7_75t_SL g1157 ( 
.A(n_1001),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1038),
.A2(n_982),
.B(n_1045),
.C(n_1037),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_1041),
.Y(n_1159)
);

AOI221x1_ASAP7_75t_L g1160 ( 
.A1(n_1056),
.A2(n_1028),
.B1(n_1040),
.B2(n_1003),
.C(n_979),
.Y(n_1160)
);

INVx6_ASAP7_75t_L g1161 ( 
.A(n_1004),
.Y(n_1161)
);

NOR4xp25_ASAP7_75t_L g1162 ( 
.A(n_1069),
.B(n_1062),
.C(n_975),
.D(n_979),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_982),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1090),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_959),
.B(n_1050),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1074),
.A2(n_1081),
.B(n_1082),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1050),
.B(n_1090),
.Y(n_1167)
);

INVxp67_ASAP7_75t_L g1168 ( 
.A(n_1050),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1074),
.A2(n_1081),
.B(n_1071),
.Y(n_1169)
);

INVx5_ASAP7_75t_L g1170 ( 
.A(n_1056),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1036),
.B(n_968),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_986),
.A2(n_1008),
.B(n_1050),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1050),
.A2(n_1042),
.B(n_1079),
.Y(n_1173)
);

AOI221x1_ASAP7_75t_L g1174 ( 
.A1(n_1036),
.A2(n_1087),
.B1(n_1085),
.B2(n_841),
.C(n_1006),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_1088),
.A2(n_1087),
.A3(n_1085),
.B(n_1094),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1088),
.A2(n_994),
.B(n_810),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1088),
.A2(n_1087),
.A3(n_1085),
.B(n_1094),
.Y(n_1177)
);

O2A1O1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1085),
.A2(n_1087),
.B(n_1089),
.C(n_1083),
.Y(n_1178)
);

OA21x2_ASAP7_75t_L g1179 ( 
.A1(n_1088),
.A2(n_858),
.B(n_994),
.Y(n_1179)
);

AOI22x1_ASAP7_75t_L g1180 ( 
.A1(n_1088),
.A2(n_994),
.B1(n_858),
.B2(n_1042),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1088),
.A2(n_994),
.B(n_810),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1088),
.A2(n_994),
.B(n_810),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_950),
.A2(n_1084),
.B1(n_1087),
.B2(n_1085),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1086),
.B(n_997),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_999),
.B(n_841),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_990),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_999),
.B(n_841),
.Y(n_1187)
);

AO31x2_ASAP7_75t_L g1188 ( 
.A1(n_1088),
.A2(n_1087),
.A3(n_1085),
.B(n_1094),
.Y(n_1188)
);

AO21x2_ASAP7_75t_L g1189 ( 
.A1(n_1088),
.A2(n_788),
.B(n_858),
.Y(n_1189)
);

NOR2xp67_ASAP7_75t_L g1190 ( 
.A(n_997),
.B(n_854),
.Y(n_1190)
);

OAI221xp5_ASAP7_75t_L g1191 ( 
.A1(n_1092),
.A2(n_841),
.B1(n_447),
.B2(n_1087),
.C(n_1085),
.Y(n_1191)
);

NAND3xp33_ASAP7_75t_L g1192 ( 
.A(n_950),
.B(n_841),
.C(n_1084),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_963),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1007),
.B(n_1009),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1042),
.A2(n_1079),
.B(n_1065),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1042),
.A2(n_1079),
.B(n_1065),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1088),
.A2(n_994),
.B(n_810),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_963),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1091),
.B(n_1095),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_963),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_963),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1042),
.A2(n_1079),
.B(n_1065),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1088),
.A2(n_994),
.B(n_810),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_963),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_999),
.B(n_841),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1088),
.A2(n_994),
.B(n_810),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1042),
.A2(n_1079),
.B(n_1065),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_SL g1208 ( 
.A1(n_1085),
.A2(n_1087),
.B(n_1006),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1088),
.A2(n_994),
.B(n_810),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_963),
.Y(n_1210)
);

AO31x2_ASAP7_75t_L g1211 ( 
.A1(n_1088),
.A2(n_1087),
.A3(n_1085),
.B(n_1094),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1042),
.A2(n_1079),
.B(n_1065),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1091),
.B(n_1095),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1088),
.A2(n_994),
.B(n_810),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_962),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1088),
.A2(n_994),
.B(n_810),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1085),
.A2(n_1087),
.B(n_1089),
.C(n_1083),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1042),
.A2(n_1079),
.B(n_1065),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_999),
.B(n_841),
.Y(n_1219)
);

O2A1O1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1085),
.A2(n_1087),
.B(n_1089),
.C(n_1083),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1042),
.A2(n_1079),
.B(n_1065),
.Y(n_1221)
);

AO22x2_ASAP7_75t_L g1222 ( 
.A1(n_1096),
.A2(n_1097),
.B1(n_1094),
.B2(n_520),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_SL g1223 ( 
.A1(n_1085),
.A2(n_1087),
.B(n_1006),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_963),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_SL g1225 ( 
.A1(n_1085),
.A2(n_1087),
.B(n_1006),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_963),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1086),
.B(n_997),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1042),
.A2(n_1079),
.B(n_1065),
.Y(n_1228)
);

INVx3_ASAP7_75t_SL g1229 ( 
.A(n_984),
.Y(n_1229)
);

BUFx10_ASAP7_75t_L g1230 ( 
.A(n_984),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1042),
.A2(n_1079),
.B(n_1065),
.Y(n_1231)
);

BUFx10_ASAP7_75t_L g1232 ( 
.A(n_984),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1042),
.A2(n_1079),
.B(n_1065),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1085),
.A2(n_841),
.B(n_1087),
.C(n_1083),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_963),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_1026),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1088),
.A2(n_994),
.B(n_810),
.Y(n_1237)
);

HB1xp67_ASAP7_75t_L g1238 ( 
.A(n_1020),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1088),
.A2(n_994),
.B(n_810),
.Y(n_1239)
);

NOR2xp67_ASAP7_75t_L g1240 ( 
.A(n_997),
.B(n_854),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1088),
.A2(n_994),
.B(n_810),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_962),
.Y(n_1242)
);

AO31x2_ASAP7_75t_L g1243 ( 
.A1(n_1088),
.A2(n_1087),
.A3(n_1085),
.B(n_1094),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1184),
.B(n_1227),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1141),
.Y(n_1245)
);

BUFx4f_ASAP7_75t_SL g1246 ( 
.A(n_1229),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_1101),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1185),
.B(n_1187),
.Y(n_1248)
);

OAI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1219),
.A2(n_1191),
.B1(n_1192),
.B2(n_1100),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1186),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1176),
.A2(n_1182),
.B(n_1181),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1105),
.A2(n_1205),
.B1(n_1183),
.B2(n_1149),
.Y(n_1252)
);

CKINVDCx8_ASAP7_75t_R g1253 ( 
.A(n_1132),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_1230),
.Y(n_1254)
);

CKINVDCx11_ASAP7_75t_R g1255 ( 
.A(n_1230),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1235),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_1232),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1134),
.A2(n_1153),
.B1(n_1240),
.B2(n_1190),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1199),
.B(n_1213),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1107),
.B(n_1157),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1099),
.A2(n_1222),
.B1(n_1114),
.B2(n_1139),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1108),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1242),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1222),
.A2(n_1150),
.B1(n_1124),
.B2(n_1111),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_SL g1265 ( 
.A1(n_1163),
.A2(n_1102),
.B1(n_1115),
.B2(n_1172),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1189),
.A2(n_1180),
.B1(n_1136),
.B2(n_1179),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1113),
.Y(n_1267)
);

INVx6_ASAP7_75t_L g1268 ( 
.A(n_1159),
.Y(n_1268)
);

INVx3_ASAP7_75t_L g1269 ( 
.A(n_1104),
.Y(n_1269)
);

INVxp67_ASAP7_75t_SL g1270 ( 
.A(n_1238),
.Y(n_1270)
);

BUFx12f_ASAP7_75t_L g1271 ( 
.A(n_1232),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1180),
.A2(n_1179),
.B1(n_1154),
.B2(n_1133),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1234),
.A2(n_1102),
.B1(n_1122),
.B2(n_1225),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1128),
.A2(n_1174),
.B(n_1223),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1193),
.Y(n_1275)
);

BUFx10_ASAP7_75t_L g1276 ( 
.A(n_1132),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1154),
.A2(n_1129),
.B1(n_1147),
.B2(n_1151),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1165),
.A2(n_1152),
.B1(n_1210),
.B2(n_1198),
.Y(n_1278)
);

INVx6_ASAP7_75t_L g1279 ( 
.A(n_1159),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1200),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1201),
.A2(n_1204),
.B1(n_1226),
.B2(n_1224),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1144),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1123),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1168),
.A2(n_1217),
.B1(n_1178),
.B2(n_1220),
.Y(n_1284)
);

BUFx12f_ASAP7_75t_L g1285 ( 
.A(n_1132),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1236),
.A2(n_1146),
.B1(n_1117),
.B2(n_1208),
.Y(n_1286)
);

CKINVDCx11_ASAP7_75t_R g1287 ( 
.A(n_1236),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1155),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1103),
.A2(n_1155),
.B1(n_1146),
.B2(n_1148),
.Y(n_1289)
);

CKINVDCx8_ASAP7_75t_R g1290 ( 
.A(n_1236),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1167),
.A2(n_1140),
.B1(n_1137),
.B2(n_1158),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1171),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1116),
.B(n_1175),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1104),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1161),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_1131),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1121),
.A2(n_1146),
.B1(n_1138),
.B2(n_1166),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1156),
.Y(n_1298)
);

INVx8_ASAP7_75t_L g1299 ( 
.A(n_1170),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1131),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1146),
.A2(n_1117),
.B1(n_1109),
.B2(n_1118),
.Y(n_1301)
);

CKINVDCx11_ASAP7_75t_R g1302 ( 
.A(n_1194),
.Y(n_1302)
);

BUFx12f_ASAP7_75t_L g1303 ( 
.A(n_1161),
.Y(n_1303)
);

OAI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1170),
.A2(n_1160),
.B1(n_1169),
.B2(n_1135),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1117),
.A2(n_1209),
.B1(n_1241),
.B2(n_1239),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1117),
.A2(n_1194),
.B1(n_1127),
.B2(n_1162),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1197),
.A2(n_1237),
.B1(n_1216),
.B2(n_1214),
.Y(n_1307)
);

INVx4_ASAP7_75t_L g1308 ( 
.A(n_1170),
.Y(n_1308)
);

BUFx12f_ASAP7_75t_SL g1309 ( 
.A(n_1110),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_1164),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_1164),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1203),
.A2(n_1206),
.B(n_1125),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1173),
.A2(n_1142),
.B1(n_1211),
.B2(n_1188),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1143),
.A2(n_1106),
.B1(n_1233),
.B2(n_1231),
.Y(n_1314)
);

CKINVDCx11_ASAP7_75t_R g1315 ( 
.A(n_1120),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1175),
.A2(n_1211),
.B1(n_1188),
.B2(n_1177),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1112),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1175),
.A2(n_1243),
.B1(n_1211),
.B2(n_1188),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1177),
.A2(n_1243),
.B1(n_1202),
.B2(n_1207),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1177),
.A2(n_1243),
.B1(n_1196),
.B2(n_1212),
.Y(n_1320)
);

CKINVDCx11_ASAP7_75t_R g1321 ( 
.A(n_1145),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1126),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1119),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1130),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1195),
.A2(n_1218),
.B1(n_1221),
.B2(n_1228),
.Y(n_1325)
);

BUFx10_ASAP7_75t_L g1326 ( 
.A(n_1130),
.Y(n_1326)
);

CKINVDCx6p67_ASAP7_75t_R g1327 ( 
.A(n_1145),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1119),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_1141),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_SL g1330 ( 
.A1(n_1185),
.A2(n_520),
.B(n_1187),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1215),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1185),
.A2(n_1219),
.B1(n_1187),
.B2(n_841),
.Y(n_1332)
);

INVx8_ASAP7_75t_L g1333 ( 
.A(n_1159),
.Y(n_1333)
);

OAI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1185),
.A2(n_1219),
.B1(n_1187),
.B2(n_1191),
.Y(n_1334)
);

BUFx6f_ASAP7_75t_SL g1335 ( 
.A(n_1132),
.Y(n_1335)
);

CKINVDCx11_ASAP7_75t_R g1336 ( 
.A(n_1229),
.Y(n_1336)
);

INVx4_ASAP7_75t_L g1337 ( 
.A(n_1159),
.Y(n_1337)
);

NAND2x1p5_ASAP7_75t_L g1338 ( 
.A(n_1170),
.B(n_1008),
.Y(n_1338)
);

AOI22xp5_ASAP7_75t_SL g1339 ( 
.A1(n_1185),
.A2(n_1187),
.B1(n_1219),
.B2(n_980),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1185),
.A2(n_1219),
.B1(n_1187),
.B2(n_950),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1185),
.A2(n_1219),
.B1(n_1187),
.B2(n_950),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_SL g1342 ( 
.A1(n_1185),
.A2(n_1219),
.B1(n_1187),
.B2(n_841),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1185),
.A2(n_1219),
.B1(n_1187),
.B2(n_950),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1192),
.A2(n_1187),
.B1(n_1219),
.B2(n_1185),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1215),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_1141),
.Y(n_1346)
);

INVx5_ASAP7_75t_L g1347 ( 
.A(n_1159),
.Y(n_1347)
);

INVxp67_ASAP7_75t_SL g1348 ( 
.A(n_1238),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1103),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1186),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1185),
.A2(n_1219),
.B1(n_1187),
.B2(n_841),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1192),
.A2(n_1187),
.B1(n_1219),
.B2(n_1185),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1192),
.A2(n_1187),
.B1(n_1219),
.B2(n_1185),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1293),
.B(n_1322),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1274),
.B(n_1350),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_1317),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1299),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1324),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1299),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_SL g1360 ( 
.A(n_1340),
.B(n_1341),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1344),
.B(n_1352),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_1260),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1298),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1299),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1270),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1348),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1312),
.A2(n_1251),
.B(n_1305),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1249),
.A2(n_1343),
.B1(n_1334),
.B2(n_1273),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_1328),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1292),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1323),
.Y(n_1371)
);

NAND2xp33_ASAP7_75t_R g1372 ( 
.A(n_1254),
.B(n_1245),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1344),
.B(n_1352),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1250),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1275),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1315),
.Y(n_1376)
);

INVxp33_ASAP7_75t_L g1377 ( 
.A(n_1244),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1306),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1326),
.Y(n_1379)
);

NAND2x1p5_ASAP7_75t_L g1380 ( 
.A(n_1314),
.B(n_1308),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1347),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1332),
.A2(n_1351),
.B1(n_1342),
.B2(n_1353),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1305),
.A2(n_1307),
.B(n_1325),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1261),
.B(n_1316),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1353),
.B(n_1259),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1327),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1307),
.A2(n_1320),
.B(n_1319),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1249),
.B(n_1334),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1310),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1267),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1291),
.Y(n_1391)
);

INVxp67_ASAP7_75t_R g1392 ( 
.A(n_1255),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1261),
.B(n_1316),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1318),
.B(n_1284),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1252),
.A2(n_1265),
.B1(n_1284),
.B2(n_1264),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1280),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1301),
.B(n_1256),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1281),
.Y(n_1398)
);

BUFx2_ASAP7_75t_R g1399 ( 
.A(n_1253),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1321),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1281),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1311),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1272),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1272),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1318),
.B(n_1266),
.Y(n_1405)
);

OAI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1339),
.A2(n_1330),
.B(n_1278),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1266),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1289),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1313),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1347),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1313),
.Y(n_1411)
);

BUFx12f_ASAP7_75t_L g1412 ( 
.A(n_1287),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_L g1413 ( 
.A(n_1288),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1319),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_L g1415 ( 
.A(n_1248),
.B(n_1277),
.C(n_1278),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1277),
.A2(n_1297),
.B(n_1301),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1320),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1304),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1304),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1297),
.A2(n_1338),
.B(n_1294),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1300),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1286),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1347),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1283),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1263),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1300),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1372),
.Y(n_1427)
);

A2O1A1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1360),
.A2(n_1258),
.B(n_1263),
.C(n_1296),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1362),
.B(n_1349),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1368),
.A2(n_1290),
.B1(n_1257),
.B2(n_1345),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1377),
.B(n_1346),
.Y(n_1431)
);

A2O1A1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1406),
.A2(n_1262),
.B(n_1331),
.C(n_1282),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1396),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_L g1434 ( 
.A(n_1389),
.Y(n_1434)
);

BUFx12f_ASAP7_75t_L g1435 ( 
.A(n_1412),
.Y(n_1435)
);

AOI221xp5_ASAP7_75t_L g1436 ( 
.A1(n_1382),
.A2(n_1406),
.B1(n_1391),
.B2(n_1361),
.C(n_1373),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1395),
.A2(n_1331),
.B1(n_1335),
.B2(n_1268),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1388),
.A2(n_1335),
.B1(n_1302),
.B2(n_1285),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1385),
.B(n_1329),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1389),
.B(n_1246),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1374),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1375),
.B(n_1269),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1365),
.B(n_1366),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1382),
.A2(n_1268),
.B1(n_1279),
.B2(n_1337),
.Y(n_1444)
);

A2O1A1Ixp33_ASAP7_75t_L g1445 ( 
.A1(n_1391),
.A2(n_1333),
.B(n_1295),
.C(n_1247),
.Y(n_1445)
);

A2O1A1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1416),
.A2(n_1333),
.B(n_1309),
.C(n_1279),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_SL g1447 ( 
.A(n_1399),
.B(n_1412),
.Y(n_1447)
);

INVx2_ASAP7_75t_SL g1448 ( 
.A(n_1389),
.Y(n_1448)
);

OR2x6_ASAP7_75t_L g1449 ( 
.A(n_1412),
.B(n_1416),
.Y(n_1449)
);

O2A1O1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1415),
.A2(n_1276),
.B(n_1333),
.C(n_1268),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1400),
.B(n_1276),
.Y(n_1451)
);

AO32x2_ASAP7_75t_L g1452 ( 
.A1(n_1381),
.A2(n_1423),
.A3(n_1410),
.B1(n_1354),
.B2(n_1419),
.Y(n_1452)
);

OR2x6_ASAP7_75t_L g1453 ( 
.A(n_1376),
.B(n_1271),
.Y(n_1453)
);

OR2x6_ASAP7_75t_L g1454 ( 
.A(n_1376),
.B(n_1303),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1354),
.B(n_1336),
.Y(n_1455)
);

AO32x2_ASAP7_75t_L g1456 ( 
.A1(n_1381),
.A2(n_1423),
.A3(n_1410),
.B1(n_1419),
.B2(n_1356),
.Y(n_1456)
);

NOR2x1_ASAP7_75t_SL g1457 ( 
.A(n_1376),
.B(n_1415),
.Y(n_1457)
);

INVxp33_ASAP7_75t_L g1458 ( 
.A(n_1402),
.Y(n_1458)
);

AOI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1378),
.A2(n_1422),
.B1(n_1408),
.B2(n_1376),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1378),
.A2(n_1376),
.B1(n_1422),
.B2(n_1408),
.Y(n_1460)
);

A2O1A1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1418),
.A2(n_1408),
.B(n_1356),
.C(n_1394),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1421),
.B(n_1426),
.Y(n_1462)
);

OAI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1383),
.A2(n_1420),
.B(n_1367),
.Y(n_1463)
);

OR2x6_ASAP7_75t_L g1464 ( 
.A(n_1420),
.B(n_1357),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1394),
.A2(n_1402),
.B1(n_1418),
.B2(n_1393),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1421),
.B(n_1426),
.Y(n_1466)
);

AO32x2_ASAP7_75t_L g1467 ( 
.A1(n_1355),
.A2(n_1370),
.A3(n_1409),
.B1(n_1411),
.B2(n_1371),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1383),
.A2(n_1367),
.B(n_1387),
.Y(n_1468)
);

OAI221xp5_ASAP7_75t_L g1469 ( 
.A1(n_1424),
.A2(n_1402),
.B1(n_1425),
.B2(n_1380),
.C(n_1386),
.Y(n_1469)
);

AOI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1384),
.A2(n_1393),
.B1(n_1401),
.B2(n_1398),
.Y(n_1470)
);

AOI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1384),
.A2(n_1401),
.B1(n_1398),
.B2(n_1392),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1424),
.B(n_1413),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1441),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1467),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1467),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1467),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1436),
.A2(n_1461),
.B1(n_1465),
.B2(n_1459),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1471),
.B(n_1386),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1452),
.B(n_1411),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1433),
.B(n_1407),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1452),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_SL g1482 ( 
.A1(n_1457),
.A2(n_1397),
.B1(n_1403),
.B2(n_1404),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1468),
.B(n_1387),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1463),
.B(n_1417),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1464),
.B(n_1417),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1456),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1443),
.B(n_1407),
.Y(n_1487)
);

NAND2x1_ASAP7_75t_L g1488 ( 
.A(n_1464),
.B(n_1379),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1456),
.B(n_1414),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1429),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1470),
.B(n_1404),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1469),
.B(n_1390),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1456),
.Y(n_1493)
);

CKINVDCx20_ASAP7_75t_R g1494 ( 
.A(n_1427),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1472),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1442),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1428),
.A2(n_1405),
.B1(n_1403),
.B2(n_1397),
.Y(n_1497)
);

INVx5_ASAP7_75t_L g1498 ( 
.A(n_1449),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1462),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1466),
.B(n_1369),
.Y(n_1500)
);

NOR2x1_ASAP7_75t_L g1501 ( 
.A(n_1449),
.B(n_1379),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1483),
.B(n_1363),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1487),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1478),
.B(n_1458),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1473),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1488),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1494),
.Y(n_1507)
);

INVx3_ASAP7_75t_L g1508 ( 
.A(n_1488),
.Y(n_1508)
);

INVx2_ASAP7_75t_SL g1509 ( 
.A(n_1488),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1486),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1483),
.B(n_1405),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1500),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1474),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1475),
.Y(n_1514)
);

AOI211xp5_ASAP7_75t_SL g1515 ( 
.A1(n_1477),
.A2(n_1432),
.B(n_1460),
.C(n_1446),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1498),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1476),
.B(n_1358),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1480),
.Y(n_1518)
);

OAI221xp5_ASAP7_75t_L g1519 ( 
.A1(n_1477),
.A2(n_1438),
.B1(n_1437),
.B2(n_1445),
.C(n_1430),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1482),
.A2(n_1454),
.B1(n_1453),
.B2(n_1455),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1493),
.Y(n_1521)
);

A2O1A1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1492),
.A2(n_1439),
.B(n_1450),
.C(n_1447),
.Y(n_1522)
);

AOI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1497),
.A2(n_1444),
.B1(n_1453),
.B2(n_1397),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1493),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1505),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1503),
.B(n_1481),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1510),
.B(n_1512),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1520),
.B(n_1498),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1511),
.B(n_1496),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1510),
.B(n_1479),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1521),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1512),
.B(n_1499),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1511),
.B(n_1496),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1521),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_1506),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1505),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1516),
.B(n_1485),
.Y(n_1537)
);

INVx4_ASAP7_75t_L g1538 ( 
.A(n_1507),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1518),
.B(n_1487),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1514),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1518),
.B(n_1480),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1514),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1511),
.B(n_1489),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1517),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1518),
.B(n_1480),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1519),
.A2(n_1497),
.B1(n_1478),
.B2(n_1482),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1516),
.B(n_1485),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1514),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1506),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1546),
.B(n_1511),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1538),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1531),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1546),
.B(n_1492),
.Y(n_1553)
);

INVx3_ASAP7_75t_L g1554 ( 
.A(n_1540),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1531),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1534),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1535),
.B(n_1506),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1543),
.B(n_1510),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1534),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1527),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1543),
.B(n_1521),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1537),
.B(n_1512),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1541),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1541),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1545),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1527),
.Y(n_1566)
);

OAI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1528),
.A2(n_1522),
.B(n_1515),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1537),
.B(n_1547),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1530),
.Y(n_1569)
);

NAND3xp33_ASAP7_75t_L g1570 ( 
.A(n_1538),
.B(n_1515),
.C(n_1522),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1545),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1527),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1539),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1540),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1537),
.B(n_1512),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1539),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1535),
.B(n_1506),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1537),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1529),
.B(n_1521),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1529),
.B(n_1524),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1533),
.B(n_1504),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1540),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1547),
.B(n_1512),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1547),
.B(n_1512),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1542),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1533),
.B(n_1504),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1542),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1542),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1548),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1547),
.B(n_1495),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1535),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1568),
.B(n_1549),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1557),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1568),
.B(n_1549),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1578),
.B(n_1530),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1567),
.A2(n_1519),
.B1(n_1520),
.B2(n_1538),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1552),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1552),
.Y(n_1598)
);

NAND2x1_ASAP7_75t_L g1599 ( 
.A(n_1557),
.B(n_1530),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1573),
.B(n_1526),
.Y(n_1600)
);

NAND3xp33_ASAP7_75t_SL g1601 ( 
.A(n_1570),
.B(n_1507),
.C(n_1523),
.Y(n_1601)
);

INVxp67_ASAP7_75t_SL g1602 ( 
.A(n_1578),
.Y(n_1602)
);

OAI21x1_ASAP7_75t_L g1603 ( 
.A1(n_1578),
.A2(n_1508),
.B(n_1548),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1569),
.B(n_1532),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1553),
.B(n_1538),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1557),
.B(n_1532),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1555),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1551),
.B(n_1502),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1554),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1573),
.B(n_1526),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1557),
.B(n_1509),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1550),
.B(n_1502),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1581),
.A2(n_1392),
.B(n_1494),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1577),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1576),
.B(n_1544),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1555),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1577),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1556),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1577),
.B(n_1509),
.Y(n_1619)
);

NOR2x1_ASAP7_75t_L g1620 ( 
.A(n_1577),
.B(n_1556),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1559),
.Y(n_1621)
);

OAI21xp33_ASAP7_75t_L g1622 ( 
.A1(n_1586),
.A2(n_1523),
.B(n_1491),
.Y(n_1622)
);

OAI31xp33_ASAP7_75t_L g1623 ( 
.A1(n_1591),
.A2(n_1516),
.A3(n_1448),
.B(n_1484),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1559),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1590),
.B(n_1502),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1563),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1596),
.B(n_1576),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1597),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1597),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1592),
.B(n_1594),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1620),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1598),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1592),
.B(n_1591),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1593),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1605),
.B(n_1563),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1598),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1622),
.B(n_1564),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1622),
.B(n_1564),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1607),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1607),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1601),
.A2(n_1523),
.B1(n_1516),
.B2(n_1484),
.Y(n_1641)
);

OAI21xp33_ASAP7_75t_L g1642 ( 
.A1(n_1594),
.A2(n_1571),
.B(n_1565),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1620),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1616),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1616),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1602),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1618),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1593),
.B(n_1562),
.Y(n_1648)
);

OAI21xp33_ASAP7_75t_SL g1649 ( 
.A1(n_1623),
.A2(n_1575),
.B(n_1562),
.Y(n_1649)
);

OAI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1613),
.A2(n_1501),
.B(n_1565),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1599),
.A2(n_1454),
.B1(n_1558),
.B2(n_1498),
.Y(n_1651)
);

OAI221xp5_ASAP7_75t_L g1652 ( 
.A1(n_1641),
.A2(n_1623),
.B1(n_1599),
.B2(n_1626),
.C(n_1614),
.Y(n_1652)
);

NAND4xp25_ASAP7_75t_SL g1653 ( 
.A(n_1627),
.B(n_1612),
.C(n_1606),
.D(n_1595),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1630),
.A2(n_1626),
.B1(n_1608),
.B2(n_1606),
.Y(n_1654)
);

NAND4xp25_ASAP7_75t_SL g1655 ( 
.A(n_1650),
.B(n_1595),
.C(n_1604),
.D(n_1619),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1630),
.B(n_1604),
.Y(n_1656)
);

AOI21xp33_ASAP7_75t_SL g1657 ( 
.A1(n_1643),
.A2(n_1440),
.B(n_1593),
.Y(n_1657)
);

NOR3xp33_ASAP7_75t_L g1658 ( 
.A(n_1646),
.B(n_1621),
.C(n_1618),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1628),
.Y(n_1659)
);

AOI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1637),
.A2(n_1621),
.B1(n_1624),
.B2(n_1593),
.C(n_1617),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1633),
.B(n_1614),
.Y(n_1661)
);

OAI221xp5_ASAP7_75t_SL g1662 ( 
.A1(n_1638),
.A2(n_1600),
.B1(n_1610),
.B2(n_1624),
.C(n_1558),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_1633),
.Y(n_1663)
);

AOI21xp33_ASAP7_75t_L g1664 ( 
.A1(n_1631),
.A2(n_1617),
.B(n_1614),
.Y(n_1664)
);

INVxp67_ASAP7_75t_L g1665 ( 
.A(n_1634),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1648),
.Y(n_1666)
);

A2O1A1Ixp33_ASAP7_75t_L g1667 ( 
.A1(n_1642),
.A2(n_1617),
.B(n_1614),
.C(n_1610),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1635),
.B(n_1617),
.Y(n_1668)
);

AOI21xp33_ASAP7_75t_L g1669 ( 
.A1(n_1651),
.A2(n_1600),
.B(n_1615),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1649),
.A2(n_1619),
.B(n_1611),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1665),
.Y(n_1671)
);

XOR2xp5_ASAP7_75t_L g1672 ( 
.A(n_1653),
.B(n_1434),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1663),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1666),
.B(n_1634),
.Y(n_1674)
);

O2A1O1Ixp33_ASAP7_75t_L g1675 ( 
.A1(n_1662),
.A2(n_1640),
.B(n_1636),
.C(n_1645),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1661),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1656),
.B(n_1639),
.Y(n_1677)
);

AOI211xp5_ASAP7_75t_SL g1678 ( 
.A1(n_1662),
.A2(n_1644),
.B(n_1647),
.C(n_1628),
.Y(n_1678)
);

XOR2x2_ASAP7_75t_L g1679 ( 
.A(n_1658),
.B(n_1431),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1652),
.A2(n_1648),
.B1(n_1625),
.B2(n_1509),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1665),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1670),
.B(n_1611),
.Y(n_1682)
);

NOR3xp33_ASAP7_75t_SL g1683 ( 
.A(n_1680),
.B(n_1655),
.C(n_1667),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1674),
.Y(n_1684)
);

XOR2xp5_ASAP7_75t_L g1685 ( 
.A(n_1679),
.B(n_1672),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_L g1686 ( 
.A(n_1678),
.B(n_1660),
.C(n_1657),
.Y(n_1686)
);

INVxp67_ASAP7_75t_L g1687 ( 
.A(n_1682),
.Y(n_1687)
);

O2A1O1Ixp5_ASAP7_75t_L g1688 ( 
.A1(n_1671),
.A2(n_1664),
.B(n_1669),
.C(n_1668),
.Y(n_1688)
);

NOR3xp33_ASAP7_75t_L g1689 ( 
.A(n_1673),
.B(n_1659),
.C(n_1632),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1673),
.B(n_1654),
.Y(n_1690)
);

NAND3xp33_ASAP7_75t_L g1691 ( 
.A(n_1675),
.B(n_1632),
.C(n_1629),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1681),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1685),
.B(n_1676),
.Y(n_1693)
);

NAND4xp25_ASAP7_75t_L g1694 ( 
.A(n_1686),
.B(n_1677),
.C(n_1647),
.D(n_1629),
.Y(n_1694)
);

NAND3xp33_ASAP7_75t_SL g1695 ( 
.A(n_1688),
.B(n_1615),
.C(n_1566),
.Y(n_1695)
);

OAI211xp5_ASAP7_75t_SL g1696 ( 
.A1(n_1683),
.A2(n_1609),
.B(n_1571),
.C(n_1572),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1691),
.A2(n_1609),
.B1(n_1566),
.B2(n_1572),
.C(n_1560),
.Y(n_1697)
);

OAI211xp5_ASAP7_75t_SL g1698 ( 
.A1(n_1693),
.A2(n_1687),
.B(n_1690),
.C(n_1684),
.Y(n_1698)
);

OAI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1694),
.A2(n_1689),
.B1(n_1692),
.B2(n_1609),
.C(n_1560),
.Y(n_1699)
);

AOI211xp5_ASAP7_75t_L g1700 ( 
.A1(n_1696),
.A2(n_1451),
.B(n_1603),
.C(n_1575),
.Y(n_1700)
);

OAI221xp5_ASAP7_75t_L g1701 ( 
.A1(n_1695),
.A2(n_1434),
.B1(n_1509),
.B2(n_1588),
.C(n_1589),
.Y(n_1701)
);

NOR3xp33_ASAP7_75t_L g1702 ( 
.A(n_1697),
.B(n_1435),
.C(n_1603),
.Y(n_1702)
);

AOI211xp5_ASAP7_75t_L g1703 ( 
.A1(n_1696),
.A2(n_1583),
.B(n_1584),
.C(n_1434),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1698),
.A2(n_1584),
.B1(n_1583),
.B2(n_1587),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1703),
.B(n_1561),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1699),
.Y(n_1706)
);

NAND2xp33_ASAP7_75t_SL g1707 ( 
.A(n_1701),
.B(n_1579),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1700),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1706),
.B(n_1702),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1708),
.B(n_1561),
.Y(n_1710)
);

NAND4xp75_ASAP7_75t_L g1711 ( 
.A(n_1705),
.B(n_1501),
.C(n_1588),
.D(n_1587),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1711),
.Y(n_1712)
);

AO22x2_ASAP7_75t_L g1713 ( 
.A1(n_1712),
.A2(n_1709),
.B1(n_1710),
.B2(n_1707),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1713),
.B(n_1704),
.Y(n_1714)
);

OA22x2_ASAP7_75t_L g1715 ( 
.A1(n_1713),
.A2(n_1554),
.B1(n_1574),
.B2(n_1582),
.Y(n_1715)
);

OAI22x1_ASAP7_75t_L g1716 ( 
.A1(n_1714),
.A2(n_1574),
.B1(n_1554),
.B2(n_1582),
.Y(n_1716)
);

OAI22x1_ASAP7_75t_L g1717 ( 
.A1(n_1715),
.A2(n_1554),
.B1(n_1585),
.B2(n_1589),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1716),
.Y(n_1718)
);

AOI22x1_ASAP7_75t_L g1719 ( 
.A1(n_1717),
.A2(n_1585),
.B1(n_1548),
.B2(n_1579),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1718),
.Y(n_1720)
);

OA21x2_ASAP7_75t_L g1721 ( 
.A1(n_1720),
.A2(n_1719),
.B(n_1580),
.Y(n_1721)
);

OAI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1721),
.A2(n_1580),
.B1(n_1536),
.B2(n_1525),
.Y(n_1722)
);

OAI221xp5_ASAP7_75t_L g1723 ( 
.A1(n_1722),
.A2(n_1364),
.B1(n_1359),
.B2(n_1490),
.C(n_1514),
.Y(n_1723)
);

AOI211xp5_ASAP7_75t_L g1724 ( 
.A1(n_1723),
.A2(n_1364),
.B(n_1359),
.C(n_1513),
.Y(n_1724)
);


endmodule