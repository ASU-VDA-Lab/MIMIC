module fake_jpeg_8693_n_326 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_9),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_40),
.Y(n_50)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_43),
.Y(n_57)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_44),
.Y(n_48)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_17),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_55),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_17),
.B1(n_18),
.B2(n_23),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_51),
.A2(n_62),
.B1(n_65),
.B2(n_67),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_25),
.C(n_18),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_69),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_70),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_59),
.B(n_68),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_28),
.Y(n_61)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_31),
.B1(n_18),
.B2(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

OR2x2_ASAP7_75t_SL g94 ( 
.A(n_63),
.B(n_46),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_31),
.B1(n_23),
.B2(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_17),
.Y(n_66)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_28),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_30),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_26),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_26),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_45),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_34),
.B1(n_22),
.B2(n_26),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_73),
.B1(n_45),
.B2(n_40),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_44),
.A2(n_22),
.B1(n_34),
.B2(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_43),
.B(n_34),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_52),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_27),
.B1(n_30),
.B2(n_32),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_75),
.A2(n_35),
.B1(n_29),
.B2(n_20),
.Y(n_110)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_79),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_80),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_87),
.Y(n_123)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_54),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_82),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_35),
.B1(n_32),
.B2(n_20),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_89),
.B(n_71),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_93),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_94),
.A2(n_74),
.B(n_50),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_48),
.A2(n_46),
.B1(n_45),
.B2(n_40),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_99),
.A2(n_102),
.B1(n_67),
.B2(n_51),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_45),
.B1(n_40),
.B2(n_46),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_60),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_104),
.B(n_111),
.Y(n_117)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_61),
.Y(n_119)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_58),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_60),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_112),
.B(n_50),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_48),
.C(n_47),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_128),
.C(n_134),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_119),
.A2(n_85),
.B1(n_108),
.B2(n_98),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_63),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_120),
.A2(n_134),
.B(n_139),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_125),
.B(n_141),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_68),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_133),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_97),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_49),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_86),
.A2(n_66),
.B(n_70),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_100),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_110),
.B1(n_102),
.B2(n_94),
.Y(n_148)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_96),
.A2(n_36),
.A3(n_19),
.B1(n_27),
.B2(n_30),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_92),
.A2(n_19),
.B(n_36),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g141 ( 
.A(n_78),
.B(n_19),
.CI(n_21),
.CON(n_141),
.SN(n_141)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_136),
.A2(n_88),
.B(n_111),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_144),
.A2(n_149),
.B(n_150),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_145),
.B(n_121),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_125),
.B(n_90),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_146),
.B(n_155),
.Y(n_205)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_147),
.B(n_151),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_148),
.A2(n_158),
.B1(n_159),
.B2(n_130),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_111),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_114),
.A2(n_99),
.B(n_76),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_124),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_101),
.Y(n_153)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_153),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_171),
.C(n_118),
.Y(n_179)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_114),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_157),
.Y(n_176)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_101),
.B1(n_76),
.B2(n_36),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_95),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_160),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_129),
.A2(n_29),
.B1(n_21),
.B2(n_27),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_161),
.A2(n_115),
.B(n_122),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_135),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_163),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_95),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_167),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_80),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_168),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_133),
.B(n_97),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_120),
.Y(n_168)
);

BUFx24_ASAP7_75t_SL g169 ( 
.A(n_141),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_169),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_124),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_170),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_80),
.C(n_83),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_120),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_120),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_173),
.B(n_130),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_124),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_174),
.A2(n_122),
.B(n_115),
.Y(n_177)
);

INVxp33_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_191),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_177),
.A2(n_178),
.B(n_185),
.Y(n_214)
);

AOI211xp5_ASAP7_75t_SL g178 ( 
.A1(n_166),
.A2(n_138),
.B(n_141),
.C(n_119),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_182),
.C(n_195),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_180),
.B(n_200),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_141),
.Y(n_182)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_143),
.A2(n_164),
.B1(n_172),
.B2(n_168),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_189),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_190),
.B(n_203),
.Y(n_228)
);

OAI211xp5_ASAP7_75t_L g192 ( 
.A1(n_152),
.A2(n_138),
.B(n_130),
.C(n_121),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_201),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_121),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_145),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_143),
.A2(n_135),
.B1(n_140),
.B2(n_118),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_159),
.A2(n_127),
.B1(n_113),
.B2(n_126),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_148),
.A2(n_155),
.B1(n_158),
.B2(n_166),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_162),
.Y(n_201)
);

AOI221xp5_ASAP7_75t_L g203 ( 
.A1(n_144),
.A2(n_113),
.B1(n_127),
.B2(n_21),
.C(n_126),
.Y(n_203)
);

MAJx2_ASAP7_75t_L g204 ( 
.A(n_149),
.B(n_109),
.C(n_1),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_173),
.C(n_142),
.Y(n_225)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_211),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_184),
.A2(n_201),
.B1(n_174),
.B2(n_196),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_187),
.B1(n_204),
.B2(n_145),
.Y(n_240)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_205),
.B(n_156),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_212),
.B(n_213),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_177),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_221),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_176),
.B(n_157),
.Y(n_219)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_152),
.Y(n_220)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_201),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_198),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_230),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_199),
.A2(n_189),
.B1(n_197),
.B2(n_181),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_223),
.A2(n_227),
.B1(n_187),
.B2(n_195),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_181),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_224),
.B(n_3),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_183),
.C(n_2),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_180),
.A2(n_149),
.B1(n_147),
.B2(n_150),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_229),
.B(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_185),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_0),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_161),
.Y(n_232)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_232),
.Y(n_237)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_16),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_216),
.A2(n_178),
.B1(n_179),
.B2(n_191),
.Y(n_234)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_234),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_182),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_244),
.C(n_256),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_240),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_243),
.A2(n_247),
.B(n_249),
.Y(n_257)
);

OAI322xp33_ASAP7_75t_L g245 ( 
.A1(n_220),
.A2(n_11),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_6),
.C2(n_8),
.Y(n_245)
);

NOR3xp33_ASAP7_75t_SL g271 ( 
.A(n_245),
.B(n_10),
.C(n_11),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_231),
.A2(n_82),
.B1(n_103),
.B2(n_0),
.Y(n_246)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_214),
.A2(n_0),
.B(n_2),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_208),
.A2(n_103),
.B1(n_0),
.B2(n_4),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_207),
.A2(n_3),
.B1(n_6),
.B2(n_8),
.Y(n_251)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_251),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_253),
.Y(n_265)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_219),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_211),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_214),
.B(n_8),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_209),
.Y(n_258)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_258),
.Y(n_287)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_217),
.C(n_226),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_273),
.C(n_259),
.Y(n_277)
);

AO221x1_ASAP7_75t_L g266 ( 
.A1(n_236),
.A2(n_213),
.B1(n_233),
.B2(n_207),
.C(n_227),
.Y(n_266)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_236),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_267),
.B(n_255),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_237),
.Y(n_282)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_274),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_228),
.C(n_225),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_241),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_275),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_239),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_273),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_259),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_241),
.C(n_234),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_283),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_282),
.B(n_289),
.Y(n_299)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_268),
.A2(n_223),
.B1(n_242),
.B2(n_230),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_284),
.A2(n_285),
.B(n_288),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_208),
.B1(n_256),
.B2(n_218),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_257),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_286),
.A2(n_280),
.B(n_278),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_257),
.A2(n_249),
.B(n_246),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_248),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_298),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_263),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_292),
.C(n_290),
.Y(n_308)
);

AO21x1_ASAP7_75t_L g293 ( 
.A1(n_278),
.A2(n_261),
.B(n_269),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_293),
.B(n_300),
.Y(n_304)
);

AND2x6_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_272),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_297),
.A2(n_301),
.B(n_287),
.Y(n_306)
);

FAx1_ASAP7_75t_SL g300 ( 
.A(n_285),
.B(n_251),
.CI(n_228),
.CON(n_300),
.SN(n_300)
);

INVxp33_ASAP7_75t_L g301 ( 
.A(n_288),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_261),
.B1(n_279),
.B2(n_270),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_302),
.A2(n_307),
.B1(n_293),
.B2(n_300),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_295),
.B(n_284),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_229),
.C(n_244),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_309),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_301),
.A2(n_297),
.B1(n_235),
.B2(n_281),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_310),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_277),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_247),
.C(n_260),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_312),
.A2(n_316),
.B(n_317),
.Y(n_321)
);

NAND4xp25_ASAP7_75t_SL g313 ( 
.A(n_305),
.B(n_299),
.C(n_265),
.D(n_271),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_314),
.C(n_12),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_303),
.B(n_265),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_10),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g318 ( 
.A1(n_315),
.A2(n_310),
.A3(n_308),
.B1(n_15),
.B2(n_16),
.C1(n_14),
.C2(n_12),
.Y(n_318)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_318),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_320),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_311),
.A2(n_12),
.B(n_14),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_322),
.A2(n_316),
.B(n_321),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_323),
.Y(n_325)
);

AOI21x1_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_15),
.B(n_313),
.Y(n_326)
);


endmodule