module real_aes_7681_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g233 ( .A1(n_0), .A2(n_234), .B(n_235), .C(n_239), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_1), .B(n_175), .Y(n_240) );
INVx1_ASAP7_75t_L g108 ( .A(n_2), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_3), .B(n_147), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_4), .A2(n_133), .B(n_138), .C(n_501), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_5), .A2(n_128), .B(n_539), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_6), .A2(n_128), .B(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_7), .B(n_175), .Y(n_545) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_8), .A2(n_163), .B(n_179), .Y(n_178) );
AND2x6_ASAP7_75t_L g133 ( .A(n_9), .B(n_134), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_10), .A2(n_133), .B(n_138), .C(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g483 ( .A(n_11), .Y(n_483) );
INVx1_ASAP7_75t_L g105 ( .A(n_12), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_12), .B(n_40), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_13), .B(n_238), .Y(n_503) );
INVx1_ASAP7_75t_L g157 ( .A(n_14), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_15), .B(n_147), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_16), .A2(n_148), .B(n_491), .C(n_493), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_17), .B(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_18), .B(n_175), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_19), .B(n_212), .Y(n_582) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_20), .A2(n_138), .B(n_189), .C(n_208), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_21), .A2(n_187), .B(n_237), .C(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_22), .B(n_238), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_23), .B(n_238), .Y(n_523) );
CKINVDCx16_ASAP7_75t_R g530 ( .A(n_24), .Y(n_530) );
INVx1_ASAP7_75t_L g522 ( .A(n_25), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_26), .A2(n_138), .B(n_182), .C(n_189), .Y(n_181) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_27), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_28), .Y(n_499) );
INVx1_ASAP7_75t_L g579 ( .A(n_29), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_30), .A2(n_128), .B(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g131 ( .A(n_31), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_32), .A2(n_136), .B(n_151), .C(n_197), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_33), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_34), .A2(n_237), .B(n_542), .C(n_544), .Y(n_541) );
INVxp67_ASAP7_75t_L g580 ( .A(n_35), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_36), .B(n_184), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_37), .A2(n_138), .B(n_189), .C(n_521), .Y(n_520) );
CKINVDCx14_ASAP7_75t_R g540 ( .A(n_38), .Y(n_540) );
AOI222xp33_ASAP7_75t_L g464 ( .A1(n_39), .A2(n_98), .B1(n_465), .B2(n_742), .C1(n_743), .C2(n_746), .Y(n_464) );
INVx1_ASAP7_75t_L g742 ( .A(n_39), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_40), .B(n_105), .Y(n_104) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_41), .A2(n_239), .B(n_481), .C(n_482), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_42), .B(n_206), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_43), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g119 ( .A1(n_44), .A2(n_120), .B1(n_121), .B2(n_451), .Y(n_119) );
INVx1_ASAP7_75t_L g451 ( .A(n_44), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_45), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_46), .B(n_128), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_47), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_48), .Y(n_576) );
A2O1A1Ixp33_ASAP7_75t_L g135 ( .A1(n_49), .A2(n_136), .B(n_141), .C(n_151), .Y(n_135) );
INVx1_ASAP7_75t_L g236 ( .A(n_50), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_51), .A2(n_100), .B1(n_113), .B2(n_750), .Y(n_99) );
INVx1_ASAP7_75t_L g142 ( .A(n_52), .Y(n_142) );
INVx1_ASAP7_75t_L g511 ( .A(n_53), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_54), .B(n_128), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_55), .Y(n_215) );
CKINVDCx14_ASAP7_75t_R g479 ( .A(n_56), .Y(n_479) );
INVx1_ASAP7_75t_L g134 ( .A(n_57), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_58), .B(n_128), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_59), .B(n_175), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g168 ( .A1(n_60), .A2(n_169), .B(n_171), .C(n_173), .Y(n_168) );
INVx1_ASAP7_75t_L g156 ( .A(n_61), .Y(n_156) );
INVx1_ASAP7_75t_SL g543 ( .A(n_62), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_63), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_64), .B(n_147), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_65), .B(n_175), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_66), .B(n_148), .Y(n_250) );
INVx1_ASAP7_75t_L g533 ( .A(n_67), .Y(n_533) );
CKINVDCx16_ASAP7_75t_R g232 ( .A(n_68), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_69), .B(n_144), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_70), .A2(n_138), .B(n_151), .C(n_221), .Y(n_220) );
CKINVDCx16_ASAP7_75t_R g167 ( .A(n_71), .Y(n_167) );
INVx1_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_73), .A2(n_128), .B(n_478), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_74), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_75), .A2(n_128), .B(n_488), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_76), .A2(n_206), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g489 ( .A(n_77), .Y(n_489) );
CKINVDCx16_ASAP7_75t_R g519 ( .A(n_78), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_79), .B(n_143), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_80), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_81), .A2(n_128), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g492 ( .A(n_82), .Y(n_492) );
INVx2_ASAP7_75t_L g154 ( .A(n_83), .Y(n_154) );
INVx1_ASAP7_75t_L g502 ( .A(n_84), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_85), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_86), .B(n_238), .Y(n_251) );
INVx2_ASAP7_75t_L g109 ( .A(n_87), .Y(n_109) );
OR2x2_ASAP7_75t_L g455 ( .A(n_87), .B(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g741 ( .A(n_87), .B(n_457), .Y(n_741) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_88), .A2(n_138), .B(n_151), .C(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_89), .B(n_128), .Y(n_195) );
INVx1_ASAP7_75t_L g198 ( .A(n_90), .Y(n_198) );
INVxp67_ASAP7_75t_L g172 ( .A(n_91), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_92), .B(n_163), .Y(n_484) );
INVx2_ASAP7_75t_L g514 ( .A(n_93), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_94), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g222 ( .A(n_95), .Y(n_222) );
INVx1_ASAP7_75t_L g246 ( .A(n_96), .Y(n_246) );
AND2x2_ASAP7_75t_L g158 ( .A(n_97), .B(n_153), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
INVx3_ASAP7_75t_SL g752 ( .A(n_102), .Y(n_752) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_106), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx14_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_109), .C(n_110), .Y(n_107) );
AND2x2_ASAP7_75t_L g457 ( .A(n_108), .B(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g470 ( .A(n_109), .B(n_457), .Y(n_470) );
NOR2x2_ASAP7_75t_L g745 ( .A(n_109), .B(n_456), .Y(n_745) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_118), .B(n_463), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g749 ( .A(n_117), .Y(n_749) );
OAI21xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_452), .B(n_459), .Y(n_118) );
AOI22x1_ASAP7_75t_SL g747 ( .A1(n_120), .A2(n_467), .B1(n_738), .B2(n_748), .Y(n_747) );
INVx4_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_121), .A2(n_467), .B1(n_471), .B2(n_738), .Y(n_466) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OR5x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_324), .C(n_402), .D(n_426), .E(n_443), .Y(n_122) );
OAI211xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_190), .B(n_241), .C(n_301), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_159), .Y(n_124) );
AND2x2_ASAP7_75t_L g255 ( .A(n_125), .B(n_161), .Y(n_255) );
INVx5_ASAP7_75t_SL g283 ( .A(n_125), .Y(n_283) );
AND2x2_ASAP7_75t_L g319 ( .A(n_125), .B(n_304), .Y(n_319) );
OR2x2_ASAP7_75t_L g358 ( .A(n_125), .B(n_160), .Y(n_358) );
OR2x2_ASAP7_75t_L g389 ( .A(n_125), .B(n_280), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_125), .B(n_293), .Y(n_425) );
AND2x2_ASAP7_75t_L g437 ( .A(n_125), .B(n_280), .Y(n_437) );
OR2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_158), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_135), .B(n_153), .Y(n_126) );
BUFx2_ASAP7_75t_L g206 ( .A(n_128), .Y(n_206) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_133), .Y(n_128) );
NAND2x1p5_ASAP7_75t_L g247 ( .A(n_129), .B(n_133), .Y(n_247) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_132), .Y(n_129) );
INVx1_ASAP7_75t_L g173 ( .A(n_130), .Y(n_173) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g139 ( .A(n_131), .Y(n_139) );
INVx1_ASAP7_75t_L g188 ( .A(n_131), .Y(n_188) );
INVx1_ASAP7_75t_L g140 ( .A(n_132), .Y(n_140) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_132), .Y(n_145) );
INVx3_ASAP7_75t_L g148 ( .A(n_132), .Y(n_148) );
INVx1_ASAP7_75t_L g184 ( .A(n_132), .Y(n_184) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_132), .Y(n_238) );
INVx4_ASAP7_75t_SL g152 ( .A(n_133), .Y(n_152) );
BUFx3_ASAP7_75t_L g189 ( .A(n_133), .Y(n_189) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
O2A1O1Ixp33_ASAP7_75t_L g166 ( .A1(n_137), .A2(n_152), .B(n_167), .C(n_168), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_SL g231 ( .A1(n_137), .A2(n_152), .B(n_232), .C(n_233), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_SL g478 ( .A1(n_137), .A2(n_152), .B(n_479), .C(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_SL g488 ( .A1(n_137), .A2(n_152), .B(n_489), .C(n_490), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_SL g510 ( .A1(n_137), .A2(n_152), .B(n_511), .C(n_512), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_137), .A2(n_152), .B(n_540), .C(n_541), .Y(n_539) );
O2A1O1Ixp33_ASAP7_75t_SL g575 ( .A1(n_137), .A2(n_152), .B(n_576), .C(n_577), .Y(n_575) );
INVx5_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x6_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
BUFx3_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_139), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_146), .C(n_149), .Y(n_141) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_143), .A2(n_149), .B(n_198), .C(n_199), .Y(n_197) );
O2A1O1Ixp5_ASAP7_75t_L g501 ( .A1(n_143), .A2(n_502), .B(n_503), .C(n_504), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_143), .A2(n_504), .B(n_533), .C(n_534), .Y(n_532) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx4_ASAP7_75t_L g170 ( .A(n_145), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_147), .B(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g234 ( .A(n_147), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_147), .A2(n_211), .B(n_522), .C(n_523), .Y(n_521) );
OAI22xp33_ASAP7_75t_L g578 ( .A1(n_147), .A2(n_170), .B1(n_579), .B2(n_580), .Y(n_578) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_148), .B(n_483), .Y(n_482) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g239 ( .A(n_150), .Y(n_239) );
INVx1_ASAP7_75t_L g493 ( .A(n_150), .Y(n_493) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_153), .A2(n_195), .B(n_196), .Y(n_194) );
INVx2_ASAP7_75t_L g213 ( .A(n_153), .Y(n_213) );
INVx1_ASAP7_75t_L g216 ( .A(n_153), .Y(n_216) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_153), .A2(n_477), .B(n_484), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_153), .A2(n_247), .B(n_519), .C(n_520), .Y(n_518) );
AND2x2_ASAP7_75t_SL g153 ( .A(n_154), .B(n_155), .Y(n_153) );
AND2x2_ASAP7_75t_L g164 ( .A(n_154), .B(n_155), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
AND2x2_ASAP7_75t_L g436 ( .A(n_159), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
OR2x2_ASAP7_75t_L g299 ( .A(n_160), .B(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_177), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_161), .B(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_161), .Y(n_292) );
INVx3_ASAP7_75t_L g307 ( .A(n_161), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_161), .B(n_177), .Y(n_331) );
OR2x2_ASAP7_75t_L g340 ( .A(n_161), .B(n_283), .Y(n_340) );
AND2x2_ASAP7_75t_L g344 ( .A(n_161), .B(n_304), .Y(n_344) );
AND2x2_ASAP7_75t_L g350 ( .A(n_161), .B(n_351), .Y(n_350) );
INVxp67_ASAP7_75t_L g387 ( .A(n_161), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_161), .B(n_244), .Y(n_401) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_165), .B(n_174), .Y(n_161) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_162), .A2(n_487), .B(n_494), .Y(n_486) );
OA21x2_ASAP7_75t_L g508 ( .A1(n_162), .A2(n_509), .B(n_515), .Y(n_508) );
OA21x2_ASAP7_75t_L g537 ( .A1(n_162), .A2(n_538), .B(n_545), .Y(n_537) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx4_ASAP7_75t_L g176 ( .A(n_163), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_163), .A2(n_180), .B(n_181), .Y(n_179) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g254 ( .A(n_164), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_169), .A2(n_222), .B(n_223), .C(n_224), .Y(n_221) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_170), .B(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_170), .B(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g211 ( .A(n_173), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_173), .B(n_578), .Y(n_577) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_175), .A2(n_230), .B(n_240), .Y(n_229) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_176), .B(n_201), .Y(n_200) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_176), .A2(n_219), .B(n_227), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_176), .B(n_228), .Y(n_227) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_176), .A2(n_245), .B(n_252), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_176), .B(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_176), .B(n_525), .Y(n_524) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_176), .A2(n_529), .B(n_535), .Y(n_528) );
OR2x2_ASAP7_75t_L g293 ( .A(n_177), .B(n_244), .Y(n_293) );
AND2x2_ASAP7_75t_L g304 ( .A(n_177), .B(n_280), .Y(n_304) );
AND2x2_ASAP7_75t_L g316 ( .A(n_177), .B(n_307), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g339 ( .A(n_177), .B(n_244), .Y(n_339) );
INVx1_ASAP7_75t_SL g351 ( .A(n_177), .Y(n_351) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g243 ( .A(n_178), .B(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_178), .B(n_283), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_185), .B(n_186), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_186), .A2(n_250), .B(n_251), .Y(n_249) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_202), .Y(n_191) );
AND2x2_ASAP7_75t_L g264 ( .A(n_192), .B(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_192), .B(n_217), .Y(n_268) );
AND2x2_ASAP7_75t_L g271 ( .A(n_192), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_192), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g296 ( .A(n_192), .B(n_287), .Y(n_296) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_192), .Y(n_315) );
AND2x2_ASAP7_75t_L g336 ( .A(n_192), .B(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g346 ( .A(n_192), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g392 ( .A(n_192), .B(n_275), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_192), .B(n_298), .Y(n_419) );
INVx5_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
BUFx2_ASAP7_75t_L g289 ( .A(n_193), .Y(n_289) );
AND2x2_ASAP7_75t_L g355 ( .A(n_193), .B(n_287), .Y(n_355) );
AND2x2_ASAP7_75t_L g439 ( .A(n_193), .B(n_307), .Y(n_439) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_200), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_202), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g428 ( .A(n_202), .Y(n_428) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_217), .Y(n_202) );
AND2x2_ASAP7_75t_L g258 ( .A(n_203), .B(n_259), .Y(n_258) );
AND2x4_ASAP7_75t_L g267 ( .A(n_203), .B(n_265), .Y(n_267) );
INVx5_ASAP7_75t_L g275 ( .A(n_203), .Y(n_275) );
AND2x2_ASAP7_75t_L g298 ( .A(n_203), .B(n_229), .Y(n_298) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_203), .Y(n_335) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_214), .Y(n_203) );
AOI21xp5_ASAP7_75t_SL g204 ( .A1(n_205), .A2(n_207), .B(n_212), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_211), .Y(n_208) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_213), .B(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_216), .A2(n_498), .B(n_505), .Y(n_497) );
INVx1_ASAP7_75t_L g376 ( .A(n_217), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_217), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g409 ( .A(n_217), .B(n_275), .Y(n_409) );
A2O1A1Ixp33_ASAP7_75t_L g438 ( .A1(n_217), .A2(n_332), .B(n_439), .C(n_440), .Y(n_438) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_229), .Y(n_217) );
BUFx2_ASAP7_75t_L g259 ( .A(n_218), .Y(n_259) );
INVx2_ASAP7_75t_L g263 ( .A(n_218), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_226), .Y(n_219) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx3_ASAP7_75t_L g544 ( .A(n_225), .Y(n_544) );
INVx2_ASAP7_75t_L g265 ( .A(n_229), .Y(n_265) );
AND2x2_ASAP7_75t_L g272 ( .A(n_229), .B(n_263), .Y(n_272) );
AND2x2_ASAP7_75t_L g363 ( .A(n_229), .B(n_275), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_237), .B(n_543), .Y(n_542) );
INVx4_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g481 ( .A(n_238), .Y(n_481) );
INVx2_ASAP7_75t_L g504 ( .A(n_239), .Y(n_504) );
AOI211x1_ASAP7_75t_SL g241 ( .A1(n_242), .A2(n_256), .B(n_269), .C(n_294), .Y(n_241) );
INVx1_ASAP7_75t_L g360 ( .A(n_242), .Y(n_360) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_255), .Y(n_242) );
INVx5_ASAP7_75t_SL g280 ( .A(n_244), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_244), .B(n_350), .Y(n_349) );
AOI311xp33_ASAP7_75t_L g368 ( .A1(n_244), .A2(n_369), .A3(n_371), .B(n_372), .C(n_378), .Y(n_368) );
A2O1A1Ixp33_ASAP7_75t_L g403 ( .A1(n_244), .A2(n_316), .B(n_404), .C(n_407), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_247), .B(n_248), .Y(n_245) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_247), .A2(n_499), .B(n_500), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g529 ( .A1(n_247), .A2(n_530), .B(n_531), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
INVx2_ASAP7_75t_L g572 ( .A(n_254), .Y(n_572) );
INVxp67_ASAP7_75t_L g323 ( .A(n_255), .Y(n_323) );
NAND4xp25_ASAP7_75t_SL g256 ( .A(n_257), .B(n_260), .C(n_266), .D(n_268), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_257), .B(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g314 ( .A(n_258), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_264), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_261), .B(n_267), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_261), .B(n_274), .Y(n_394) );
BUFx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_262), .B(n_275), .Y(n_412) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g287 ( .A(n_263), .Y(n_287) );
INVxp67_ASAP7_75t_L g322 ( .A(n_264), .Y(n_322) );
AND2x4_ASAP7_75t_L g274 ( .A(n_265), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g348 ( .A(n_265), .B(n_287), .Y(n_348) );
INVx1_ASAP7_75t_L g375 ( .A(n_265), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_265), .B(n_362), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_266), .B(n_336), .Y(n_356) );
INVx1_ASAP7_75t_SL g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_267), .B(n_289), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_267), .B(n_336), .Y(n_435) );
INVx1_ASAP7_75t_L g446 ( .A(n_268), .Y(n_446) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_273), .B(n_276), .C(n_284), .Y(n_269) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g288 ( .A(n_272), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g326 ( .A(n_272), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g308 ( .A(n_273), .Y(n_308) );
AND2x2_ASAP7_75t_L g285 ( .A(n_274), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_274), .B(n_336), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_274), .B(n_355), .Y(n_379) );
OR2x2_ASAP7_75t_L g295 ( .A(n_275), .B(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g327 ( .A(n_275), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_275), .B(n_287), .Y(n_342) );
AND2x2_ASAP7_75t_L g399 ( .A(n_275), .B(n_355), .Y(n_399) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_275), .Y(n_406) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_277), .A2(n_289), .B1(n_411), .B2(n_413), .C(n_416), .Y(n_410) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_281), .Y(n_277) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g300 ( .A(n_280), .B(n_283), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_280), .B(n_350), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_280), .B(n_307), .Y(n_415) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g400 ( .A(n_282), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g414 ( .A(n_282), .B(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_283), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g311 ( .A(n_283), .B(n_304), .Y(n_311) );
AND2x2_ASAP7_75t_L g381 ( .A(n_283), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_283), .B(n_330), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_283), .B(n_431), .Y(n_430) );
OAI21xp5_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_288), .B(n_290), .Y(n_284) );
INVx2_ASAP7_75t_L g317 ( .A(n_285), .Y(n_317) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g337 ( .A(n_287), .Y(n_337) );
OR2x2_ASAP7_75t_L g341 ( .A(n_289), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g444 ( .A(n_289), .B(n_412), .Y(n_444) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AOI21xp33_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_297), .B(n_299), .Y(n_294) );
INVx1_ASAP7_75t_L g448 ( .A(n_295), .Y(n_448) );
INVx2_ASAP7_75t_SL g362 ( .A(n_296), .Y(n_362) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_L g443 ( .A1(n_299), .A2(n_380), .B(n_444), .C(n_445), .Y(n_443) );
OAI322xp33_ASAP7_75t_SL g312 ( .A1(n_300), .A2(n_313), .A3(n_316), .B1(n_317), .B2(n_318), .C1(n_320), .C2(n_323), .Y(n_312) );
INVx2_ASAP7_75t_L g332 ( .A(n_300), .Y(n_332) );
AOI221xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_308), .B1(n_309), .B2(n_311), .C(n_312), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI22xp33_ASAP7_75t_SL g378 ( .A1(n_303), .A2(n_379), .B1(n_380), .B2(n_383), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_304), .B(n_307), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_304), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g377 ( .A(n_306), .B(n_339), .Y(n_377) );
INVx1_ASAP7_75t_L g367 ( .A(n_307), .Y(n_367) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_311), .A2(n_421), .B(n_423), .Y(n_420) );
AOI21xp33_ASAP7_75t_L g345 ( .A1(n_313), .A2(n_346), .B(n_349), .Y(n_345) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NOR2xp67_ASAP7_75t_SL g374 ( .A(n_315), .B(n_375), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_315), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g431 ( .A(n_316), .Y(n_431) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND4xp25_ASAP7_75t_L g324 ( .A(n_325), .B(n_352), .C(n_368), .D(n_384), .Y(n_324) );
AOI211xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_328), .B(n_333), .C(n_345), .Y(n_325) );
INVx1_ASAP7_75t_L g417 ( .A(n_326), .Y(n_417) );
AND2x2_ASAP7_75t_L g365 ( .A(n_327), .B(n_348), .Y(n_365) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_332), .B(n_367), .Y(n_366) );
OAI22xp33_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_338), .B1(n_341), .B2(n_343), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_335), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g383 ( .A(n_336), .Y(n_383) );
O2A1O1Ixp33_ASAP7_75t_L g397 ( .A1(n_336), .A2(n_375), .B(n_398), .C(n_400), .Y(n_397) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx1_ASAP7_75t_L g382 ( .A(n_339), .Y(n_382) );
INVx1_ASAP7_75t_L g442 ( .A(n_340), .Y(n_442) );
NAND2xp33_ASAP7_75t_SL g432 ( .A(n_341), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g371 ( .A(n_350), .Y(n_371) );
O2A1O1Ixp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_356), .B(n_357), .C(n_359), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_361), .B1(n_364), .B2(n_366), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_362), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_367), .B(n_388), .Y(n_450) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AOI21xp33_ASAP7_75t_SL g372 ( .A1(n_373), .A2(n_376), .B(n_377), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
AOI221xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_390), .B1(n_393), .B2(n_395), .C(n_397), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_400), .A2(n_417), .B1(n_418), .B2(n_419), .Y(n_416) );
NAND3xp33_ASAP7_75t_SL g402 ( .A(n_403), .B(n_410), .C(n_420), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
CKINVDCx16_ASAP7_75t_R g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVxp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI211xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B(n_429), .C(n_438), .Y(n_426) );
INVx1_ASAP7_75t_L g447 ( .A(n_427), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_432), .B1(n_434), .B2(n_436), .Y(n_429) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B1(n_448), .B2(n_449), .Y(n_445) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g462 ( .A(n_455), .Y(n_462) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND3xp33_ASAP7_75t_L g463 ( .A(n_459), .B(n_464), .C(n_749), .Y(n_463) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g748 ( .A(n_471), .Y(n_748) );
OR2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_668), .Y(n_471) );
NAND5xp2_ASAP7_75t_L g472 ( .A(n_473), .B(n_583), .C(n_615), .D(n_632), .E(n_655), .Y(n_472) );
AOI221xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_516), .B1(n_546), .B2(n_550), .C(n_554), .Y(n_473) );
INVx1_ASAP7_75t_L g695 ( .A(n_474), .Y(n_695) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_495), .Y(n_474) );
AND3x2_ASAP7_75t_L g670 ( .A(n_475), .B(n_497), .C(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_485), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_476), .B(n_552), .Y(n_551) );
BUFx3_ASAP7_75t_L g561 ( .A(n_476), .Y(n_561) );
AND2x2_ASAP7_75t_L g565 ( .A(n_476), .B(n_507), .Y(n_565) );
INVx2_ASAP7_75t_L g592 ( .A(n_476), .Y(n_592) );
OR2x2_ASAP7_75t_L g603 ( .A(n_476), .B(n_508), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_476), .B(n_496), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_476), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g682 ( .A(n_476), .B(n_508), .Y(n_682) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_485), .Y(n_564) );
AND2x2_ASAP7_75t_L g623 ( .A(n_485), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_485), .B(n_496), .Y(n_642) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
OR2x2_ASAP7_75t_L g553 ( .A(n_486), .B(n_496), .Y(n_553) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_486), .Y(n_560) );
AND2x2_ASAP7_75t_L g609 ( .A(n_486), .B(n_508), .Y(n_609) );
NAND3xp33_ASAP7_75t_L g634 ( .A(n_486), .B(n_495), .C(n_592), .Y(n_634) );
AND2x2_ASAP7_75t_L g699 ( .A(n_486), .B(n_497), .Y(n_699) );
AND2x2_ASAP7_75t_L g733 ( .A(n_486), .B(n_496), .Y(n_733) );
INVxp67_ASAP7_75t_L g562 ( .A(n_495), .Y(n_562) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_507), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_496), .B(n_592), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_496), .B(n_623), .Y(n_631) );
AND2x2_ASAP7_75t_L g681 ( .A(n_496), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g709 ( .A(n_496), .Y(n_709) );
INVx4_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g616 ( .A(n_497), .B(n_609), .Y(n_616) );
BUFx3_ASAP7_75t_L g648 ( .A(n_497), .Y(n_648) );
INVx2_ASAP7_75t_L g624 ( .A(n_507), .Y(n_624) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_508), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_516), .A2(n_684), .B1(n_686), .B2(n_687), .Y(n_683) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_526), .Y(n_516) );
AND2x2_ASAP7_75t_L g546 ( .A(n_517), .B(n_547), .Y(n_546) );
INVx3_ASAP7_75t_SL g557 ( .A(n_517), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_517), .B(n_587), .Y(n_619) );
OR2x2_ASAP7_75t_L g638 ( .A(n_517), .B(n_527), .Y(n_638) );
AND2x2_ASAP7_75t_L g643 ( .A(n_517), .B(n_595), .Y(n_643) );
AND2x2_ASAP7_75t_L g646 ( .A(n_517), .B(n_588), .Y(n_646) );
AND2x2_ASAP7_75t_L g658 ( .A(n_517), .B(n_537), .Y(n_658) );
AND2x2_ASAP7_75t_L g674 ( .A(n_517), .B(n_528), .Y(n_674) );
AND2x4_ASAP7_75t_L g677 ( .A(n_517), .B(n_548), .Y(n_677) );
OR2x2_ASAP7_75t_L g694 ( .A(n_517), .B(n_630), .Y(n_694) );
OR2x2_ASAP7_75t_L g725 ( .A(n_517), .B(n_570), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g727 ( .A(n_517), .B(n_653), .Y(n_727) );
OR2x6_ASAP7_75t_L g517 ( .A(n_518), .B(n_524), .Y(n_517) );
AND2x2_ASAP7_75t_L g601 ( .A(n_526), .B(n_568), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_526), .B(n_588), .Y(n_720) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_537), .Y(n_526) );
AND2x2_ASAP7_75t_L g556 ( .A(n_527), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g587 ( .A(n_527), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g595 ( .A(n_527), .B(n_570), .Y(n_595) );
AND2x2_ASAP7_75t_L g613 ( .A(n_527), .B(n_548), .Y(n_613) );
OR2x2_ASAP7_75t_L g630 ( .A(n_527), .B(n_588), .Y(n_630) );
INVx2_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
BUFx2_ASAP7_75t_L g549 ( .A(n_528), .Y(n_549) );
AND2x2_ASAP7_75t_L g653 ( .A(n_528), .B(n_537), .Y(n_653) );
INVx2_ASAP7_75t_L g548 ( .A(n_537), .Y(n_548) );
INVx1_ASAP7_75t_L g665 ( .A(n_537), .Y(n_665) );
AND2x2_ASAP7_75t_L g715 ( .A(n_537), .B(n_557), .Y(n_715) );
AND2x2_ASAP7_75t_L g567 ( .A(n_547), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g599 ( .A(n_547), .B(n_557), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_547), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
AND2x2_ASAP7_75t_L g586 ( .A(n_548), .B(n_557), .Y(n_586) );
OR2x2_ASAP7_75t_L g702 ( .A(n_549), .B(n_676), .Y(n_702) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_552), .B(n_682), .Y(n_688) );
INVx2_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
OAI32xp33_ASAP7_75t_L g644 ( .A1(n_553), .A2(n_645), .A3(n_647), .B1(n_649), .B2(n_650), .Y(n_644) );
OR2x2_ASAP7_75t_L g661 ( .A(n_553), .B(n_603), .Y(n_661) );
OAI21xp33_ASAP7_75t_SL g686 ( .A1(n_553), .A2(n_563), .B(n_591), .Y(n_686) );
OAI22xp33_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_558), .B1(n_563), .B2(n_566), .Y(n_554) );
INVxp33_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_556), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_557), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g612 ( .A(n_557), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g712 ( .A(n_557), .B(n_653), .Y(n_712) );
OR2x2_ASAP7_75t_L g736 ( .A(n_557), .B(n_630), .Y(n_736) );
AOI21xp33_ASAP7_75t_L g719 ( .A1(n_558), .A2(n_618), .B(n_720), .Y(n_719) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_562), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g596 ( .A(n_560), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_560), .B(n_565), .Y(n_614) );
AND2x2_ASAP7_75t_L g636 ( .A(n_561), .B(n_609), .Y(n_636) );
INVx1_ASAP7_75t_L g649 ( .A(n_561), .Y(n_649) );
OR2x2_ASAP7_75t_L g654 ( .A(n_561), .B(n_588), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_564), .B(n_603), .Y(n_602) );
OAI22xp33_ASAP7_75t_L g584 ( .A1(n_565), .A2(n_585), .B1(n_590), .B2(n_594), .Y(n_584) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_568), .A2(n_627), .B1(n_634), .B2(n_635), .Y(n_633) );
AND2x2_ASAP7_75t_L g711 ( .A(n_568), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_570), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g730 ( .A(n_570), .B(n_613), .Y(n_730) );
AO21x2_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_573), .B(n_581), .Y(n_570) );
INVx1_ASAP7_75t_L g589 ( .A(n_571), .Y(n_589) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OA21x2_ASAP7_75t_L g588 ( .A1(n_574), .A2(n_582), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AOI221xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_596), .B1(n_597), .B2(n_602), .C(n_604), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_586), .B(n_588), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_586), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g605 ( .A(n_587), .Y(n_605) );
O2A1O1Ixp33_ASAP7_75t_L g692 ( .A1(n_587), .A2(n_693), .B(n_694), .C(n_695), .Y(n_692) );
AND2x2_ASAP7_75t_L g697 ( .A(n_587), .B(n_677), .Y(n_697) );
O2A1O1Ixp33_ASAP7_75t_SL g735 ( .A1(n_587), .A2(n_676), .B(n_736), .C(n_737), .Y(n_735) );
BUFx3_ASAP7_75t_L g627 ( .A(n_588), .Y(n_627) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_591), .B(n_648), .Y(n_691) );
AOI211xp5_ASAP7_75t_L g710 ( .A1(n_591), .A2(n_711), .B(n_713), .C(n_719), .Y(n_710) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVxp67_ASAP7_75t_L g671 ( .A(n_593), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_595), .B(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_598), .B(n_600), .Y(n_597) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
AOI211xp5_ASAP7_75t_L g615 ( .A1(n_599), .A2(n_616), .B(n_617), .C(n_625), .Y(n_615) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g700 ( .A(n_603), .Y(n_700) );
OR2x2_ASAP7_75t_L g717 ( .A(n_603), .B(n_647), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_606), .B1(n_611), .B2(n_614), .Y(n_604) );
OAI22xp33_ASAP7_75t_L g617 ( .A1(n_606), .A2(n_618), .B1(n_619), .B2(n_620), .Y(n_617) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
OR2x2_ASAP7_75t_L g704 ( .A(n_608), .B(n_648), .Y(n_704) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g659 ( .A(n_609), .B(n_649), .Y(n_659) );
INVx1_ASAP7_75t_L g667 ( .A(n_610), .Y(n_667) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_613), .B(n_627), .Y(n_675) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_623), .B(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g732 ( .A(n_624), .Y(n_732) );
AOI21xp33_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_628), .B(n_631), .Y(n_625) );
INVx1_ASAP7_75t_L g662 ( .A(n_626), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_627), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_627), .B(n_658), .Y(n_657) );
NAND2x1p5_ASAP7_75t_L g678 ( .A(n_627), .B(n_653), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_627), .B(n_674), .Y(n_685) );
OAI211xp5_ASAP7_75t_L g689 ( .A1(n_627), .A2(n_637), .B(n_677), .C(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
AOI221xp5_ASAP7_75t_SL g632 ( .A1(n_633), .A2(n_637), .B1(n_639), .B2(n_643), .C(n_644), .Y(n_632) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVxp67_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_641), .B(n_649), .Y(n_723) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
O2A1O1Ixp33_ASAP7_75t_L g734 ( .A1(n_643), .A2(n_658), .B(n_660), .C(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_646), .B(n_653), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g737 ( .A(n_647), .B(n_700), .Y(n_737) );
CKINVDCx16_ASAP7_75t_R g647 ( .A(n_648), .Y(n_647) );
INVxp33_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
AOI21xp33_ASAP7_75t_SL g663 ( .A1(n_652), .A2(n_664), .B(n_666), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_652), .B(n_725), .Y(n_724) );
INVx2_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_653), .B(n_707), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_659), .B1(n_660), .B2(n_662), .C(n_663), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_659), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g693 ( .A(n_665), .Y(n_693) );
NAND5xp2_ASAP7_75t_L g668 ( .A(n_669), .B(n_696), .C(n_710), .D(n_721), .E(n_734), .Y(n_668) );
AOI211xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_672), .B(n_679), .C(n_692), .Y(n_669) );
INVx2_ASAP7_75t_SL g716 ( .A(n_670), .Y(n_716) );
NAND4xp25_ASAP7_75t_SL g672 ( .A(n_673), .B(n_675), .C(n_676), .D(n_678), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx3_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI211xp5_ASAP7_75t_SL g679 ( .A1(n_678), .A2(n_680), .B(n_683), .C(n_689), .Y(n_679) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_681), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_681), .A2(n_722), .B1(n_724), .B2(n_726), .C(n_728), .Y(n_721) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI221xp5_ASAP7_75t_SL g696 ( .A1(n_697), .A2(n_698), .B1(n_701), .B2(n_703), .C(n_705), .Y(n_696) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_704), .A2(n_727), .B1(n_729), .B2(n_731), .Y(n_728) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_713) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_752), .Y(n_751) );
endmodule