module fake_jpeg_16846_n_317 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_16),
.B(n_7),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_31),
.B(n_34),
.Y(n_52)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_7),
.B(n_12),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_37),
.Y(n_46)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_16),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_32),
.A2(n_15),
.B1(n_18),
.B2(n_25),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_25),
.B(n_23),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_32),
.A2(n_18),
.B1(n_15),
.B2(n_26),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_26),
.B1(n_23),
.B2(n_30),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_29),
.B(n_33),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_18),
.B1(n_21),
.B2(n_17),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_25),
.B1(n_23),
.B2(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_51),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_14),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_30),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_20),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_49),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_35),
.B1(n_18),
.B2(n_30),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_69),
.B1(n_47),
.B2(n_51),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_57),
.A2(n_77),
.B(n_42),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_52),
.B(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_60),
.A2(n_65),
.B1(n_68),
.B2(n_74),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_72),
.Y(n_90)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_37),
.B1(n_36),
.B2(n_21),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_37),
.B1(n_36),
.B2(n_17),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

BUFx2_ASAP7_75t_SL g71 ( 
.A(n_51),
.Y(n_71)
);

BUFx2_ASAP7_75t_SL g91 ( 
.A(n_71),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_28),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_39),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_27),
.B1(n_36),
.B2(n_37),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_28),
.B1(n_14),
.B2(n_17),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_41),
.B1(n_40),
.B2(n_45),
.Y(n_93)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_47),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_42),
.A2(n_28),
.B(n_14),
.C(n_22),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_40),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_85),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_49),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_72),
.B(n_56),
.Y(n_112)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_96),
.B1(n_65),
.B2(n_76),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_67),
.B(n_46),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_100),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_39),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_103),
.Y(n_117)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_44),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_83),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_77),
.C(n_69),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_120),
.C(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_90),
.B(n_63),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_88),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_111),
.A2(n_113),
.B1(n_125),
.B2(n_79),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_112),
.B(n_95),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_68),
.B1(n_74),
.B2(n_57),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_99),
.A2(n_68),
.B1(n_40),
.B2(n_57),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_127),
.B1(n_86),
.B2(n_91),
.Y(n_133)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_46),
.C(n_58),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_88),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_103),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_73),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_82),
.B(n_75),
.Y(n_146)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_60),
.B1(n_78),
.B2(n_50),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_91),
.A2(n_50),
.B1(n_78),
.B2(n_51),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_46),
.C(n_75),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_131),
.B(n_139),
.Y(n_158)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_133),
.A2(n_136),
.B1(n_123),
.B2(n_119),
.Y(n_167)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_149),
.B1(n_155),
.B2(n_156),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_104),
.B1(n_93),
.B2(n_83),
.Y(n_136)
);

INVxp67_ASAP7_75t_SL g137 ( 
.A(n_114),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_80),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_128),
.Y(n_168)
);

XOR2x1_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_85),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_141),
.A2(n_142),
.B(n_146),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_82),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_144),
.B(n_147),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_60),
.B1(n_85),
.B2(n_87),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_145),
.A2(n_151),
.B1(n_109),
.B2(n_108),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_110),
.B(n_87),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_86),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_148),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_87),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_129),
.A2(n_85),
.B1(n_39),
.B2(n_86),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_79),
.Y(n_152)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_135),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_159),
.B(n_160),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_108),
.C(n_109),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_171),
.C(n_173),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_135),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_163),
.B(n_164),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_138),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_155),
.A2(n_125),
.B1(n_113),
.B2(n_115),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_166),
.A2(n_167),
.B1(n_170),
.B2(n_176),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_101),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_136),
.A2(n_107),
.B1(n_128),
.B2(n_123),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_107),
.C(n_123),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_138),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_178),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_140),
.C(n_141),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_133),
.A2(n_141),
.B1(n_152),
.B2(n_154),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_130),
.A2(n_132),
.B1(n_139),
.B2(n_148),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_134),
.B1(n_47),
.B2(n_44),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_153),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_66),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_146),
.C(n_145),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_142),
.Y(n_187)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_193),
.C(n_197),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_166),
.B1(n_175),
.B2(n_165),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_195),
.B1(n_185),
.B2(n_184),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_142),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_SL g222 ( 
.A(n_192),
.B(n_199),
.C(n_205),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_151),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_157),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_202),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_131),
.B1(n_147),
.B2(n_106),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_106),
.C(n_144),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_105),
.C(n_126),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_210),
.C(n_24),
.Y(n_231)
);

A2O1A1Ixp33_ASAP7_75t_SL g199 ( 
.A1(n_167),
.A2(n_176),
.B(n_179),
.C(n_161),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_182),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_203),
.B(n_172),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_134),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_206),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_124),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_163),
.A2(n_101),
.B(n_118),
.C(n_121),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_160),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_97),
.C(n_84),
.Y(n_210)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_180),
.Y(n_214)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_170),
.B1(n_178),
.B2(n_164),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_217),
.A2(n_218),
.B1(n_220),
.B2(n_228),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_183),
.B1(n_185),
.B2(n_181),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_224),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_174),
.B1(n_97),
.B2(n_2),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_187),
.B(n_94),
.Y(n_223)
);

AOI21xp33_ASAP7_75t_L g251 ( 
.A1(n_223),
.A2(n_8),
.B(n_13),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_94),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_22),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_227),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_193),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_199),
.A2(n_10),
.B(n_13),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_199),
.A2(n_198),
.B1(n_197),
.B2(n_205),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_22),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_186),
.Y(n_230)
);

INVx11_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_188),
.C(n_211),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_24),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_213),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_240),
.C(n_242),
.Y(n_258)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_188),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_195),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_249),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_211),
.C(n_200),
.Y(n_242)
);

AOI21x1_ASAP7_75t_L g243 ( 
.A1(n_222),
.A2(n_199),
.B(n_206),
.Y(n_243)
);

NAND2xp33_ASAP7_75t_SL g264 ( 
.A(n_243),
.B(n_249),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_221),
.C(n_227),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_245),
.C(n_246),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_200),
.C(n_207),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_196),
.C(n_21),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_17),
.B(n_14),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_21),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_251),
.A2(n_8),
.B(n_13),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_248),
.A2(n_215),
.B1(n_226),
.B2(n_233),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_253),
.B(n_255),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_257),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_250),
.A2(n_217),
.B1(n_218),
.B2(n_228),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_234),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_261),
.B1(n_264),
.B2(n_265),
.Y(n_273)
);

BUFx24_ASAP7_75t_SL g257 ( 
.A(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_220),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_246),
.Y(n_271)
);

BUFx4f_ASAP7_75t_SL g261 ( 
.A(n_252),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_233),
.B1(n_9),
.B2(n_2),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_247),
.Y(n_277)
);

OAI321xp33_ASAP7_75t_L g274 ( 
.A1(n_266),
.A2(n_265),
.A3(n_261),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_262),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_278),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_235),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_7),
.Y(n_292)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_274),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_267),
.A2(n_235),
.B(n_261),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_277),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_238),
.C(n_244),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_279),
.C(n_14),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_267),
.A2(n_236),
.B(n_240),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_236),
.C(n_20),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_20),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_280),
.B(n_14),
.Y(n_281)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_281),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_292),
.C(n_20),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_270),
.Y(n_285)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_285),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_268),
.A2(n_7),
.B(n_13),
.Y(n_287)
);

A2O1A1Ixp33_ASAP7_75t_SL g297 ( 
.A1(n_287),
.A2(n_5),
.B(n_11),
.C(n_3),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_20),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_288),
.B(n_290),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_20),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_279),
.B(n_272),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_3),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_286),
.B1(n_284),
.B2(n_282),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_293),
.A2(n_298),
.B1(n_4),
.B2(n_5),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_292),
.A2(n_6),
.B(n_12),
.Y(n_294)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_294),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_287),
.A2(n_6),
.B(n_11),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

OAI321xp33_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_295),
.A3(n_0),
.B1(n_1),
.B2(n_5),
.C(n_10),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_299),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_301),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_304),
.A2(n_306),
.B(n_308),
.Y(n_313)
);

NOR3xp33_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_4),
.C(n_10),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_309),
.A2(n_297),
.B(n_1),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_305),
.A2(n_300),
.B(n_297),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_312),
.C(n_307),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_311),
.A2(n_0),
.B1(n_1),
.B2(n_313),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_10),
.B(n_0),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_314),
.B(n_315),
.C(n_1),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_316),
.Y(n_317)
);


endmodule