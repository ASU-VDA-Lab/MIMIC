module fake_jpeg_28498_n_309 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_309);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_40),
.B(n_48),
.Y(n_74)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_16),
.B(n_14),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_54),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_24),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_36),
.B1(n_28),
.B2(n_22),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_60),
.A2(n_63),
.B1(n_65),
.B2(n_76),
.Y(n_126)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_36),
.B1(n_18),
.B2(n_22),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_29),
.B(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_73),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_36),
.B1(n_35),
.B2(n_25),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_23),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_66),
.B(n_83),
.Y(n_118)
);

CKINVDCx6p67_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_35),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_75),
.B(n_81),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_39),
.A2(n_36),
.B1(n_18),
.B2(n_22),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_87),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_45),
.A2(n_52),
.B1(n_35),
.B2(n_25),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_79),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_43),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_17),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_16),
.B1(n_34),
.B2(n_33),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_104),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_19),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_58),
.A2(n_29),
.B1(n_21),
.B2(n_33),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_88),
.A2(n_95),
.B1(n_101),
.B2(n_1),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_40),
.B(n_19),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_91),
.Y(n_131)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_40),
.B(n_34),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_102),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_58),
.A2(n_21),
.B1(n_27),
.B2(n_23),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_31),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_37),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_58),
.A2(n_27),
.B1(n_17),
.B2(n_37),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_40),
.B(n_31),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_40),
.B(n_8),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_10),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_54),
.B(n_37),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_105),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_106),
.B(n_9),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_24),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_114),
.Y(n_140)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_109),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_70),
.A2(n_24),
.B1(n_13),
.B2(n_11),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_113),
.A2(n_132),
.B1(n_65),
.B2(n_97),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_0),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_1),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_81),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_59),
.A2(n_74),
.B(n_84),
.C(n_81),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_116),
.B(n_2),
.Y(n_167)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_75),
.A2(n_13),
.B(n_11),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_135),
.C(n_69),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_122),
.A2(n_67),
.B1(n_77),
.B2(n_100),
.Y(n_142)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_130),
.Y(n_143)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_71),
.B(n_1),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_127),
.A2(n_93),
.B1(n_70),
.B2(n_97),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_137),
.A2(n_139),
.B1(n_159),
.B2(n_105),
.Y(n_181)
);

AO21x1_ASAP7_75t_L g201 ( 
.A1(n_142),
.A2(n_163),
.B(n_167),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_145),
.B(n_148),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_77),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_147),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_82),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_82),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_153),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_L g150 ( 
.A1(n_107),
.A2(n_67),
.B(n_8),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_150),
.B(n_154),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_86),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_86),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_118),
.B(n_8),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_96),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_162),
.Y(n_176)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_67),
.C(n_80),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_6),
.C(n_165),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_93),
.B1(n_96),
.B2(n_90),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_157),
.A2(n_160),
.B1(n_149),
.B2(n_153),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_132),
.A2(n_130),
.B1(n_126),
.B2(n_127),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_135),
.B1(n_116),
.B2(n_112),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_90),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_111),
.A2(n_69),
.B1(n_62),
.B2(n_80),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_165),
.B(n_135),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_62),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_119),
.B(n_2),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_169),
.B(n_171),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_121),
.B(n_2),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_197),
.C(n_193),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_134),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_175),
.B(n_199),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_128),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_179),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_160),
.B(n_128),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_178),
.B(n_193),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_129),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_110),
.B(n_109),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_180),
.A2(n_194),
.B(n_198),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_181),
.A2(n_184),
.B1(n_186),
.B2(n_168),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_139),
.A2(n_124),
.B1(n_136),
.B2(n_92),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_117),
.B1(n_110),
.B2(n_5),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_187),
.A2(n_195),
.B1(n_161),
.B2(n_158),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_3),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_191),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_4),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_138),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_140),
.B(n_4),
.Y(n_191)
);

OAI21x1_ASAP7_75t_SL g194 ( 
.A1(n_156),
.A2(n_6),
.B(n_167),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_144),
.Y(n_196)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_156),
.B(n_140),
.C(n_143),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_171),
.A2(n_148),
.B(n_154),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_161),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_144),
.Y(n_200)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_168),
.B(n_141),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_202),
.A2(n_177),
.B(n_203),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_152),
.B(n_170),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_204),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_170),
.B(n_164),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_205),
.A2(n_206),
.B1(n_211),
.B2(n_228),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_201),
.A2(n_158),
.B1(n_161),
.B2(n_138),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_208),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_204),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_202),
.B(n_189),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_195),
.B1(n_181),
.B2(n_194),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_225),
.C(n_182),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_190),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_216),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_190),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_188),
.B(n_174),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_173),
.Y(n_232)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_224),
.A2(n_229),
.B(n_189),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_172),
.C(n_178),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_179),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_226),
.B(n_185),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_184),
.A2(n_173),
.B1(n_176),
.B2(n_174),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_176),
.A2(n_192),
.B(n_201),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_239),
.C(n_248),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_223),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_231),
.B(n_242),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_232),
.B(n_244),
.Y(n_253)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_182),
.C(n_191),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_243),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_205),
.A2(n_201),
.B1(n_187),
.B2(n_183),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_241),
.A2(n_235),
.B1(n_236),
.B2(n_207),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_223),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_214),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_247),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_183),
.C(n_198),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_226),
.Y(n_255)
);

XOR2x1_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_185),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_250),
.B(n_218),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_255),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_234),
.A2(n_228),
.B1(n_208),
.B2(n_211),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_258),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_229),
.B1(n_206),
.B2(n_227),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_263),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_209),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_220),
.Y(n_271)
);

OA22x2_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_210),
.B1(n_224),
.B2(n_186),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_264),
.B(n_253),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_248),
.B(n_217),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_232),
.Y(n_270)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_262),
.Y(n_268)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_239),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_269),
.B(n_270),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_273),
.C(n_274),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_241),
.C(n_209),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_250),
.C(n_218),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_245),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_275),
.A2(n_252),
.B(n_222),
.Y(n_280)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_276),
.A2(n_263),
.B1(n_237),
.B2(n_238),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g282 ( 
.A(n_277),
.B(n_278),
.CI(n_253),
.CON(n_282),
.SN(n_282)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_222),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_276),
.A2(n_258),
.B(n_251),
.Y(n_279)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_279),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_280),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_272),
.A2(n_267),
.B(n_259),
.Y(n_281)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_285),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_277),
.A2(n_263),
.B1(n_256),
.B2(n_261),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_287),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_278),
.A2(n_233),
.B1(n_249),
.B2(n_240),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_252),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_271),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_266),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_295),
.B(n_283),
.Y(n_297)
);

NAND2xp33_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_233),
.Y(n_296)
);

AOI21x1_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_217),
.B(n_210),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_298),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_292),
.A2(n_281),
.B1(n_279),
.B2(n_285),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_299),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_273),
.B(n_284),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_301),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_304),
.A2(n_294),
.B(n_289),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_305),
.B(n_306),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_302),
.A2(n_294),
.B(n_284),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_293),
.B(n_303),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_290),
.Y(n_309)
);


endmodule