module fake_jpeg_30461_n_309 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_309);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_2),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_40),
.Y(n_54)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_29),
.B1(n_33),
.B2(n_31),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_45),
.A2(n_63),
.B1(n_34),
.B2(n_19),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_17),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_56),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_25),
.B(n_28),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_30),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_16),
.B1(n_23),
.B2(n_27),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_39),
.B1(n_24),
.B2(n_27),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_62),
.Y(n_102)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_21),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_33),
.B1(n_31),
.B2(n_16),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_70),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_61),
.A2(n_18),
.B1(n_28),
.B2(n_25),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_69),
.A2(n_72),
.B1(n_78),
.B2(n_79),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_18),
.B1(n_32),
.B2(n_28),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_73),
.A2(n_91),
.B1(n_106),
.B2(n_44),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_18),
.B1(n_16),
.B2(n_23),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_74),
.A2(n_99),
.B1(n_44),
.B2(n_42),
.Y(n_112)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_60),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_77),
.B(n_0),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_52),
.A2(n_25),
.B1(n_32),
.B2(n_26),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_52),
.A2(n_32),
.B1(n_26),
.B2(n_35),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_52),
.A2(n_26),
.B1(n_35),
.B2(n_23),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_80),
.A2(n_83),
.B1(n_86),
.B2(n_101),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_81),
.B(n_87),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_22),
.B(n_42),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_35),
.B1(n_16),
.B2(n_23),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_46),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_84),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_51),
.A2(n_35),
.B1(n_27),
.B2(n_24),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_54),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_90),
.Y(n_135)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_39),
.B1(n_27),
.B2(n_24),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_95),
.Y(n_124)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_96),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_46),
.A2(n_19),
.B(n_34),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_97),
.A2(n_91),
.B(n_84),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_65),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_41),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_46),
.A2(n_35),
.B1(n_19),
.B2(n_34),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_50),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_105),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_44),
.C(n_42),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_92),
.C(n_77),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_112),
.A2(n_113),
.B1(n_118),
.B2(n_132),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_81),
.A2(n_30),
.B1(n_44),
.B2(n_42),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_89),
.B1(n_76),
.B2(n_84),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_106),
.A2(n_35),
.B1(n_22),
.B2(n_12),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_117),
.B(n_113),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_102),
.A2(n_22),
.B1(n_41),
.B2(n_66),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_0),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_126),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_75),
.B(n_0),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_95),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_97),
.B(n_8),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_134),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_67),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_88),
.B(n_1),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_139),
.A2(n_148),
.B(n_152),
.Y(n_194)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_146),
.B1(n_166),
.B2(n_111),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_149),
.Y(n_174)
);

INVx2_ASAP7_75t_R g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_143),
.Y(n_197)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_114),
.A2(n_107),
.B1(n_93),
.B2(n_103),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_107),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_155),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_SL g152 ( 
.A(n_117),
.B(n_11),
.C(n_14),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_123),
.Y(n_177)
);

OAI32xp33_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_126),
.A3(n_130),
.B1(n_134),
.B2(n_115),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_168),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_93),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_119),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_160),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_92),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_118),
.B(n_103),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_161),
.B(n_164),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_96),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_167),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_120),
.A2(n_90),
.B(n_14),
.C(n_13),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_165),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_120),
.A2(n_98),
.B1(n_104),
.B2(n_105),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_116),
.B(n_94),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_111),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_159),
.A2(n_127),
.B1(n_112),
.B2(n_128),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_170),
.A2(n_182),
.B1(n_197),
.B2(n_180),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_136),
.C(n_137),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_177),
.C(n_179),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_172),
.A2(n_173),
.B1(n_147),
.B2(n_152),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_127),
.B1(n_132),
.B2(n_123),
.Y(n_173)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_185),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_136),
.C(n_122),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

BUFx24_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_181),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_123),
.B1(n_128),
.B2(n_101),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_139),
.A2(n_94),
.B(n_71),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_183),
.A2(n_160),
.B(n_161),
.Y(n_204)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_SL g199 ( 
.A1(n_184),
.A2(n_183),
.B(n_198),
.Y(n_199)
);

NAND3xp33_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_12),
.C(n_11),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_138),
.B(n_150),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_189),
.B(n_191),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_133),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_190),
.B(n_165),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_138),
.B(n_133),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_199),
.A2(n_202),
.B(n_209),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_178),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_158),
.Y(n_201)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_170),
.A2(n_166),
.B1(n_163),
.B2(n_164),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_189),
.B(n_145),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_205),
.B(n_217),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_151),
.C(n_145),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_208),
.C(n_220),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_151),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_196),
.A2(n_154),
.B(n_141),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_168),
.Y(n_210)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_146),
.Y(n_211)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_211),
.Y(n_232)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_187),
.B(n_157),
.Y(n_217)
);

AOI22x1_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_71),
.B1(n_108),
.B2(n_105),
.Y(n_218)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_219),
.A2(n_173),
.B1(n_172),
.B2(n_197),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_108),
.C(n_101),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_188),
.A2(n_108),
.B(n_85),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_175),
.B(n_169),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_85),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_223),
.B(n_181),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_1),
.Y(n_224)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_194),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_228),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_227),
.A2(n_230),
.B1(n_213),
.B2(n_216),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_201),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_231),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_192),
.B1(n_181),
.B2(n_178),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_184),
.Y(n_234)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_238),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_169),
.C(n_11),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_204),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_250),
.B1(n_262),
.B2(n_235),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_203),
.C(n_206),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_258),
.C(n_226),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_244),
.A2(n_209),
.B1(n_221),
.B2(n_215),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_212),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_232),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_224),
.Y(n_252)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_234),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_263),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_233),
.A2(n_215),
.B(n_220),
.Y(n_254)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_255),
.B(n_237),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_212),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_257),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_223),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_219),
.C(n_211),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_222),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_231),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_227),
.A2(n_226),
.B1(n_235),
.B2(n_242),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_1),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_267),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_274),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_269),
.A2(n_275),
.B1(n_218),
.B2(n_257),
.Y(n_278)
);

AO22x1_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_259),
.B1(n_261),
.B2(n_260),
.Y(n_270)
);

AOI21x1_ASAP7_75t_SL g287 ( 
.A1(n_270),
.A2(n_3),
.B(n_4),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_238),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_272),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_240),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_240),
.Y(n_273)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_273),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_247),
.A2(n_232),
.B1(n_236),
.B2(n_218),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_286),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_251),
.C(n_256),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_280),
.C(n_264),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_249),
.C(n_236),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g282 ( 
.A1(n_277),
.A2(n_2),
.B(n_3),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_282),
.A2(n_266),
.B(n_270),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_2),
.Y(n_286)
);

FAx1_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_3),
.CI(n_4),
.CON(n_294),
.SN(n_294)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_291),
.Y(n_300)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_283),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_268),
.C(n_265),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_293),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_285),
.Y(n_293)
);

AOI31xp33_ASAP7_75t_L g296 ( 
.A1(n_294),
.A2(n_295),
.A3(n_4),
.B(n_5),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_287),
.A2(n_273),
.B(n_264),
.Y(n_295)
);

AOI31xp67_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_6),
.A3(n_4),
.B(n_5),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_280),
.C(n_284),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_298),
.B(n_289),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_301),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_297),
.B(n_294),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_302),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_304),
.A2(n_299),
.B(n_300),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_305),
.C(n_298),
.Y(n_307)
);

OA21x2_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_303),
.B(n_5),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_6),
.Y(n_309)
);


endmodule