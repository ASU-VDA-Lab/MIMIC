module fake_jpeg_288_n_112 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_112);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_43),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_44),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_35),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_34),
.B(n_32),
.Y(n_50)
);

AO22x1_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_34),
.B1(n_32),
.B2(n_29),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_31),
.B1(n_30),
.B2(n_36),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_29),
.B1(n_33),
.B2(n_2),
.Y(n_60)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_59),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_62),
.Y(n_66)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_63),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_71),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_50),
.B(n_48),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_14),
.B(n_26),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_52),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_73),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_0),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_12),
.Y(n_73)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_77),
.B(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_74),
.B(n_73),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_63),
.B1(n_3),
.B2(n_4),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_1),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_81),
.B1(n_83),
.B2(n_75),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_13),
.B(n_24),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_92),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_11),
.C(n_23),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_20),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_94),
.B1(n_76),
.B2(n_8),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_27),
.B(n_22),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_96),
.B(n_100),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_101),
.C(n_87),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_89),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_88),
.B(n_9),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_97),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_93),
.B1(n_98),
.B2(n_103),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_102),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_108),
.B(n_90),
.Y(n_109)
);

NOR3xp33_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_94),
.C(n_10),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_110),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_21),
.Y(n_112)
);


endmodule