module real_aes_18285_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_1601, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_1601;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_571;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_1049;
wire n_559;
wire n_1277;
wire n_1584;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
OAI22xp33_ASAP7_75t_L g1197 ( .A1(n_0), .A2(n_90), .B1(n_690), .B2(n_693), .Y(n_1197) );
INVxp67_ASAP7_75t_SL g1211 ( .A(n_0), .Y(n_1211) );
CKINVDCx5p33_ASAP7_75t_R g855 ( .A(n_1), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g1330 ( .A1(n_2), .A2(n_7), .B1(n_1292), .B2(n_1295), .Y(n_1330) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_3), .Y(n_815) );
INVx1_ASAP7_75t_L g1248 ( .A(n_4), .Y(n_1248) );
AOI221xp5_ASAP7_75t_L g1265 ( .A1(n_4), .A2(n_148), .B1(n_714), .B2(n_1262), .C(n_1266), .Y(n_1265) );
CKINVDCx5p33_ASAP7_75t_R g1134 ( .A(n_5), .Y(n_1134) );
INVx1_ASAP7_75t_L g1183 ( .A(n_6), .Y(n_1183) );
INVx1_ASAP7_75t_L g336 ( .A(n_8), .Y(n_336) );
OAI221xp5_ASAP7_75t_SL g427 ( .A1(n_8), .A2(n_91), .B1(n_428), .B2(n_429), .C(n_433), .Y(n_427) );
INVx1_ASAP7_75t_L g502 ( .A(n_9), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_9), .A2(n_113), .B1(n_334), .B2(n_552), .Y(n_551) );
OAI221xp5_ASAP7_75t_L g491 ( .A1(n_10), .A2(n_226), .B1(n_428), .B2(n_429), .C(n_450), .Y(n_491) );
OA222x2_ASAP7_75t_L g567 ( .A1(n_10), .A2(n_50), .B1(n_229), .B2(n_568), .C1(n_572), .C2(n_576), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_11), .A2(n_73), .B1(n_562), .B2(n_611), .Y(n_924) );
OAI22xp33_ASAP7_75t_L g967 ( .A1(n_11), .A2(n_38), .B1(n_690), .B2(n_693), .Y(n_967) );
CKINVDCx5p33_ASAP7_75t_R g1077 ( .A(n_12), .Y(n_1077) );
INVx1_ASAP7_75t_L g297 ( .A(n_13), .Y(n_297) );
AND2x2_ASAP7_75t_L g338 ( .A(n_13), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g350 ( .A(n_13), .B(n_235), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_13), .B(n_307), .Y(n_530) );
INVx1_ASAP7_75t_L g1494 ( .A(n_14), .Y(n_1494) );
OAI221xp5_ASAP7_75t_SL g1522 ( .A1(n_14), .A2(n_272), .B1(n_1523), .B2(n_1526), .C(n_1529), .Y(n_1522) );
INVx1_ASAP7_75t_L g609 ( .A(n_15), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_15), .A2(n_263), .B1(n_627), .B2(n_630), .Y(n_626) );
INVx1_ASAP7_75t_L g1044 ( .A(n_16), .Y(n_1044) );
AOI22xp5_ASAP7_75t_L g1062 ( .A1(n_16), .A2(n_39), .B1(n_715), .B2(n_907), .Y(n_1062) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_17), .A2(n_122), .B1(n_673), .B2(n_675), .Y(n_672) );
INVxp67_ASAP7_75t_SL g723 ( .A(n_17), .Y(n_723) );
INVx2_ASAP7_75t_L g1288 ( .A(n_18), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_18), .B(n_108), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_18), .B(n_1294), .Y(n_1296) );
AOI21xp5_ASAP7_75t_L g1194 ( .A1(n_19), .A2(n_426), .B(n_1195), .Y(n_1194) );
INVx1_ASAP7_75t_L g1222 ( .A(n_19), .Y(n_1222) );
INVx1_ASAP7_75t_L g852 ( .A(n_20), .Y(n_852) );
OAI22xp5_ASAP7_75t_L g1235 ( .A1(n_21), .A2(n_240), .B1(n_673), .B2(n_675), .Y(n_1235) );
INVxp67_ASAP7_75t_SL g1269 ( .A(n_21), .Y(n_1269) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_22), .A2(n_154), .B1(n_521), .B2(n_638), .Y(n_1204) );
AOI32xp33_ASAP7_75t_L g1213 ( .A1(n_22), .A2(n_333), .A3(n_1214), .B1(n_1216), .B2(n_1601), .Y(n_1213) );
AOI22xp5_ASAP7_75t_L g1308 ( .A1(n_23), .A2(n_241), .B1(n_1292), .B2(n_1295), .Y(n_1308) );
CKINVDCx5p33_ASAP7_75t_R g1086 ( .A(n_24), .Y(n_1086) );
INVx1_ASAP7_75t_L g688 ( .A(n_25), .Y(n_688) );
OAI22xp33_ASAP7_75t_L g1111 ( .A1(n_26), .A2(n_267), .B1(n_299), .B2(n_1112), .Y(n_1111) );
OAI22xp33_ASAP7_75t_L g1143 ( .A1(n_26), .A2(n_267), .B1(n_1144), .B2(n_1147), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_27), .B(n_876), .Y(n_1196) );
AOI221xp5_ASAP7_75t_L g1225 ( .A1(n_27), .A2(n_154), .B1(n_329), .B2(n_839), .C(n_1067), .Y(n_1225) );
INVx1_ASAP7_75t_L g1004 ( .A(n_28), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1576 ( .A1(n_29), .A2(n_193), .B1(n_955), .B2(n_1505), .Y(n_1576) );
AOI22xp33_ASAP7_75t_L g1593 ( .A1(n_29), .A2(n_132), .B1(n_380), .B2(n_905), .Y(n_1593) );
AOI22xp33_ASAP7_75t_L g1575 ( .A1(n_30), .A2(n_132), .B1(n_955), .B2(n_1505), .Y(n_1575) );
AOI22xp33_ASAP7_75t_SL g1588 ( .A1(n_30), .A2(n_193), .B1(n_714), .B2(n_1514), .Y(n_1588) );
CKINVDCx5p33_ASAP7_75t_R g1091 ( .A(n_31), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_32), .A2(n_172), .B1(n_687), .B2(n_876), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_32), .A2(n_143), .B1(n_899), .B2(n_905), .Y(n_904) );
AOI222xp33_ASAP7_75t_L g700 ( .A1(n_33), .A2(n_181), .B1(n_223), .B2(n_479), .C1(n_512), .C2(n_648), .Y(n_700) );
INVx1_ASAP7_75t_L g734 ( .A(n_33), .Y(n_734) );
CKINVDCx5p33_ASAP7_75t_R g762 ( .A(n_34), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_35), .B(n_1193), .Y(n_1192) );
AOI22xp33_ASAP7_75t_L g1224 ( .A1(n_35), .A2(n_279), .B1(n_603), .B2(n_730), .Y(n_1224) );
AOI22xp5_ASAP7_75t_L g1300 ( .A1(n_36), .A2(n_271), .B1(n_1285), .B2(n_1301), .Y(n_1300) );
INVx1_ASAP7_75t_L g592 ( .A(n_37), .Y(n_592) );
OAI211xp5_ASAP7_75t_L g921 ( .A1(n_38), .A2(n_922), .B(n_923), .C(n_945), .Y(n_921) );
INVx1_ASAP7_75t_L g1052 ( .A(n_39), .Y(n_1052) );
INVx1_ASAP7_75t_L g1049 ( .A(n_40), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_40), .A2(n_179), .B1(n_603), .B2(n_715), .Y(n_1065) );
INVx1_ASAP7_75t_L g860 ( .A(n_41), .Y(n_860) );
INVx1_ASAP7_75t_L g1069 ( .A(n_42), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g1499 ( .A1(n_43), .A2(n_78), .B1(n_878), .B2(n_1500), .Y(n_1499) );
INVxp67_ASAP7_75t_SL g1531 ( .A(n_43), .Y(n_1531) );
AOI22xp5_ASAP7_75t_L g1320 ( .A1(n_44), .A2(n_250), .B1(n_1292), .B2(n_1295), .Y(n_1320) );
OAI21xp33_ASAP7_75t_L g594 ( .A1(n_45), .A2(n_568), .B(n_595), .Y(n_594) );
OAI221xp5_ASAP7_75t_L g650 ( .A1(n_45), .A2(n_53), .B1(n_651), .B2(n_652), .C(n_654), .Y(n_650) );
AO22x1_ASAP7_75t_L g1305 ( .A1(n_46), .A2(n_62), .B1(n_1285), .B2(n_1289), .Y(n_1305) );
OAI22xp33_ASAP7_75t_L g825 ( .A1(n_47), .A2(n_170), .B1(n_630), .B2(n_671), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_47), .A2(n_82), .B1(n_560), .B2(n_565), .Y(n_844) );
AOI221xp5_ASAP7_75t_L g1237 ( .A1(n_48), .A2(n_118), .B1(n_883), .B2(n_1238), .C(n_1240), .Y(n_1237) );
INVx1_ASAP7_75t_L g1264 ( .A(n_48), .Y(n_1264) );
INVx1_ASAP7_75t_L g396 ( .A(n_49), .Y(n_396) );
INVx1_ASAP7_75t_L g417 ( .A(n_49), .Y(n_417) );
INVx1_ASAP7_75t_L g489 ( .A(n_50), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_51), .A2(n_156), .B1(n_344), .B2(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g448 ( .A(n_51), .Y(n_448) );
INVx1_ASAP7_75t_L g612 ( .A(n_52), .Y(n_612) );
INVxp67_ASAP7_75t_SL g662 ( .A(n_53), .Y(n_662) );
CKINVDCx5p33_ASAP7_75t_R g752 ( .A(n_54), .Y(n_752) );
CKINVDCx5p33_ASAP7_75t_R g767 ( .A(n_55), .Y(n_767) );
INVx1_ASAP7_75t_L g995 ( .A(n_56), .Y(n_995) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_57), .A2(n_163), .B1(n_679), .B2(n_681), .C(n_683), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_57), .A2(n_228), .B1(n_728), .B2(n_730), .C(n_732), .Y(n_727) );
OAI221xp5_ASAP7_75t_L g1033 ( .A1(n_58), .A2(n_110), .B1(n_673), .B2(n_675), .C(n_1034), .Y(n_1033) );
INVxp67_ASAP7_75t_SL g1057 ( .A(n_58), .Y(n_1057) );
OAI221xp5_ASAP7_75t_L g670 ( .A1(n_59), .A2(n_254), .B1(n_630), .B2(n_634), .C(n_671), .Y(n_670) );
OAI21xp33_ASAP7_75t_SL g711 ( .A1(n_59), .A2(n_554), .B(n_576), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_60), .A2(n_248), .B1(n_673), .B2(n_675), .Y(n_952) );
INVxp67_ASAP7_75t_SL g972 ( .A(n_60), .Y(n_972) );
INVx1_ASAP7_75t_L g290 ( .A(n_61), .Y(n_290) );
INVx2_ASAP7_75t_L g403 ( .A(n_63), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g1087 ( .A(n_64), .Y(n_1087) );
INVx1_ASAP7_75t_L g812 ( .A(n_65), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_65), .A2(n_231), .B1(n_344), .B2(n_373), .Y(n_838) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_66), .Y(n_824) );
OAI22xp33_ASAP7_75t_L g689 ( .A1(n_67), .A2(n_72), .B1(n_690), .B2(n_693), .Y(n_689) );
INVxp67_ASAP7_75t_SL g706 ( .A(n_67), .Y(n_706) );
AOI21xp33_ASAP7_75t_L g999 ( .A1(n_68), .A2(n_454), .B(n_642), .Y(n_999) );
INVxp67_ASAP7_75t_L g1017 ( .A(n_68), .Y(n_1017) );
INVx1_ASAP7_75t_L g773 ( .A(n_69), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g1321 ( .A1(n_70), .A2(n_182), .B1(n_1285), .B2(n_1289), .Y(n_1321) );
INVx1_ASAP7_75t_L g1175 ( .A(n_71), .Y(n_1175) );
AO221x2_ASAP7_75t_L g1362 ( .A1(n_71), .A2(n_225), .B1(n_1292), .B2(n_1295), .C(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g710 ( .A(n_72), .Y(n_710) );
OAI221xp5_ASAP7_75t_L g951 ( .A1(n_73), .A2(n_125), .B1(n_630), .B2(n_634), .C(n_671), .Y(n_951) );
INVx1_ASAP7_75t_L g1249 ( .A(n_74), .Y(n_1249) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_75), .A2(n_183), .B1(n_363), .B2(n_369), .C(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g449 ( .A(n_75), .Y(n_449) );
INVx1_ASAP7_75t_L g669 ( .A(n_76), .Y(n_669) );
OAI21xp33_ASAP7_75t_L g707 ( .A1(n_76), .A2(n_572), .B(n_708), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g1501 ( .A1(n_77), .A2(n_252), .B1(n_648), .B2(n_1502), .Y(n_1501) );
AOI22xp33_ASAP7_75t_L g1516 ( .A1(n_77), .A2(n_221), .B1(n_329), .B2(n_1067), .Y(n_1516) );
AOI221xp5_ASAP7_75t_L g1513 ( .A1(n_78), .A2(n_102), .B1(n_896), .B2(n_908), .C(n_1514), .Y(n_1513) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_79), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_80), .A2(n_260), .B1(n_1116), .B2(n_1119), .Y(n_1115) );
OAI22xp33_ASAP7_75t_L g1164 ( .A1(n_80), .A2(n_260), .B1(n_1165), .B2(n_1167), .Y(n_1164) );
INVx1_ASAP7_75t_L g506 ( .A(n_81), .Y(n_506) );
AOI221x1_ASAP7_75t_SL g531 ( .A1(n_81), .A2(n_99), .B1(n_363), .B2(n_373), .C(n_532), .Y(n_531) );
OAI221xp5_ASAP7_75t_L g820 ( .A1(n_82), .A2(n_169), .B1(n_821), .B2(n_822), .C(n_823), .Y(n_820) );
OAI222xp33_ASAP7_75t_L g779 ( .A1(n_83), .A2(n_133), .B1(n_246), .B2(n_408), .C1(n_505), .C2(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g797 ( .A(n_83), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g1503 ( .A1(n_84), .A2(n_221), .B1(n_1504), .B2(n_1505), .Y(n_1503) );
AOI221xp5_ASAP7_75t_L g1533 ( .A1(n_84), .A2(n_252), .B1(n_333), .B2(n_714), .C(n_1534), .Y(n_1533) );
INVx1_ASAP7_75t_L g1050 ( .A(n_85), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_85), .A2(n_237), .B1(n_344), .B2(n_373), .Y(n_1063) );
AOI22xp33_ASAP7_75t_SL g866 ( .A1(n_86), .A2(n_96), .B1(n_867), .B2(n_869), .Y(n_866) );
AOI221xp5_ASAP7_75t_L g895 ( .A1(n_86), .A2(n_131), .B1(n_333), .B2(n_730), .C(n_896), .Y(n_895) );
XOR2x1_ASAP7_75t_L g1178 ( .A(n_87), .B(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g940 ( .A(n_88), .Y(n_940) );
AOI221xp5_ASAP7_75t_L g1245 ( .A1(n_89), .A2(n_100), .B1(n_520), .B2(n_1246), .C(n_1247), .Y(n_1245) );
INVx1_ASAP7_75t_L g1268 ( .A(n_89), .Y(n_1268) );
INVx1_ASAP7_75t_L g1180 ( .A(n_90), .Y(n_1180) );
INVx1_ASAP7_75t_L g355 ( .A(n_91), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g1040 ( .A(n_92), .Y(n_1040) );
INVx1_ASAP7_75t_L g484 ( .A(n_93), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_93), .A2(n_226), .B1(n_560), .B2(n_565), .Y(n_559) );
INVx1_ASAP7_75t_L g1553 ( .A(n_94), .Y(n_1553) );
OAI22xp5_ASAP7_75t_L g1005 ( .A1(n_95), .A2(n_186), .B1(n_690), .B2(n_693), .Y(n_1005) );
INVxp67_ASAP7_75t_SL g1007 ( .A(n_95), .Y(n_1007) );
AOI221xp5_ASAP7_75t_L g906 ( .A1(n_96), .A2(n_211), .B1(n_907), .B2(n_908), .C(n_912), .Y(n_906) );
INVx1_ASAP7_75t_L g766 ( .A(n_97), .Y(n_766) );
AOI221xp5_ASAP7_75t_L g784 ( .A1(n_97), .A2(n_153), .B1(n_478), .B2(n_785), .C(n_788), .Y(n_784) );
OAI221xp5_ASAP7_75t_L g320 ( .A1(n_98), .A2(n_280), .B1(n_321), .B2(n_323), .C(n_328), .Y(n_320) );
INVx1_ASAP7_75t_L g387 ( .A(n_98), .Y(n_387) );
INVx1_ASAP7_75t_L g522 ( .A(n_99), .Y(n_522) );
AOI221xp5_ASAP7_75t_L g1261 ( .A1(n_100), .A2(n_195), .B1(n_714), .B2(n_1262), .C(n_1263), .Y(n_1261) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_101), .Y(n_292) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_101), .B(n_290), .Y(n_1286) );
AOI22xp33_ASAP7_75t_SL g1506 ( .A1(n_102), .A2(n_166), .B1(n_389), .B2(n_1507), .Y(n_1506) );
INVx1_ASAP7_75t_L g1556 ( .A(n_103), .Y(n_1556) );
OAI22xp5_ASAP7_75t_L g1563 ( .A1(n_103), .A2(n_264), .B1(n_1564), .B2(n_1566), .Y(n_1563) );
OAI21xp5_ASAP7_75t_SL g915 ( .A1(n_104), .A2(n_916), .B(n_917), .Y(n_915) );
INVx1_ASAP7_75t_L g974 ( .A(n_105), .Y(n_974) );
XNOR2xp5_ASAP7_75t_L g1487 ( .A(n_106), .B(n_1488), .Y(n_1487) );
AOI22xp33_ASAP7_75t_SL g602 ( .A1(n_107), .A2(n_188), .B1(n_365), .B2(n_603), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g639 ( .A1(n_107), .A2(n_173), .B1(n_640), .B2(n_641), .C(n_642), .Y(n_639) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_108), .B(n_1288), .Y(n_1287) );
INVx1_ASAP7_75t_L g1294 ( .A(n_108), .Y(n_1294) );
INVx1_ASAP7_75t_L g1497 ( .A(n_109), .Y(n_1497) );
INVx1_ASAP7_75t_L g1068 ( .A(n_110), .Y(n_1068) );
AOI221xp5_ASAP7_75t_L g1198 ( .A1(n_111), .A2(n_279), .B1(n_1199), .B2(n_1202), .C(n_1203), .Y(n_1198) );
INVx1_ASAP7_75t_L g1223 ( .A(n_111), .Y(n_1223) );
INVx1_ASAP7_75t_L g1558 ( .A(n_112), .Y(n_1558) );
INVx1_ASAP7_75t_L g513 ( .A(n_113), .Y(n_513) );
XNOR2xp5_ASAP7_75t_L g846 ( .A(n_114), .B(n_847), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g1185 ( .A1(n_115), .A2(n_269), .B1(n_673), .B2(n_675), .Y(n_1185) );
INVxp33_ASAP7_75t_L g1227 ( .A(n_115), .Y(n_1227) );
INVx1_ASAP7_75t_L g347 ( .A(n_116), .Y(n_347) );
OAI21xp33_ASAP7_75t_L g420 ( .A1(n_116), .A2(n_421), .B(n_425), .Y(n_420) );
OAI22xp33_ASAP7_75t_L g1244 ( .A1(n_117), .A2(n_161), .B1(n_690), .B2(n_693), .Y(n_1244) );
INVxp67_ASAP7_75t_SL g1271 ( .A(n_117), .Y(n_1271) );
INVx1_ASAP7_75t_L g1267 ( .A(n_118), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_119), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g440 ( .A(n_119), .Y(n_440) );
INVx1_ASAP7_75t_L g468 ( .A(n_119), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g807 ( .A(n_120), .Y(n_807) );
INVx1_ASAP7_75t_L g774 ( .A(n_121), .Y(n_774) );
OAI22xp33_ASAP7_75t_L g782 ( .A1(n_121), .A2(n_160), .B1(n_630), .B2(n_671), .Y(n_782) );
INVxp67_ASAP7_75t_SL g703 ( .A(n_122), .Y(n_703) );
INVx1_ASAP7_75t_L g997 ( .A(n_123), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g1329 ( .A1(n_124), .A2(n_219), .B1(n_1285), .B2(n_1289), .Y(n_1329) );
INVxp67_ASAP7_75t_SL g947 ( .A(n_125), .Y(n_947) );
INVx1_ASAP7_75t_L g1550 ( .A(n_126), .Y(n_1550) );
AOI22xp33_ASAP7_75t_SL g1572 ( .A1(n_127), .A2(n_147), .B1(n_1573), .B2(n_1574), .Y(n_1572) );
AOI22xp33_ASAP7_75t_SL g1589 ( .A1(n_127), .A2(n_222), .B1(n_714), .B2(n_1590), .Y(n_1589) );
OAI221xp5_ASAP7_75t_L g1184 ( .A1(n_128), .A2(n_157), .B1(n_630), .B2(n_634), .C(n_671), .Y(n_1184) );
NOR2xp33_ASAP7_75t_L g1215 ( .A(n_128), .B(n_599), .Y(n_1215) );
XOR2xp5_ASAP7_75t_L g469 ( .A(n_129), .B(n_470), .Y(n_469) );
AOI221xp5_ASAP7_75t_L g941 ( .A1(n_130), .A2(n_149), .B1(n_935), .B2(n_942), .C(n_944), .Y(n_941) );
AOI221xp5_ASAP7_75t_L g963 ( .A1(n_130), .A2(n_159), .B1(n_426), .B2(n_956), .C(n_964), .Y(n_963) );
AOI221xp5_ASAP7_75t_L g877 ( .A1(n_131), .A2(n_143), .B1(n_869), .B2(n_878), .C(n_879), .Y(n_877) );
OAI221xp5_ASAP7_75t_L g770 ( .A1(n_133), .A2(n_160), .B1(n_554), .B2(n_560), .C(n_565), .Y(n_770) );
INVx1_ASAP7_75t_L g741 ( .A(n_134), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_135), .A2(n_315), .B1(n_316), .B2(n_317), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_135), .Y(n_315) );
AOI22xp33_ASAP7_75t_SL g604 ( .A1(n_136), .A2(n_265), .B1(n_379), .B2(n_605), .Y(n_604) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_136), .A2(n_217), .B1(n_426), .B2(n_640), .C(n_644), .Y(n_643) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_137), .Y(n_509) );
INVx1_ASAP7_75t_L g938 ( .A(n_138), .Y(n_938) );
AOI221xp5_ASAP7_75t_L g954 ( .A1(n_138), .A2(n_281), .B1(n_955), .B2(n_956), .C(n_957), .Y(n_954) );
INVx1_ASAP7_75t_L g1053 ( .A(n_139), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_139), .A2(n_190), .B1(n_329), .B2(n_1067), .Y(n_1066) );
OAI221xp5_ASAP7_75t_L g1234 ( .A1(n_140), .A2(n_196), .B1(n_630), .B2(n_634), .C(n_671), .Y(n_1234) );
OAI21xp33_ASAP7_75t_L g1257 ( .A1(n_140), .A2(n_554), .B(n_576), .Y(n_1257) );
OAI22xp33_ASAP7_75t_L g485 ( .A1(n_141), .A2(n_146), .B1(n_486), .B2(n_487), .Y(n_485) );
INVx1_ASAP7_75t_L g585 ( .A(n_141), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_142), .A2(n_191), .B1(n_379), .B2(n_380), .Y(n_378) );
INVx1_ASAP7_75t_L g462 ( .A(n_142), .Y(n_462) );
XOR2x2_ASAP7_75t_L g981 ( .A(n_144), .B(n_982), .Y(n_981) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_145), .A2(n_675), .B1(n_810), .B2(n_813), .Y(n_809) );
INVx1_ASAP7_75t_L g831 ( .A(n_145), .Y(n_831) );
INVx1_ASAP7_75t_L g581 ( .A(n_146), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g1585 ( .A1(n_147), .A2(n_275), .B1(n_905), .B2(n_1586), .Y(n_1585) );
INVx1_ASAP7_75t_L g1241 ( .A(n_148), .Y(n_1241) );
INVx1_ASAP7_75t_L g960 ( .A(n_149), .Y(n_960) );
AO22x1_ASAP7_75t_L g1306 ( .A1(n_150), .A2(n_239), .B1(n_1292), .B2(n_1295), .Y(n_1306) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_151), .A2(n_216), .B1(n_379), .B2(n_615), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_151), .A2(n_265), .B1(n_426), .B2(n_638), .Y(n_637) );
AOI221xp5_ASAP7_75t_SL g362 ( .A1(n_152), .A2(n_174), .B1(n_363), .B2(n_369), .C(n_370), .Y(n_362) );
INVx1_ASAP7_75t_L g452 ( .A(n_152), .Y(n_452) );
INVx1_ASAP7_75t_L g748 ( .A(n_153), .Y(n_748) );
BUFx3_ASAP7_75t_L g393 ( .A(n_155), .Y(n_393) );
INVx1_ASAP7_75t_L g464 ( .A(n_156), .Y(n_464) );
INVxp67_ASAP7_75t_SL g1210 ( .A(n_157), .Y(n_1210) );
INVx1_ASAP7_75t_L g1233 ( .A(n_158), .Y(n_1233) );
AOI221xp5_ASAP7_75t_L g932 ( .A1(n_159), .A2(n_209), .B1(n_839), .B2(n_933), .C(n_935), .Y(n_932) );
OAI22xp5_ASAP7_75t_L g1258 ( .A1(n_161), .A2(n_196), .B1(n_565), .B2(n_1259), .Y(n_1258) );
INVx1_ASAP7_75t_L g985 ( .A(n_162), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_163), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g685 ( .A(n_164), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g1291 ( .A1(n_165), .A2(n_177), .B1(n_1292), .B2(n_1295), .Y(n_1291) );
INVxp67_ASAP7_75t_SL g1532 ( .A(n_166), .Y(n_1532) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_167), .Y(n_304) );
INVx1_ASAP7_75t_L g596 ( .A(n_168), .Y(n_596) );
OAI211xp5_ASAP7_75t_L g829 ( .A1(n_169), .A2(n_661), .B(n_830), .C(n_833), .Y(n_829) );
INVx1_ASAP7_75t_L g832 ( .A(n_170), .Y(n_832) );
CKINVDCx5p33_ASAP7_75t_R g806 ( .A(n_171), .Y(n_806) );
AOI22xp33_ASAP7_75t_SL g897 ( .A1(n_172), .A2(n_270), .B1(n_898), .B2(n_899), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_173), .A2(n_217), .B1(n_618), .B2(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g461 ( .A(n_174), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g990 ( .A1(n_175), .A2(n_426), .B(n_644), .Y(n_990) );
INVxp67_ASAP7_75t_SL g1014 ( .A(n_175), .Y(n_1014) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_176), .Y(n_360) );
OAI222xp33_ASAP7_75t_L g1508 ( .A1(n_178), .A2(n_220), .B1(n_244), .B2(n_850), .C1(n_854), .C2(n_916), .Y(n_1508) );
OAI211xp5_ASAP7_75t_L g1510 ( .A1(n_178), .A2(n_1511), .B(n_1512), .C(n_1517), .Y(n_1510) );
INVx1_ASAP7_75t_L g1043 ( .A(n_179), .Y(n_1043) );
INVx1_ASAP7_75t_L g1138 ( .A(n_180), .Y(n_1138) );
OAI211xp5_ASAP7_75t_L g1150 ( .A1(n_180), .A2(n_1151), .B(n_1153), .C(n_1155), .Y(n_1150) );
INVx1_ASAP7_75t_L g719 ( .A(n_181), .Y(n_719) );
INVx1_ASAP7_75t_L g465 ( .A(n_183), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g761 ( .A(n_184), .Y(n_761) );
INVx1_ASAP7_75t_L g817 ( .A(n_185), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_185), .A2(n_194), .B1(n_344), .B2(n_381), .Y(n_843) );
OAI221xp5_ASAP7_75t_L g1025 ( .A1(n_186), .A2(n_212), .B1(n_554), .B2(n_560), .C(n_565), .Y(n_1025) );
AOI22xp5_ASAP7_75t_L g1309 ( .A1(n_187), .A2(n_249), .B1(n_1285), .B2(n_1289), .Y(n_1309) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_188), .A2(n_216), .B1(n_638), .B2(n_646), .Y(n_645) );
CKINVDCx5p33_ASAP7_75t_R g1078 ( .A(n_189), .Y(n_1078) );
INVx1_ASAP7_75t_L g1047 ( .A(n_190), .Y(n_1047) );
INVx1_ASAP7_75t_L g458 ( .A(n_191), .Y(n_458) );
INVx1_ASAP7_75t_L g1003 ( .A(n_192), .Y(n_1003) );
AOI221xp5_ASAP7_75t_L g804 ( .A1(n_194), .A2(n_231), .B1(n_638), .B2(n_787), .C(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g1243 ( .A(n_195), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1284 ( .A1(n_197), .A2(n_245), .B1(n_1285), .B2(n_1289), .Y(n_1284) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_198), .Y(n_303) );
INVx1_ASAP7_75t_L g992 ( .A(n_199), .Y(n_992) );
INVx1_ASAP7_75t_L g1036 ( .A(n_200), .Y(n_1036) );
OAI22xp5_ASAP7_75t_L g1060 ( .A1(n_200), .A2(n_202), .B1(n_562), .B2(n_611), .Y(n_1060) );
OAI211xp5_ASAP7_75t_L g1125 ( .A1(n_201), .A2(n_1126), .B(n_1129), .C(n_1132), .Y(n_1125) );
INVx1_ASAP7_75t_L g1163 ( .A(n_201), .Y(n_1163) );
INVx1_ASAP7_75t_L g1039 ( .A(n_202), .Y(n_1039) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_203), .Y(n_499) );
XNOR2x1_ASAP7_75t_L g1229 ( .A(n_204), .B(n_1230), .Y(n_1229) );
CKINVDCx5p33_ASAP7_75t_R g811 ( .A(n_205), .Y(n_811) );
CKINVDCx5p33_ASAP7_75t_R g1093 ( .A(n_206), .Y(n_1093) );
CKINVDCx5p33_ASAP7_75t_R g756 ( .A(n_207), .Y(n_756) );
INVxp67_ASAP7_75t_SL g772 ( .A(n_208), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_208), .A2(n_675), .B1(n_790), .B2(n_791), .Y(n_789) );
INVx1_ASAP7_75t_L g958 ( .A(n_209), .Y(n_958) );
INVx1_ASAP7_75t_L g946 ( .A(n_210), .Y(n_946) );
AOI22xp33_ASAP7_75t_SL g882 ( .A1(n_211), .A2(n_270), .B1(n_867), .B2(n_883), .Y(n_882) );
OAI221xp5_ASAP7_75t_L g986 ( .A1(n_212), .A2(n_243), .B1(n_630), .B2(n_634), .C(n_671), .Y(n_986) );
CKINVDCx5p33_ASAP7_75t_R g1084 ( .A(n_213), .Y(n_1084) );
INVx1_ASAP7_75t_L g1189 ( .A(n_214), .Y(n_1189) );
AO22x1_ASAP7_75t_L g1339 ( .A1(n_215), .A2(n_242), .B1(n_1285), .B2(n_1340), .Y(n_1339) );
AOI22xp33_ASAP7_75t_L g1538 ( .A1(n_215), .A2(n_1539), .B1(n_1541), .B2(n_1594), .Y(n_1538) );
XNOR2xp5_ASAP7_75t_L g1543 ( .A(n_215), .B(n_1544), .Y(n_1543) );
CKINVDCx16_ASAP7_75t_R g1364 ( .A(n_218), .Y(n_1364) );
AOI22xp33_ASAP7_75t_SL g1578 ( .A1(n_222), .A2(n_275), .B1(n_426), .B2(n_1579), .Y(n_1578) );
AOI21xp33_ASAP7_75t_L g721 ( .A1(n_223), .A2(n_333), .B(n_722), .Y(n_721) );
OAI211xp5_ASAP7_75t_L g1037 ( .A1(n_224), .A2(n_634), .B(n_659), .C(n_1038), .Y(n_1037) );
INVxp33_ASAP7_75t_SL g1059 ( .A(n_224), .Y(n_1059) );
INVx1_ASAP7_75t_L g887 ( .A(n_227), .Y(n_887) );
AOI21xp33_ASAP7_75t_L g695 ( .A1(n_228), .A2(n_696), .B(n_699), .Y(n_695) );
INVx1_ASAP7_75t_L g480 ( .A(n_229), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g749 ( .A(n_230), .Y(n_749) );
INVx1_ASAP7_75t_L g858 ( .A(n_232), .Y(n_858) );
AOI22xp5_ASAP7_75t_L g1299 ( .A1(n_233), .A2(n_258), .B1(n_1292), .B2(n_1295), .Y(n_1299) );
INVx1_ASAP7_75t_L g1548 ( .A(n_234), .Y(n_1548) );
BUFx3_ASAP7_75t_L g307 ( .A(n_235), .Y(n_307) );
INVx1_ASAP7_75t_L g339 ( .A(n_235), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g1082 ( .A(n_236), .Y(n_1082) );
INVx1_ASAP7_75t_L g1046 ( .A(n_237), .Y(n_1046) );
CKINVDCx20_ASAP7_75t_R g1366 ( .A(n_238), .Y(n_1366) );
INVxp67_ASAP7_75t_SL g1252 ( .A(n_240), .Y(n_1252) );
INVxp67_ASAP7_75t_SL g1027 ( .A(n_243), .Y(n_1027) );
INVx1_ASAP7_75t_L g776 ( .A(n_246), .Y(n_776) );
INVx2_ASAP7_75t_L g384 ( .A(n_247), .Y(n_384) );
INVx1_ASAP7_75t_L g401 ( .A(n_247), .Y(n_401) );
INVx1_ASAP7_75t_L g436 ( .A(n_247), .Y(n_436) );
INVxp67_ASAP7_75t_SL g948 ( .A(n_248), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_251), .A2(n_262), .B1(n_479), .B2(n_787), .Y(n_1000) );
INVxp67_ASAP7_75t_SL g1023 ( .A(n_251), .Y(n_1023) );
INVx1_ASAP7_75t_L g890 ( .A(n_253), .Y(n_890) );
INVx1_ASAP7_75t_L g709 ( .A(n_254), .Y(n_709) );
AO22x1_ASAP7_75t_L g1341 ( .A1(n_255), .A2(n_273), .B1(n_1292), .B2(n_1295), .Y(n_1341) );
INVx1_ASAP7_75t_L g800 ( .A(n_256), .Y(n_800) );
INVx1_ASAP7_75t_L g1496 ( .A(n_257), .Y(n_1496) );
XOR2x2_ASAP7_75t_L g665 ( .A(n_258), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g819 ( .A(n_259), .Y(n_819) );
INVx1_ASAP7_75t_L g989 ( .A(n_261), .Y(n_989) );
INVxp67_ASAP7_75t_SL g1013 ( .A(n_262), .Y(n_1013) );
INVx1_ASAP7_75t_L g597 ( .A(n_263), .Y(n_597) );
INVx1_ASAP7_75t_L g1555 ( .A(n_264), .Y(n_1555) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_266), .Y(n_517) );
OAI21xp33_ASAP7_75t_SL g1031 ( .A1(n_268), .A2(n_922), .B(n_1032), .Y(n_1031) );
INVx1_ASAP7_75t_L g1035 ( .A(n_268), .Y(n_1035) );
INVxp67_ASAP7_75t_SL g1206 ( .A(n_269), .Y(n_1206) );
INVx1_ASAP7_75t_L g1493 ( .A(n_272), .Y(n_1493) );
INVx1_ASAP7_75t_L g1552 ( .A(n_274), .Y(n_1552) );
INVxp67_ASAP7_75t_SL g588 ( .A(n_276), .Y(n_588) );
NAND2xp33_ASAP7_75t_SL g930 ( .A(n_277), .B(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g965 ( .A(n_277), .Y(n_965) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_278), .Y(n_332) );
INVx1_ASAP7_75t_L g405 ( .A(n_280), .Y(n_405) );
INVx1_ASAP7_75t_L g927 ( .A(n_281), .Y(n_927) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_308), .B(n_1276), .Y(n_282) );
INVx2_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_293), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g1540 ( .A(n_287), .B(n_296), .Y(n_1540) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g1537 ( .A(n_289), .B(n_292), .Y(n_1537) );
INVx1_ASAP7_75t_L g1597 ( .A(n_289), .Y(n_1597) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g1599 ( .A(n_292), .B(n_1597), .Y(n_1599) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_298), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g1140 ( .A(n_296), .B(n_1141), .Y(n_1140) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_L g371 ( .A(n_297), .B(n_306), .Y(n_371) );
AND2x4_ASAP7_75t_L g377 ( .A(n_297), .B(n_307), .Y(n_377) );
AND2x4_ASAP7_75t_SL g1539 ( .A(n_298), .B(n_1540), .Y(n_1539) );
AOI22xp33_ASAP7_75t_L g1551 ( .A1(n_298), .A2(n_1113), .B1(n_1552), .B2(n_1553), .Y(n_1551) );
INVx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x6_ASAP7_75t_L g299 ( .A(n_300), .B(n_305), .Y(n_299) );
BUFx4f_ASAP7_75t_L g718 ( .A(n_300), .Y(n_718) );
INVxp67_ASAP7_75t_L g765 ( .A(n_300), .Y(n_765) );
OR2x6_ASAP7_75t_L g1118 ( .A(n_300), .B(n_1114), .Y(n_1118) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx4f_ASAP7_75t_L g322 ( .A(n_301), .Y(n_322) );
INVx3_ASAP7_75t_L g534 ( .A(n_301), .Y(n_534) );
INVx3_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx2_ASAP7_75t_L g327 ( .A(n_303), .Y(n_327) );
INVx2_ASAP7_75t_L g331 ( .A(n_303), .Y(n_331) );
AND2x2_ASAP7_75t_L g335 ( .A(n_303), .B(n_304), .Y(n_335) );
INVx1_ASAP7_75t_L g359 ( .A(n_303), .Y(n_359) );
AND2x2_ASAP7_75t_L g367 ( .A(n_303), .B(n_368), .Y(n_367) );
NAND2x1_ASAP7_75t_L g537 ( .A(n_303), .B(n_304), .Y(n_537) );
OR2x2_ASAP7_75t_L g326 ( .A(n_304), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g330 ( .A(n_304), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g346 ( .A(n_304), .Y(n_346) );
BUFx2_ASAP7_75t_L g354 ( .A(n_304), .Y(n_354) );
INVx2_ASAP7_75t_L g368 ( .A(n_304), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_304), .B(n_331), .Y(n_550) );
INVxp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g1131 ( .A(n_306), .Y(n_1131) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx2_ASAP7_75t_L g1124 ( .A(n_307), .Y(n_1124) );
AND2x4_ASAP7_75t_L g1137 ( .A(n_307), .B(n_358), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_977), .B1(n_1274), .B2(n_1275), .Y(n_308) );
INVx1_ASAP7_75t_L g1274 ( .A(n_309), .Y(n_1274) );
BUFx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
XOR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_737), .Y(n_310) );
XNOR2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_586), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
XNOR2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_469), .Y(n_313) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_385), .Y(n_317) );
AOI21xp5_ASAP7_75t_SL g318 ( .A1(n_319), .A2(n_361), .B(n_382), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_337), .B(n_340), .Y(n_319) );
INVx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx6f_ASAP7_75t_L g1098 ( .A(n_322), .Y(n_1098) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx4_ASAP7_75t_L g755 ( .A(n_324), .Y(n_755) );
INVx4_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g545 ( .A(n_326), .Y(n_545) );
INVx2_ASAP7_75t_L g760 ( .A(n_326), .Y(n_760) );
BUFx3_ASAP7_75t_L g836 ( .A(n_326), .Y(n_836) );
BUFx2_ASAP7_75t_L g1019 ( .A(n_326), .Y(n_1019) );
AND2x2_ASAP7_75t_L g345 ( .A(n_327), .B(n_346), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_332), .B1(n_333), .B2(n_336), .Y(n_328) );
BUFx3_ASAP7_75t_L g899 ( .A(n_329), .Y(n_899) );
INVx1_ASAP7_75t_SL g1587 ( .A(n_329), .Y(n_1587) );
BUFx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g374 ( .A(n_330), .Y(n_374) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_330), .Y(n_381) );
BUFx3_ASAP7_75t_L g605 ( .A(n_330), .Y(n_605) );
A2O1A1Ixp33_ASAP7_75t_L g425 ( .A1(n_332), .A2(n_426), .B(n_427), .C(n_434), .Y(n_425) );
A2O1A1Ixp33_ASAP7_75t_L g341 ( .A1(n_333), .A2(n_342), .B(n_347), .C(n_348), .Y(n_341) );
BUFx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx3_ASAP7_75t_L g369 ( .A(n_334), .Y(n_369) );
BUFx3_ASAP7_75t_L g603 ( .A(n_334), .Y(n_603) );
BUFx6f_ASAP7_75t_L g729 ( .A(n_334), .Y(n_729) );
AND2x6_ASAP7_75t_L g900 ( .A(n_334), .B(n_350), .Y(n_900) );
AND2x4_ASAP7_75t_SL g903 ( .A(n_334), .B(n_338), .Y(n_903) );
BUFx3_ASAP7_75t_L g907 ( .A(n_334), .Y(n_907) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_334), .B(n_1131), .Y(n_1130) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g621 ( .A(n_335), .Y(n_621) );
BUFx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_338), .B(n_436), .Y(n_575) );
AND2x2_ASAP7_75t_L g580 ( .A(n_338), .B(n_345), .Y(n_580) );
AND2x2_ASAP7_75t_L g583 ( .A(n_338), .B(n_584), .Y(n_583) );
AND2x4_ASAP7_75t_L g892 ( .A(n_338), .B(n_584), .Y(n_892) );
AND2x4_ASAP7_75t_L g894 ( .A(n_338), .B(n_381), .Y(n_894) );
HB1xp67_ASAP7_75t_L g1114 ( .A(n_339), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_351), .Y(n_340) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_344), .Y(n_379) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_344), .B(n_1124), .Y(n_1549) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx3_ASAP7_75t_L g553 ( .A(n_345), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_345), .B(n_350), .Y(n_571) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NOR2x1_ASAP7_75t_L g1527 ( .A(n_349), .B(n_1528), .Y(n_1527) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g352 ( .A(n_350), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_350), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_350), .B(n_384), .Y(n_558) );
AOI22xp33_ASAP7_75t_SL g351 ( .A1(n_352), .A2(n_355), .B1(n_356), .B2(n_360), .Y(n_351) );
INVx1_ASAP7_75t_L g914 ( .A(n_352), .Y(n_914) );
BUFx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g564 ( .A(n_354), .Y(n_564) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_354), .B(n_1124), .Y(n_1133) );
INVx1_ASAP7_75t_L g1528 ( .A(n_354), .Y(n_1528) );
AND2x4_ASAP7_75t_L g1557 ( .A(n_354), .B(n_1124), .Y(n_1557) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g565 ( .A(n_357), .B(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g611 ( .A(n_357), .B(n_566), .Y(n_611) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_360), .A2(n_405), .B1(n_406), .B2(n_412), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_372), .B1(n_375), .B2(n_378), .Y(n_361) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g618 ( .A(n_364), .Y(n_618) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_367), .Y(n_584) );
BUFx3_ASAP7_75t_L g731 ( .A(n_367), .Y(n_731) );
AND2x4_ASAP7_75t_L g1113 ( .A(n_367), .B(n_1114), .Y(n_1113) );
INVx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g912 ( .A(n_371), .Y(n_912) );
INVx2_ASAP7_75t_L g1534 ( .A(n_371), .Y(n_1534) );
AND2x4_ASAP7_75t_L g573 ( .A(n_373), .B(n_574), .Y(n_573) );
AOI332xp33_ASAP7_75t_L g830 ( .A1(n_373), .A2(n_574), .A3(n_598), .B1(n_725), .B2(n_726), .B3(n_819), .C1(n_831), .C2(n_832), .Y(n_830) );
INVx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx4_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g540 ( .A(n_377), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_SL g769 ( .A(n_377), .B(n_399), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_377), .B(n_541), .Y(n_839) );
INVx4_ASAP7_75t_L g896 ( .A(n_377), .Y(n_896) );
BUFx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g616 ( .A(n_381), .Y(n_616) );
INVx1_ASAP7_75t_L g526 ( .A(n_382), .Y(n_526) );
BUFx2_ASAP7_75t_L g795 ( .A(n_382), .Y(n_795) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g466 ( .A(n_383), .B(n_467), .Y(n_466) );
AND2x4_ASAP7_75t_L g529 ( .A(n_383), .B(n_530), .Y(n_529) );
BUFx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g623 ( .A(n_384), .Y(n_623) );
NAND3xp33_ASAP7_75t_SL g385 ( .A(n_386), .B(n_404), .C(n_419), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_388), .A2(n_887), .B1(n_890), .B2(n_918), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g1495 ( .A1(n_388), .A2(n_918), .B1(n_1496), .B2(n_1497), .Y(n_1495) );
AND2x4_ASAP7_75t_L g388 ( .A(n_389), .B(n_397), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx8_ASAP7_75t_L g426 ( .A(n_390), .Y(n_426) );
INVx3_ASAP7_75t_L g490 ( .A(n_390), .Y(n_490) );
INVx2_ASAP7_75t_L g878 ( .A(n_390), .Y(n_878) );
INVx8_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2x1p5_ASAP7_75t_L g659 ( .A(n_391), .B(n_437), .Y(n_659) );
BUFx3_ASAP7_75t_L g687 ( .A(n_391), .Y(n_687) );
AND2x2_ASAP7_75t_L g691 ( .A(n_391), .B(n_692), .Y(n_691) );
BUFx3_ASAP7_75t_L g787 ( .A(n_391), .Y(n_787) );
AND2x4_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
AND2x4_ASAP7_75t_L g409 ( .A(n_392), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_393), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_393), .B(n_417), .Y(n_424) );
OR2x2_ASAP7_75t_L g447 ( .A(n_393), .B(n_395), .Y(n_447) );
AND2x4_ASAP7_75t_L g483 ( .A(n_393), .B(n_432), .Y(n_483) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVxp67_ASAP7_75t_L g410 ( .A(n_396), .Y(n_410) );
AND2x4_ASAP7_75t_L g918 ( .A(n_397), .B(n_648), .Y(n_918) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g411 ( .A(n_398), .Y(n_411) );
OR2x2_ASAP7_75t_L g413 ( .A(n_398), .B(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g421 ( .A(n_398), .B(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_402), .Y(n_398) );
OR2x2_ASAP7_75t_L g443 ( .A(n_399), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g542 ( .A(n_399), .Y(n_542) );
HB1xp67_ASAP7_75t_L g1174 ( .A(n_399), .Y(n_1174) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx2_ASAP7_75t_L g566 ( .A(n_400), .Y(n_566) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g476 ( .A(n_402), .Y(n_476) );
INVx1_ASAP7_75t_L g692 ( .A(n_402), .Y(n_692) );
INVx3_ASAP7_75t_L g438 ( .A(n_403), .Y(n_438) );
NAND2xp33_ASAP7_75t_SL g444 ( .A(n_403), .B(n_440), .Y(n_444) );
BUFx3_ASAP7_75t_L g524 ( .A(n_403), .Y(n_524) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_411), .Y(n_406) );
INVx2_ASAP7_75t_L g460 ( .A(n_407), .Y(n_460) );
INVx2_ASAP7_75t_L g821 ( .A(n_407), .Y(n_821) );
INVx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OR2x6_ASAP7_75t_SL g673 ( .A(n_408), .B(n_674), .Y(n_673) );
BUFx2_ASAP7_75t_L g868 ( .A(n_408), .Y(n_868) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_409), .Y(n_454) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_409), .Y(n_521) );
BUFx8_ASAP7_75t_L g648 ( .A(n_409), .Y(n_648) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g916 ( .A(n_413), .B(n_611), .Y(n_916) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_414), .Y(n_450) );
INVx4_ASAP7_75t_L g504 ( .A(n_414), .Y(n_504) );
INVx3_ASAP7_75t_L g781 ( .A(n_414), .Y(n_781) );
OAI221xp5_ASAP7_75t_L g805 ( .A1(n_414), .A2(n_523), .B1(n_806), .B2(n_807), .C(n_808), .Y(n_805) );
HB1xp67_ASAP7_75t_L g1092 ( .A(n_414), .Y(n_1092) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx3_ASAP7_75t_L g433 ( .A(n_415), .Y(n_433) );
BUFx2_ASAP7_75t_L g635 ( .A(n_415), .Y(n_635) );
NAND2x1p5_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
BUFx2_ASAP7_75t_L g1162 ( .A(n_416), .Y(n_1162) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g432 ( .A(n_417), .Y(n_432) );
INVx2_ASAP7_75t_L g428 ( .A(n_418), .Y(n_428) );
AND2x4_ASAP7_75t_L g479 ( .A(n_418), .B(n_431), .Y(n_479) );
BUFx2_ASAP7_75t_L g1159 ( .A(n_418), .Y(n_1159) );
NOR2xp33_ASAP7_75t_SL g419 ( .A(n_420), .B(n_441), .Y(n_419) );
AND2x4_ASAP7_75t_L g854 ( .A(n_421), .B(n_570), .Y(n_854) );
INVx1_ASAP7_75t_L g994 ( .A(n_422), .Y(n_994) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_423), .Y(n_653) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx2_ASAP7_75t_L g457 ( .A(n_424), .Y(n_457) );
INVx3_ASAP7_75t_L g632 ( .A(n_428), .Y(n_632) );
INVx2_ASAP7_75t_L g862 ( .A(n_429), .Y(n_862) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g629 ( .A(n_430), .B(n_437), .Y(n_629) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI22xp33_ASAP7_75t_L g463 ( .A1(n_433), .A2(n_446), .B1(n_464), .B2(n_465), .Y(n_463) );
OAI221xp5_ASAP7_75t_L g788 ( .A1(n_433), .A2(n_460), .B1(n_523), .B2(n_756), .C(n_761), .Y(n_788) );
OAI221xp5_ASAP7_75t_L g790 ( .A1(n_433), .A2(n_486), .B1(n_507), .B2(n_749), .C(n_762), .Y(n_790) );
INVx2_ASAP7_75t_L g1080 ( .A(n_433), .Y(n_1080) );
AND2x2_ASAP7_75t_L g859 ( .A(n_434), .B(n_632), .Y(n_859) );
AND2x4_ASAP7_75t_L g861 ( .A(n_434), .B(n_862), .Y(n_861) );
AND2x4_ASAP7_75t_L g864 ( .A(n_434), .B(n_655), .Y(n_864) );
AND2x4_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
OR2x2_ASAP7_75t_L g570 ( .A(n_435), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g725 ( .A(n_435), .Y(n_725) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g874 ( .A(n_436), .Y(n_874) );
INVx1_ASAP7_75t_L g493 ( .A(n_437), .Y(n_493) );
AND2x6_ASAP7_75t_L g631 ( .A(n_437), .B(n_632), .Y(n_631) );
AND2x4_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
NAND2x1p5_ASAP7_75t_L g467 ( .A(n_438), .B(n_468), .Y(n_467) );
NAND3x1_ASAP7_75t_L g873 ( .A(n_438), .B(n_468), .C(n_874), .Y(n_873) );
OR2x4_ASAP7_75t_L g1146 ( .A(n_438), .B(n_447), .Y(n_1146) );
INVx1_ASAP7_75t_L g1149 ( .A(n_438), .Y(n_1149) );
AND2x4_ASAP7_75t_L g1154 ( .A(n_438), .B(n_483), .Y(n_1154) );
OR2x6_ASAP7_75t_L g1169 ( .A(n_438), .B(n_457), .Y(n_1169) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g523 ( .A(n_440), .B(n_524), .Y(n_523) );
AND3x4_ASAP7_75t_L g881 ( .A(n_440), .B(n_524), .C(n_623), .Y(n_881) );
HB1xp67_ASAP7_75t_L g1172 ( .A(n_440), .Y(n_1172) );
OAI33xp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_445), .A3(n_451), .B1(n_459), .B2(n_463), .B3(n_466), .Y(n_441) );
BUFx4f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx8_ASAP7_75t_L g1075 ( .A(n_443), .Y(n_1075) );
BUFx2_ASAP7_75t_L g642 ( .A(n_444), .Y(n_642) );
OAI22xp33_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_448), .B1(n_449), .B2(n_450), .Y(n_445) );
OAI221xp5_ASAP7_75t_L g810 ( .A1(n_446), .A2(n_507), .B1(n_635), .B2(n_811), .C(n_812), .Y(n_810) );
INVx1_ASAP7_75t_L g962 ( .A(n_446), .Y(n_962) );
BUFx4f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g486 ( .A(n_447), .Y(n_486) );
BUFx3_ASAP7_75t_L g505 ( .A(n_447), .Y(n_505) );
INVx2_ASAP7_75t_L g512 ( .A(n_447), .Y(n_512) );
OR2x4_ASAP7_75t_L g1166 ( .A(n_447), .B(n_1149), .Y(n_1166) );
OAI221xp5_ASAP7_75t_L g1042 ( .A1(n_450), .A2(n_523), .B1(n_647), .B2(n_1043), .C(n_1044), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B1(n_455), .B2(n_458), .Y(n_451) );
INVx8_ASAP7_75t_L g641 ( .A(n_453), .Y(n_641) );
INVx5_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_SL g487 ( .A(n_454), .Y(n_487) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_454), .Y(n_498) );
INVx3_ASAP7_75t_L g814 ( .A(n_454), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_455), .A2(n_460), .B1(n_461), .B2(n_462), .Y(n_459) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx2_ASAP7_75t_L g515 ( .A(n_456), .Y(n_515) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g500 ( .A(n_457), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g1085 ( .A1(n_460), .A2(n_500), .B1(n_1086), .B2(n_1087), .Y(n_1085) );
INVx3_ASAP7_75t_L g507 ( .A(n_467), .Y(n_507) );
NAND4xp75_ASAP7_75t_L g470 ( .A(n_471), .B(n_527), .C(n_567), .D(n_577), .Y(n_470) );
OAI21x1_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_494), .B(n_525), .Y(n_471) );
OAI21xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_477), .B(n_488), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_474), .A2(n_596), .B1(n_650), .B2(n_656), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g778 ( .A1(n_474), .A2(n_658), .B1(n_773), .B2(n_779), .C(n_782), .Y(n_778) );
AOI221xp5_ASAP7_75t_L g818 ( .A1(n_474), .A2(n_658), .B1(n_819), .B2(n_820), .C(n_825), .Y(n_818) );
BUFx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g674 ( .A(n_476), .Y(n_674) );
AND2x4_ASAP7_75t_L g676 ( .A(n_476), .B(n_479), .Y(n_676) );
AOI221xp5_ASAP7_75t_SL g477 ( .A1(n_478), .A2(n_480), .B1(n_481), .B2(n_484), .C(n_485), .Y(n_477) );
BUFx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx12f_ASAP7_75t_L g638 ( .A(n_479), .Y(n_638) );
INVx5_ASAP7_75t_L g684 ( .A(n_479), .Y(n_684) );
BUFx3_ASAP7_75t_L g876 ( .A(n_479), .Y(n_876) );
BUFx2_ASAP7_75t_L g956 ( .A(n_479), .Y(n_956) );
AOI211xp5_ASAP7_75t_L g1562 ( .A1(n_481), .A2(n_1154), .B(n_1558), .C(n_1563), .Y(n_1562) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g869 ( .A(n_482), .Y(n_869) );
INVx2_ASAP7_75t_L g1500 ( .A(n_482), .Y(n_1500) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx3_ASAP7_75t_L g640 ( .A(n_483), .Y(n_640) );
BUFx2_ASAP7_75t_L g655 ( .A(n_483), .Y(n_655) );
AND2x2_ASAP7_75t_L g694 ( .A(n_483), .B(n_692), .Y(n_694) );
BUFx2_ASAP7_75t_L g1574 ( .A(n_483), .Y(n_1574) );
BUFx2_ASAP7_75t_L g1580 ( .A(n_483), .Y(n_1580) );
OAI221xp5_ASAP7_75t_L g1048 ( .A1(n_486), .A2(n_507), .B1(n_518), .B2(n_1049), .C(n_1050), .Y(n_1048) );
INVx1_ASAP7_75t_L g1201 ( .A(n_486), .Y(n_1201) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B(n_491), .C(n_492), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_490), .A2(n_592), .B1(n_612), .B2(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OR2x6_ASAP7_75t_L g634 ( .A(n_493), .B(n_635), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_501), .B1(n_508), .B2(n_516), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B1(n_499), .B2(n_500), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_496), .A2(n_509), .B1(n_533), .B2(n_535), .Y(n_532) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OAI221xp5_ASAP7_75t_L g543 ( .A1(n_499), .A2(n_517), .B1(n_544), .B2(n_546), .C(n_551), .Y(n_543) );
OAI221xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_503), .B1(n_505), .B2(n_506), .C(n_507), .Y(n_501) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g518 ( .A(n_504), .Y(n_518) );
INVx2_ASAP7_75t_L g682 ( .A(n_504), .Y(n_682) );
INVx2_ASAP7_75t_L g959 ( .A(n_504), .Y(n_959) );
OAI22xp33_ASAP7_75t_L g1076 ( .A1(n_505), .A2(n_1077), .B1(n_1078), .B2(n_1079), .Y(n_1076) );
OAI22xp33_ASAP7_75t_L g1090 ( .A1(n_505), .A2(n_1091), .B1(n_1092), .B2(n_1093), .Y(n_1090) );
OAI221xp5_ASAP7_75t_L g1247 ( .A1(n_505), .A2(n_507), .B1(n_998), .B2(n_1248), .C(n_1249), .Y(n_1247) );
INVx3_ASAP7_75t_L g644 ( .A(n_507), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_507), .B(n_700), .Y(n_699) );
OAI221xp5_ASAP7_75t_L g957 ( .A1(n_507), .A2(n_958), .B1(n_959), .B2(n_960), .C(n_961), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_507), .B(n_1204), .Y(n_1203) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B1(n_513), .B2(n_514), .Y(n_508) );
BUFx4f_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g1045 ( .A1(n_511), .A2(n_793), .B1(n_1046), .B2(n_1047), .Y(n_1045) );
INVx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OAI221xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B1(n_519), .B2(n_522), .C(n_523), .Y(n_516) );
OAI21xp33_ASAP7_75t_L g988 ( .A1(n_518), .A2(n_989), .B(n_990), .Y(n_988) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g651 ( .A(n_521), .Y(n_651) );
INVx1_ASAP7_75t_L g680 ( .A(n_521), .Y(n_680) );
INVx2_ASAP7_75t_L g808 ( .A(n_521), .Y(n_808) );
BUFx6f_ASAP7_75t_L g955 ( .A(n_521), .Y(n_955) );
AND2x4_ASAP7_75t_L g1148 ( .A(n_521), .B(n_1149), .Y(n_1148) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_523), .A2(n_684), .B1(n_685), .B2(n_686), .C(n_688), .Y(n_683) );
OAI221xp5_ASAP7_75t_L g964 ( .A1(n_523), .A2(n_940), .B1(n_959), .B2(n_965), .C(n_966), .Y(n_964) );
INVx1_ASAP7_75t_L g1195 ( .A(n_523), .Y(n_1195) );
OAI221xp5_ASAP7_75t_L g1240 ( .A1(n_523), .A2(n_998), .B1(n_1241), .B2(n_1242), .C(n_1243), .Y(n_1240) );
INVx3_ASAP7_75t_L g1158 ( .A(n_524), .Y(n_1158) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AOI211x1_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_531), .B(n_538), .C(n_559), .Y(n_527) );
AOI222xp33_ASAP7_75t_L g1260 ( .A1(n_528), .A2(n_540), .B1(n_724), .B2(n_1261), .C1(n_1265), .C2(n_1269), .Y(n_1260) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AOI31xp33_ASAP7_75t_L g601 ( .A1(n_529), .A2(n_602), .A3(n_604), .B(n_606), .Y(n_601) );
INVx2_ASAP7_75t_L g722 ( .A(n_529), .Y(n_722) );
INVx2_ASAP7_75t_L g746 ( .A(n_529), .Y(n_746) );
INVx4_ASAP7_75t_L g944 ( .A(n_529), .Y(n_944) );
INVx1_ASAP7_75t_L g1095 ( .A(n_529), .Y(n_1095) );
INVx2_ASAP7_75t_L g1584 ( .A(n_529), .Y(n_1584) );
BUFx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx3_ASAP7_75t_L g733 ( .A(n_534), .Y(n_733) );
BUFx6f_ASAP7_75t_L g936 ( .A(n_534), .Y(n_936) );
INVx2_ASAP7_75t_SL g1022 ( .A(n_534), .Y(n_1022) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_535), .A2(n_758), .B1(n_761), .B2(n_762), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g1016 ( .A1(n_535), .A2(n_544), .B1(n_992), .B2(n_1017), .Y(n_1016) );
BUFx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g576 ( .A(n_536), .B(n_575), .Y(n_576) );
OR2x2_ASAP7_75t_L g599 ( .A(n_536), .B(n_575), .Y(n_599) );
INVx2_ASAP7_75t_SL g1105 ( .A(n_536), .Y(n_1105) );
BUFx3_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_537), .Y(n_555) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_543), .B(n_554), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_540), .Y(n_539) );
NAND3xp33_ASAP7_75t_L g613 ( .A(n_540), .B(n_614), .C(n_617), .Y(n_613) );
AOI322xp5_ASAP7_75t_L g712 ( .A1(n_540), .A2(n_713), .A3(n_716), .B1(n_721), .B2(n_723), .C1(n_724), .C2(n_727), .Y(n_712) );
AOI332xp33_ASAP7_75t_L g1061 ( .A1(n_540), .A2(n_724), .A3(n_1062), .B1(n_1063), .B2(n_1064), .B3(n_1065), .C1(n_1066), .C2(n_1068), .Y(n_1061) );
INVx2_ASAP7_75t_L g1106 ( .A(n_540), .Y(n_1106) );
AOI33xp33_ASAP7_75t_L g1581 ( .A1(n_540), .A2(n_1582), .A3(n_1585), .B1(n_1588), .B2(n_1589), .B3(n_1593), .Y(n_1581) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g1096 ( .A1(n_546), .A2(n_1077), .B1(n_1091), .B2(n_1097), .Y(n_1096) );
OAI221xp5_ASAP7_75t_L g1529 ( .A1(n_546), .A2(n_1530), .B1(n_1531), .B2(n_1532), .C(n_1533), .Y(n_1529) );
INVx6_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx5_ASAP7_75t_L g720 ( .A(n_547), .Y(n_720) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g735 ( .A(n_548), .Y(n_735) );
INVx2_ASAP7_75t_SL g750 ( .A(n_548), .Y(n_750) );
INVx4_ASAP7_75t_L g929 ( .A(n_548), .Y(n_929) );
INVx2_ASAP7_75t_L g943 ( .A(n_548), .Y(n_943) );
INVx1_ASAP7_75t_L g1109 ( .A(n_548), .Y(n_1109) );
INVx8_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx2_ASAP7_75t_L g1015 ( .A(n_549), .Y(n_1015) );
OR2x2_ASAP7_75t_L g1123 ( .A(n_549), .B(n_1124), .Y(n_1123) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g898 ( .A(n_553), .Y(n_898) );
INVx1_ASAP7_75t_L g905 ( .A(n_553), .Y(n_905) );
INVx2_ASAP7_75t_SL g1067 ( .A(n_553), .Y(n_1067) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_554), .Y(n_606) );
OR2x6_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
INVx4_ASAP7_75t_L g754 ( .A(n_555), .Y(n_754) );
BUFx4f_ASAP7_75t_L g837 ( .A(n_555), .Y(n_837) );
BUFx6f_ASAP7_75t_L g842 ( .A(n_555), .Y(n_842) );
BUFx4f_ASAP7_75t_L g1128 ( .A(n_555), .Y(n_1128) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2x2_ASAP7_75t_L g562 ( .A(n_557), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g608 ( .A(n_562), .Y(n_608) );
HB1xp67_ASAP7_75t_L g1259 ( .A(n_562), .Y(n_1259) );
INVx2_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g579 ( .A(n_566), .Y(n_579) );
INVxp67_ASAP7_75t_L g851 ( .A(n_566), .Y(n_851) );
INVx1_ASAP7_75t_L g1141 ( .A(n_566), .Y(n_1141) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g726 ( .A(n_571), .Y(n_726) );
INVxp67_ASAP7_75t_L g1209 ( .A(n_572), .Y(n_1209) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_573), .A2(n_596), .B1(n_597), .B2(n_598), .Y(n_595) );
AOI222xp33_ASAP7_75t_L g771 ( .A1(n_573), .A2(n_598), .B1(n_724), .B2(n_772), .C1(n_773), .C2(n_774), .Y(n_771) );
AOI222xp33_ASAP7_75t_L g945 ( .A1(n_573), .A2(n_598), .B1(n_724), .B2(n_946), .C1(n_947), .C2(n_948), .Y(n_945) );
AOI222xp33_ASAP7_75t_L g1026 ( .A1(n_573), .A2(n_598), .B1(n_724), .B2(n_985), .C1(n_1004), .C2(n_1027), .Y(n_1026) );
AOI21xp33_ASAP7_75t_L g1058 ( .A1(n_573), .A2(n_1059), .B(n_1060), .Y(n_1058) );
AOI211xp5_ASAP7_75t_L g1256 ( .A1(n_573), .A2(n_1233), .B(n_1257), .C(n_1258), .Y(n_1256) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_SL g577 ( .A1(n_578), .A2(n_581), .B1(n_582), .B2(n_585), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_578), .B(n_592), .Y(n_591) );
AOI211xp5_ASAP7_75t_L g705 ( .A1(n_578), .A2(n_706), .B(n_707), .C(n_711), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_578), .B(n_776), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_578), .B(n_824), .Y(n_828) );
INVx3_ASAP7_75t_L g922 ( .A(n_578), .Y(n_922) );
AO211x2_ASAP7_75t_L g1179 ( .A1(n_578), .A2(n_1180), .B(n_1181), .C(n_1207), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1270 ( .A(n_578), .B(n_1271), .Y(n_1270) );
AND2x4_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
AND2x4_ASAP7_75t_L g582 ( .A(n_579), .B(n_583), .Y(n_582) );
BUFx6f_ASAP7_75t_L g889 ( .A(n_580), .Y(n_889) );
INVx1_ASAP7_75t_L g1519 ( .A(n_580), .Y(n_1519) );
INVx1_ASAP7_75t_L g661 ( .A(n_582), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_582), .B(n_703), .Y(n_702) );
NAND2xp33_ASAP7_75t_SL g796 ( .A(n_582), .B(n_797), .Y(n_796) );
HB1xp67_ASAP7_75t_L g973 ( .A(n_582), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_582), .B(n_1003), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_582), .B(n_1057), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_582), .B(n_1206), .Y(n_1205) );
INVx1_ASAP7_75t_L g1254 ( .A(n_582), .Y(n_1254) );
BUFx6f_ASAP7_75t_L g715 ( .A(n_584), .Y(n_715) );
INVx2_ASAP7_75t_L g911 ( .A(n_584), .Y(n_911) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_664), .B1(n_665), .B2(n_736), .Y(n_586) );
INVx1_ASAP7_75t_L g736 ( .A(n_587), .Y(n_736) );
OAI21x1_ASAP7_75t_SL g587 ( .A1(n_588), .A2(n_589), .B(n_663), .Y(n_587) );
NAND4xp25_ASAP7_75t_L g663 ( .A(n_588), .B(n_591), .C(n_593), .D(n_622), .Y(n_663) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND3xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .C(n_622), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_594), .B(n_600), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g1055 ( .A1(n_598), .A2(n_606), .B(n_1040), .Y(n_1055) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND3xp33_ASAP7_75t_SL g600 ( .A(n_601), .B(n_607), .C(n_613), .Y(n_600) );
AOI222xp33_ASAP7_75t_L g1554 ( .A1(n_603), .A2(n_1555), .B1(n_1556), .B2(n_1557), .C1(n_1558), .C2(n_1559), .Y(n_1554) );
NOR3xp33_ASAP7_75t_L g833 ( .A(n_606), .B(n_834), .C(n_844), .Y(n_833) );
NOR3xp33_ASAP7_75t_L g923 ( .A(n_606), .B(n_924), .C(n_925), .Y(n_923) );
AOI21xp33_ASAP7_75t_L g1226 ( .A1(n_606), .A2(n_724), .B(n_1227), .Y(n_1226) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_608), .A2(n_609), .B1(n_610), .B2(n_612), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_608), .A2(n_610), .B1(n_709), .B2(n_710), .Y(n_708) );
AOI222xp33_ASAP7_75t_L g1208 ( .A1(n_608), .A2(n_610), .B1(n_1183), .B2(n_1209), .C1(n_1210), .C2(n_1211), .Y(n_1208) );
INVx2_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g1262 ( .A(n_620), .Y(n_1262) );
BUFx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g1592 ( .A(n_621), .Y(n_1592) );
AOI22xp33_ASAP7_75t_SL g622 ( .A1(n_623), .A2(n_624), .B1(n_660), .B2(n_662), .Y(n_622) );
INVx2_ASAP7_75t_SL g701 ( .A(n_623), .Y(n_701) );
INVx1_ASAP7_75t_L g827 ( .A(n_623), .Y(n_827) );
OAI31xp33_ASAP7_75t_SL g1032 ( .A1(n_623), .A2(n_1033), .A3(n_1037), .B(n_1041), .Y(n_1032) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_636), .C(n_649), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_633), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g671 ( .A(n_629), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_629), .A2(n_631), .B1(n_1039), .B2(n_1040), .Y(n_1038) );
INVx4_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NOR3xp33_ASAP7_75t_L g783 ( .A(n_633), .B(n_784), .C(n_789), .Y(n_783) );
NOR3xp33_ASAP7_75t_L g803 ( .A(n_633), .B(n_804), .C(n_809), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g698 ( .A(n_635), .Y(n_698) );
INVx1_ASAP7_75t_L g1152 ( .A(n_635), .Y(n_1152) );
INVx1_ASAP7_75t_L g1202 ( .A(n_635), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_639), .B1(n_643), .B2(n_645), .Y(n_636) );
BUFx2_ASAP7_75t_L g883 ( .A(n_638), .Y(n_883) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_647), .A2(n_993), .B1(n_1052), .B2(n_1053), .Y(n_1051) );
INVx3_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx3_ASAP7_75t_L g792 ( .A(n_648), .Y(n_792) );
INVx2_ASAP7_75t_SL g966 ( .A(n_648), .Y(n_966) );
INVx2_ASAP7_75t_SL g1242 ( .A(n_648), .Y(n_1242) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_652), .A2(n_1082), .B1(n_1083), .B2(n_1084), .Y(n_1081) );
CKINVDCx8_ASAP7_75t_R g652 ( .A(n_653), .Y(n_652) );
INVx3_ASAP7_75t_L g793 ( .A(n_653), .Y(n_793) );
INVx3_ASAP7_75t_L g816 ( .A(n_653), .Y(n_816) );
BUFx2_ASAP7_75t_L g1507 ( .A(n_655), .Y(n_1507) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI211xp5_ASAP7_75t_SL g668 ( .A1(n_658), .A2(n_669), .B(n_670), .C(n_672), .Y(n_668) );
AOI211xp5_ASAP7_75t_SL g950 ( .A1(n_658), .A2(n_946), .B(n_951), .C(n_952), .Y(n_950) );
AOI211xp5_ASAP7_75t_L g984 ( .A1(n_658), .A2(n_985), .B(n_986), .C(n_987), .Y(n_984) );
AOI211xp5_ASAP7_75t_SL g1182 ( .A1(n_658), .A2(n_1183), .B(n_1184), .C(n_1185), .Y(n_1182) );
AOI211xp5_ASAP7_75t_L g1232 ( .A1(n_658), .A2(n_1233), .B(n_1234), .C(n_1235), .Y(n_1232) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OR2x6_ASAP7_75t_L g850 ( .A(n_659), .B(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NOR2x1_ASAP7_75t_L g666 ( .A(n_667), .B(n_704), .Y(n_666) );
A2O1A1Ixp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_677), .B(n_701), .C(n_702), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g1002 ( .A(n_673), .Y(n_1002) );
INVx3_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI221xp5_ASAP7_75t_L g1001 ( .A1(n_676), .A2(n_1002), .B1(n_1003), .B2(n_1004), .C(n_1005), .Y(n_1001) );
NOR3xp33_ASAP7_75t_SL g677 ( .A(n_678), .B(n_689), .C(n_695), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx2_ASAP7_75t_R g1246 ( .A(n_684), .Y(n_1246) );
INVx1_ASAP7_75t_L g1502 ( .A(n_684), .Y(n_1502) );
INVx2_ASAP7_75t_L g1505 ( .A(n_684), .Y(n_1505) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_685), .A2(n_733), .B1(n_734), .B2(n_735), .Y(n_732) );
INVx2_ASAP7_75t_L g1239 ( .A(n_686), .Y(n_1239) );
INVx2_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_687), .B(n_824), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_688), .A2(n_718), .B1(n_719), .B2(n_720), .Y(n_717) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g1034 ( .A1(n_691), .A2(n_694), .B1(n_1035), .B2(n_1036), .Y(n_1034) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_712), .Y(n_704) );
BUFx3_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_718), .A2(n_748), .B1(n_749), .B2(n_750), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g1221 ( .A1(n_718), .A2(n_720), .B1(n_1222), .B2(n_1223), .Y(n_1221) );
OAI22xp5_ASAP7_75t_L g1266 ( .A1(n_718), .A2(n_1015), .B1(n_1267), .B2(n_1268), .Y(n_1266) );
AND2x4_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
BUFx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
BUFx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
XNOR2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_845), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
XNOR2x1_ASAP7_75t_L g739 ( .A(n_740), .B(n_798), .Y(n_739) );
XNOR2x1_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
NOR2x1_ASAP7_75t_L g742 ( .A(n_743), .B(n_777), .Y(n_742) );
NAND3xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_771), .C(n_775), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_770), .Y(n_744) );
OAI33xp33_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_747), .A3(n_751), .B1(n_757), .B2(n_763), .B3(n_768), .Y(n_745) );
OAI22xp5_ASAP7_75t_SL g834 ( .A1(n_746), .A2(n_835), .B1(n_839), .B2(n_840), .Y(n_834) );
OAI33xp33_ASAP7_75t_L g1011 ( .A1(n_746), .A2(n_1012), .A3(n_1016), .B1(n_1018), .B2(n_1020), .B3(n_1024), .Y(n_1011) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_750), .A2(n_764), .B1(n_766), .B2(n_767), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_753), .B1(n_755), .B2(n_756), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_752), .A2(n_767), .B1(n_792), .B2(n_793), .Y(n_791) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g934 ( .A(n_754), .Y(n_934) );
INVx4_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
BUFx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g841 ( .A(n_760), .Y(n_841) );
INVx2_ASAP7_75t_L g1100 ( .A(n_760), .Y(n_1100) );
OAI22xp33_ASAP7_75t_L g1263 ( .A1(n_764), .A2(n_1015), .B1(n_1249), .B2(n_1264), .Y(n_1263) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx2_ASAP7_75t_L g1024 ( .A(n_769), .Y(n_1024) );
A2O1A1Ixp33_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_783), .B(n_794), .C(n_796), .Y(n_777) );
INVx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g822 ( .A(n_781), .Y(n_822) );
INVx3_ASAP7_75t_L g998 ( .A(n_781), .Y(n_998) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
BUFx2_ASAP7_75t_L g1573 ( .A(n_787), .Y(n_1573) );
INVx1_ASAP7_75t_L g1504 ( .A(n_792), .Y(n_1504) );
AOI21xp5_ASAP7_75t_L g884 ( .A1(n_794), .A2(n_885), .B(n_915), .Y(n_884) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g1250 ( .A(n_795), .Y(n_1250) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
XNOR2x1_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
OR2x2_ASAP7_75t_L g801 ( .A(n_802), .B(n_829), .Y(n_801) );
A2O1A1Ixp33_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_818), .B(n_826), .C(n_828), .Y(n_802) );
OAI221xp5_ASAP7_75t_L g840 ( .A1(n_806), .A2(n_811), .B1(n_841), .B2(n_842), .C(n_843), .Y(n_840) );
OAI221xp5_ASAP7_75t_L g835 ( .A1(n_807), .A2(n_815), .B1(n_836), .B2(n_837), .C(n_838), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_815), .B1(n_816), .B2(n_817), .Y(n_813) );
A2O1A1Ixp33_ASAP7_75t_SL g1181 ( .A1(n_826), .A2(n_1182), .B(n_1186), .C(n_1205), .Y(n_1181) );
HB1xp67_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
BUFx2_ASAP7_75t_L g970 ( .A(n_827), .Y(n_970) );
INVx2_ASAP7_75t_L g931 ( .A(n_836), .Y(n_931) );
OAI221xp5_ASAP7_75t_L g937 ( .A1(n_837), .A2(n_938), .B1(n_939), .B2(n_940), .C(n_941), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g1099 ( .A1(n_837), .A2(n_1082), .B1(n_1086), .B2(n_1100), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_842), .A2(n_989), .B1(n_997), .B2(n_1019), .Y(n_1018) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_919), .B1(n_975), .B2(n_976), .Y(n_845) );
INVx1_ASAP7_75t_L g976 ( .A(n_846), .Y(n_976) );
NAND2xp67_ASAP7_75t_L g847 ( .A(n_848), .B(n_884), .Y(n_847) );
AOI221xp5_ASAP7_75t_L g848 ( .A1(n_849), .A2(n_852), .B1(n_853), .B2(n_855), .C(n_856), .Y(n_848) );
INVx3_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
AOI221xp5_ASAP7_75t_L g893 ( .A1(n_852), .A2(n_894), .B1(n_895), .B2(n_897), .C(n_900), .Y(n_893) );
INVx8_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
NAND3xp33_ASAP7_75t_SL g856 ( .A(n_857), .B(n_863), .C(n_865), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_858), .A2(n_859), .B1(n_860), .B2(n_861), .Y(n_857) );
AOI222xp33_ASAP7_75t_L g901 ( .A1(n_858), .A2(n_860), .B1(n_902), .B2(n_904), .C1(n_906), .C2(n_913), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g1492 ( .A1(n_859), .A2(n_861), .B1(n_1493), .B2(n_1494), .Y(n_1492) );
INVx3_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
NOR3xp33_ASAP7_75t_L g1490 ( .A(n_864), .B(n_1491), .C(n_1508), .Y(n_1490) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_866), .A2(n_870), .B1(n_877), .B2(n_882), .Y(n_865) );
INVx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
AND2x2_ASAP7_75t_L g870 ( .A(n_871), .B(n_875), .Y(n_870) );
BUFx2_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
BUFx2_ASAP7_75t_L g1577 ( .A(n_872), .Y(n_1577) );
INVx3_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx3_ASAP7_75t_L g1089 ( .A(n_873), .Y(n_1089) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
AOI33xp33_ASAP7_75t_L g1498 ( .A1(n_880), .A2(n_1089), .A3(n_1499), .B1(n_1501), .B2(n_1503), .B3(n_1506), .Y(n_1498) );
AOI33xp33_ASAP7_75t_L g1571 ( .A1(n_880), .A2(n_1572), .A3(n_1575), .B1(n_1576), .B2(n_1577), .B3(n_1578), .Y(n_1571) );
BUFx3_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
NAND3xp33_ASAP7_75t_SL g885 ( .A(n_886), .B(n_893), .C(n_901), .Y(n_885) );
AOI22xp5_ASAP7_75t_L g886 ( .A1(n_887), .A2(n_888), .B1(n_890), .B2(n_891), .Y(n_886) );
HB1xp67_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
BUFx6f_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g1521 ( .A(n_892), .Y(n_1521) );
INVx3_ASAP7_75t_L g1511 ( .A(n_894), .Y(n_1511) );
AOI21xp5_ASAP7_75t_SL g1512 ( .A1(n_900), .A2(n_1513), .B(n_1516), .Y(n_1512) );
BUFx3_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx2_ASAP7_75t_L g1525 ( .A(n_903), .Y(n_1525) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
HB1xp67_ASAP7_75t_L g1220 ( .A(n_910), .Y(n_1220) );
INVx2_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g975 ( .A(n_919), .Y(n_975) );
XOR2x2_ASAP7_75t_L g919 ( .A(n_920), .B(n_974), .Y(n_919) );
NOR2x1_ASAP7_75t_SL g920 ( .A(n_921), .B(n_949), .Y(n_920) );
INVx1_ASAP7_75t_L g1008 ( .A(n_922), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_926), .B(n_937), .Y(n_925) );
OAI211xp5_ASAP7_75t_L g926 ( .A1(n_927), .A2(n_928), .B(n_930), .C(n_932), .Y(n_926) );
HB1xp67_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
INVx3_ASAP7_75t_L g939 ( .A(n_931), .Y(n_939) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
INVx2_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g1012 ( .A1(n_936), .A2(n_1013), .B1(n_1014), .B2(n_1015), .Y(n_1012) );
INVxp33_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx2_ASAP7_75t_SL g1064 ( .A(n_944), .Y(n_1064) );
INVx2_ASAP7_75t_SL g1217 ( .A(n_944), .Y(n_1217) );
A2O1A1Ixp33_ASAP7_75t_SL g949 ( .A1(n_950), .A2(n_953), .B(n_968), .C(n_971), .Y(n_949) );
NOR3xp33_ASAP7_75t_L g953 ( .A(n_954), .B(n_963), .C(n_967), .Y(n_953) );
INVx1_ASAP7_75t_L g1083 ( .A(n_955), .Y(n_1083) );
INVx1_ASAP7_75t_L g1190 ( .A(n_955), .Y(n_1190) );
INVx2_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_966), .A2(n_992), .B1(n_993), .B2(n_995), .Y(n_991) );
OAI21xp5_ASAP7_75t_L g1509 ( .A1(n_968), .A2(n_1510), .B(n_1522), .Y(n_1509) );
INVx2_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
A2O1A1Ixp33_ASAP7_75t_SL g983 ( .A1(n_970), .A2(n_984), .B(n_1001), .C(n_1006), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_972), .B(n_973), .Y(n_971) );
INVxp67_ASAP7_75t_SL g1275 ( .A(n_977), .Y(n_1275) );
XNOR2xp5_ASAP7_75t_L g977 ( .A(n_978), .B(n_1070), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
XNOR2xp5_ASAP7_75t_L g980 ( .A(n_981), .B(n_1029), .Y(n_980) );
OR2x2_ASAP7_75t_L g982 ( .A(n_983), .B(n_1009), .Y(n_982) );
OAI21xp33_ASAP7_75t_L g987 ( .A1(n_988), .A2(n_991), .B(n_996), .Y(n_987) );
INVx1_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
OAI22xp5_ASAP7_75t_L g1020 ( .A1(n_995), .A2(n_1015), .B1(n_1021), .B2(n_1023), .Y(n_1020) );
OAI211xp5_ASAP7_75t_L g996 ( .A1(n_997), .A2(n_998), .B(n_999), .C(n_1000), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1008), .Y(n_1006) );
NAND3xp33_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1026), .C(n_1028), .Y(n_1009) );
NOR2xp33_ASAP7_75t_SL g1010 ( .A(n_1011), .B(n_1025), .Y(n_1010) );
INVx2_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
XOR2x2_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1069), .Y(n_1029) );
NOR2xp33_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1054), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_1042), .A2(n_1045), .B1(n_1048), .B2(n_1051), .Y(n_1041) );
NAND4xp25_ASAP7_75t_SL g1054 ( .A(n_1055), .B(n_1056), .C(n_1058), .D(n_1061), .Y(n_1054) );
XNOR2xp5_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1176), .Y(n_1070) );
XOR2x2_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1175), .Y(n_1071) );
AND3x1_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1110), .C(n_1142), .Y(n_1072) );
NOR2xp33_ASAP7_75t_SL g1073 ( .A(n_1074), .B(n_1094), .Y(n_1073) );
OAI33xp33_ASAP7_75t_L g1074 ( .A1(n_1075), .A2(n_1076), .A3(n_1081), .B1(n_1085), .B2(n_1088), .B3(n_1090), .Y(n_1074) );
OAI22xp5_ASAP7_75t_L g1101 ( .A1(n_1078), .A2(n_1093), .B1(n_1102), .B2(n_1104), .Y(n_1101) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_1084), .A2(n_1087), .B1(n_1097), .B2(n_1108), .Y(n_1107) );
INVx2_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1092), .Y(n_1193) );
OAI33xp33_ASAP7_75t_L g1094 ( .A1(n_1095), .A2(n_1096), .A3(n_1099), .B1(n_1101), .B2(n_1106), .B3(n_1107), .Y(n_1094) );
INVx2_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
INVx2_ASAP7_75t_L g1530 ( .A(n_1098), .Y(n_1530) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1100), .Y(n_1103) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
INVx5_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
BUFx3_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
OAI31xp33_ASAP7_75t_L g1110 ( .A1(n_1111), .A2(n_1115), .A3(n_1125), .B(n_1139), .Y(n_1110) );
INVx4_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
INVx2_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
INVx2_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
INVx2_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g1547 ( .A1(n_1122), .A2(n_1548), .B1(n_1549), .B2(n_1550), .Y(n_1547) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
NAND4xp25_ASAP7_75t_L g1546 ( .A(n_1129), .B(n_1547), .C(n_1551), .D(n_1554), .Y(n_1546) );
INVx3_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_1133), .A2(n_1134), .B1(n_1135), .B2(n_1138), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_1134), .A2(n_1156), .B1(n_1160), .B2(n_1163), .Y(n_1155) );
INVx2_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
INVx2_ASAP7_75t_L g1559 ( .A(n_1136), .Y(n_1559) );
INVx2_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
BUFx3_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
AOI22xp5_ASAP7_75t_L g1545 ( .A1(n_1140), .A2(n_1546), .B1(n_1560), .B2(n_1561), .Y(n_1545) );
OAI31xp33_ASAP7_75t_L g1142 ( .A1(n_1143), .A2(n_1150), .A3(n_1164), .B(n_1170), .Y(n_1142) );
INVx2_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g1570 ( .A1(n_1145), .A2(n_1148), .B1(n_1552), .B2(n_1553), .Y(n_1570) );
INVx2_ASAP7_75t_SL g1145 ( .A(n_1146), .Y(n_1145) );
INVx2_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
INVxp67_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
CKINVDCx8_ASAP7_75t_R g1153 ( .A(n_1154), .Y(n_1153) );
BUFx3_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1159), .Y(n_1157) );
AND2x4_ASAP7_75t_L g1161 ( .A(n_1158), .B(n_1162), .Y(n_1161) );
AND2x4_ASAP7_75t_L g1565 ( .A(n_1158), .B(n_1159), .Y(n_1565) );
BUFx6f_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1161), .Y(n_1566) );
BUFx2_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
BUFx3_ASAP7_75t_L g1569 ( .A(n_1166), .Y(n_1569) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
AOI22xp33_ASAP7_75t_L g1567 ( .A1(n_1168), .A2(n_1548), .B1(n_1550), .B2(n_1568), .Y(n_1567) );
INVx2_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
AND2x2_ASAP7_75t_SL g1170 ( .A(n_1171), .B(n_1173), .Y(n_1170) );
AND2x4_ASAP7_75t_L g1560 ( .A(n_1171), .B(n_1173), .Y(n_1560) );
INVx1_ASAP7_75t_SL g1171 ( .A(n_1172), .Y(n_1171) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
AOI22xp5_ASAP7_75t_L g1176 ( .A1(n_1177), .A2(n_1228), .B1(n_1272), .B2(n_1273), .Y(n_1176) );
HB1xp67_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
INVx2_ASAP7_75t_L g1272 ( .A(n_1178), .Y(n_1272) );
NOR3xp33_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1197), .C(n_1198), .Y(n_1186) );
NOR3xp33_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1191), .C(n_1196), .Y(n_1187) );
NOR2xp33_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1190), .Y(n_1188) );
NOR2xp33_ASAP7_75t_L g1219 ( .A(n_1189), .B(n_1215), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1194), .Y(n_1191) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
INVx2_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
NAND3xp33_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1212), .C(n_1226), .Y(n_1207) );
AOI22xp5_ASAP7_75t_L g1212 ( .A1(n_1213), .A2(n_1218), .B1(n_1224), .B2(n_1225), .Y(n_1212) );
AOI22xp5_ASAP7_75t_L g1218 ( .A1(n_1214), .A2(n_1219), .B1(n_1220), .B2(n_1221), .Y(n_1218) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1228), .Y(n_1273) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
OR2x2_ASAP7_75t_L g1230 ( .A(n_1231), .B(n_1255), .Y(n_1230) );
A2O1A1Ixp33_ASAP7_75t_SL g1231 ( .A1(n_1232), .A2(n_1236), .B(n_1250), .C(n_1251), .Y(n_1231) );
NOR3xp33_ASAP7_75t_L g1236 ( .A(n_1237), .B(n_1244), .C(n_1245), .Y(n_1236) );
BUFx2_ASAP7_75t_SL g1238 ( .A(n_1239), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1252), .B(n_1253), .Y(n_1251) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
NAND3xp33_ASAP7_75t_L g1255 ( .A(n_1256), .B(n_1260), .C(n_1270), .Y(n_1255) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1262), .Y(n_1515) );
OAI221xp5_ASAP7_75t_L g1276 ( .A1(n_1277), .A2(n_1483), .B1(n_1487), .B2(n_1535), .C(n_1538), .Y(n_1276) );
NOR2xp67_ASAP7_75t_L g1277 ( .A(n_1278), .B(n_1430), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1394), .Y(n_1278) );
O2A1O1Ixp33_ASAP7_75t_SL g1279 ( .A1(n_1280), .A2(n_1331), .B(n_1360), .C(n_1368), .Y(n_1279) );
O2A1O1Ixp33_ASAP7_75t_L g1280 ( .A1(n_1281), .A2(n_1297), .B(n_1310), .C(n_1326), .Y(n_1280) );
INVx2_ASAP7_75t_L g1313 ( .A(n_1281), .Y(n_1313) );
NAND2xp5_ASAP7_75t_L g1357 ( .A(n_1281), .B(n_1353), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1281), .B(n_1337), .Y(n_1382) );
AND2x2_ASAP7_75t_L g1397 ( .A(n_1281), .B(n_1398), .Y(n_1397) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1281), .B(n_1338), .Y(n_1406) );
OAI221xp5_ASAP7_75t_L g1463 ( .A1(n_1281), .A2(n_1313), .B1(n_1464), .B2(n_1466), .C(n_1468), .Y(n_1463) );
INVx2_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_1282), .B(n_1328), .Y(n_1410) );
NAND2xp5_ASAP7_75t_L g1439 ( .A(n_1282), .B(n_1319), .Y(n_1439) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1283), .B(n_1336), .Y(n_1335) );
OR2x2_ASAP7_75t_L g1344 ( .A(n_1283), .B(n_1328), .Y(n_1344) );
AND2x2_ASAP7_75t_L g1386 ( .A(n_1283), .B(n_1328), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1419 ( .A(n_1283), .B(n_1319), .Y(n_1419) );
OR2x2_ASAP7_75t_L g1444 ( .A(n_1283), .B(n_1319), .Y(n_1444) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1284), .B(n_1291), .Y(n_1283) );
INVx2_ASAP7_75t_L g1365 ( .A(n_1285), .Y(n_1365) );
AND2x6_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1287), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1286), .B(n_1290), .Y(n_1289) );
AND2x4_ASAP7_75t_L g1292 ( .A(n_1286), .B(n_1293), .Y(n_1292) );
AND2x6_ASAP7_75t_L g1295 ( .A(n_1286), .B(n_1296), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1286), .B(n_1290), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1286), .B(n_1290), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1288), .B(n_1294), .Y(n_1293) );
INVxp67_ASAP7_75t_L g1367 ( .A(n_1289), .Y(n_1367) );
HB1xp67_ASAP7_75t_L g1486 ( .A(n_1289), .Y(n_1486) );
OAI21xp5_ASAP7_75t_L g1596 ( .A1(n_1290), .A2(n_1597), .B(n_1598), .Y(n_1596) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1297), .Y(n_1401) );
OR2x2_ASAP7_75t_L g1297 ( .A(n_1298), .B(n_1302), .Y(n_1297) );
BUFx2_ASAP7_75t_L g1318 ( .A(n_1298), .Y(n_1318) );
INVx2_ASAP7_75t_L g1352 ( .A(n_1298), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1298), .B(n_1399), .Y(n_1398) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1298), .B(n_1323), .Y(n_1408) );
AOI222xp33_ASAP7_75t_L g1468 ( .A1(n_1298), .A2(n_1398), .B1(n_1410), .B2(n_1418), .C1(n_1469), .C2(n_1470), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1299), .B(n_1300), .Y(n_1298) );
OAI221xp5_ASAP7_75t_L g1331 ( .A1(n_1302), .A2(n_1332), .B1(n_1342), .B2(n_1345), .C(n_1347), .Y(n_1331) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1380 ( .A(n_1303), .B(n_1351), .Y(n_1380) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_1303), .B(n_1317), .Y(n_1465) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_1303), .B(n_1353), .Y(n_1467) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1307), .Y(n_1303) );
INVx2_ASAP7_75t_L g1324 ( .A(n_1304), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_1304), .B(n_1325), .Y(n_1399) );
OAI222xp33_ASAP7_75t_L g1457 ( .A1(n_1304), .A2(n_1327), .B1(n_1385), .B2(n_1450), .C1(n_1458), .C2(n_1460), .Y(n_1457) );
NAND2xp5_ASAP7_75t_L g1482 ( .A(n_1304), .B(n_1318), .Y(n_1482) );
OR2x2_ASAP7_75t_L g1304 ( .A(n_1305), .B(n_1306), .Y(n_1304) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1307), .Y(n_1325) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1307), .B(n_1324), .Y(n_1358) );
AND3x1_ASAP7_75t_L g1376 ( .A(n_1307), .B(n_1324), .C(n_1352), .Y(n_1376) );
OR2x2_ASAP7_75t_L g1415 ( .A(n_1307), .B(n_1318), .Y(n_1415) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_1307), .B(n_1318), .Y(n_1417) );
NOR2xp33_ASAP7_75t_L g1438 ( .A(n_1307), .B(n_1439), .Y(n_1438) );
NAND2xp5_ASAP7_75t_L g1472 ( .A(n_1307), .B(n_1352), .Y(n_1472) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1309), .Y(n_1307) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1312), .B(n_1314), .Y(n_1311) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1312), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_1312), .B(n_1350), .Y(n_1369) );
INVx2_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
A2O1A1Ixp33_ASAP7_75t_L g1381 ( .A1(n_1313), .A2(n_1361), .B(n_1382), .C(n_1383), .Y(n_1381) );
A2O1A1Ixp33_ASAP7_75t_L g1412 ( .A1(n_1313), .A2(n_1371), .B(n_1413), .C(n_1414), .Y(n_1412) );
NAND2xp5_ASAP7_75t_L g1426 ( .A(n_1313), .B(n_1427), .Y(n_1426) );
NAND2xp5_ASAP7_75t_L g1480 ( .A(n_1313), .B(n_1371), .Y(n_1480) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
OR2x2_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1322), .Y(n_1315) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1459 ( .A(n_1317), .B(n_1399), .Y(n_1459) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_1318), .B(n_1319), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1318), .B(n_1325), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1318), .B(n_1358), .Y(n_1390) );
OR2x2_ASAP7_75t_L g1391 ( .A(n_1318), .B(n_1324), .Y(n_1391) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_1318), .B(n_1324), .Y(n_1413) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1319), .B(n_1338), .Y(n_1348) );
INVx2_ASAP7_75t_L g1353 ( .A(n_1319), .Y(n_1353) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1319), .Y(n_1375) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_1319), .B(n_1328), .Y(n_1425) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_1319), .B(n_1471), .Y(n_1470) );
OR2x2_ASAP7_75t_L g1481 ( .A(n_1319), .B(n_1482), .Y(n_1481) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1320), .B(n_1321), .Y(n_1319) );
OAI221xp5_ASAP7_75t_L g1420 ( .A1(n_1322), .A2(n_1342), .B1(n_1421), .B2(n_1425), .C(n_1426), .Y(n_1420) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_1323), .B(n_1351), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1323), .B(n_1352), .Y(n_1424) );
AND2x2_ASAP7_75t_L g1323 ( .A(n_1324), .B(n_1325), .Y(n_1323) );
AOI321xp33_ASAP7_75t_L g1347 ( .A1(n_1324), .A2(n_1326), .A3(n_1348), .B1(n_1349), .B2(n_1350), .C(n_1354), .Y(n_1347) );
CKINVDCx14_ASAP7_75t_R g1326 ( .A(n_1327), .Y(n_1326) );
NAND2xp5_ASAP7_75t_L g1377 ( .A(n_1327), .B(n_1361), .Y(n_1377) );
INVx3_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1328), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1328), .B(n_1338), .Y(n_1371) );
OR2x2_ASAP7_75t_L g1383 ( .A(n_1328), .B(n_1337), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_1328), .B(n_1419), .Y(n_1418) );
OR2x2_ASAP7_75t_L g1436 ( .A(n_1328), .B(n_1338), .Y(n_1436) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_1328), .B(n_1337), .Y(n_1441) );
AND2x4_ASAP7_75t_L g1328 ( .A(n_1329), .B(n_1330), .Y(n_1328) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1333), .Y(n_1332) );
NOR2xp33_ASAP7_75t_SL g1333 ( .A(n_1334), .B(n_1337), .Y(n_1333) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_1335), .B(n_1353), .Y(n_1393) );
AND2x2_ASAP7_75t_L g1434 ( .A(n_1335), .B(n_1337), .Y(n_1434) );
NOR2xp33_ASAP7_75t_L g1343 ( .A(n_1337), .B(n_1344), .Y(n_1343) );
NAND3xp33_ASAP7_75t_L g1442 ( .A(n_1337), .B(n_1358), .C(n_1443), .Y(n_1442) );
NAND2xp5_ASAP7_75t_L g1474 ( .A(n_1337), .B(n_1429), .Y(n_1474) );
CKINVDCx6p67_ASAP7_75t_R g1337 ( .A(n_1338), .Y(n_1337) );
OR2x2_ASAP7_75t_L g1449 ( .A(n_1338), .B(n_1447), .Y(n_1449) );
NAND2xp5_ASAP7_75t_L g1462 ( .A(n_1338), .B(n_1362), .Y(n_1462) );
OR2x6_ASAP7_75t_L g1338 ( .A(n_1339), .B(n_1341), .Y(n_1338) );
OR2x2_ASAP7_75t_L g1359 ( .A(n_1339), .B(n_1341), .Y(n_1359) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
INVx2_ASAP7_75t_L g1469 ( .A(n_1344), .Y(n_1469) );
OAI332xp33_ASAP7_75t_L g1475 ( .A1(n_1344), .A2(n_1375), .A3(n_1436), .B1(n_1476), .B2(n_1478), .B3(n_1479), .C1(n_1480), .C2(n_1481), .Y(n_1475) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
CKINVDCx14_ASAP7_75t_R g1479 ( .A(n_1348), .Y(n_1479) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1351), .B(n_1358), .Y(n_1409) );
AND2x2_ASAP7_75t_L g1351 ( .A(n_1352), .B(n_1353), .Y(n_1351) );
AND2x2_ASAP7_75t_L g1455 ( .A(n_1352), .B(n_1399), .Y(n_1455) );
OR2x2_ASAP7_75t_L g1466 ( .A(n_1352), .B(n_1467), .Y(n_1466) );
NAND2xp5_ASAP7_75t_SL g1476 ( .A(n_1352), .B(n_1477), .Y(n_1476) );
NOR2xp33_ASAP7_75t_L g1414 ( .A(n_1353), .B(n_1415), .Y(n_1414) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
NAND3xp33_ASAP7_75t_L g1355 ( .A(n_1356), .B(n_1358), .C(n_1359), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1454 ( .A(n_1356), .B(n_1455), .Y(n_1454) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
OR2x2_ASAP7_75t_L g1477 ( .A(n_1358), .B(n_1399), .Y(n_1477) );
NOR2xp33_ASAP7_75t_L g1453 ( .A(n_1359), .B(n_1454), .Y(n_1453) );
AOI221xp5_ASAP7_75t_L g1378 ( .A1(n_1360), .A2(n_1379), .B1(n_1381), .B2(n_1384), .C(n_1388), .Y(n_1378) );
A2O1A1Ixp33_ASAP7_75t_L g1431 ( .A1(n_1360), .A2(n_1374), .B(n_1432), .C(n_1435), .Y(n_1431) );
AOI311xp33_ASAP7_75t_L g1445 ( .A1(n_1360), .A2(n_1446), .A3(n_1447), .B(n_1448), .C(n_1453), .Y(n_1445) );
INVx3_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
INVx2_ASAP7_75t_SL g1361 ( .A(n_1362), .Y(n_1361) );
INVx2_ASAP7_75t_SL g1429 ( .A(n_1362), .Y(n_1429) );
OAI22xp5_ASAP7_75t_SL g1363 ( .A1(n_1364), .A2(n_1365), .B1(n_1366), .B2(n_1367), .Y(n_1363) );
OAI221xp5_ASAP7_75t_L g1368 ( .A1(n_1369), .A2(n_1370), .B1(n_1372), .B2(n_1377), .C(n_1378), .Y(n_1368) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
AND2x2_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1376), .Y(n_1373) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1374), .Y(n_1404) );
NAND2xp5_ASAP7_75t_L g1428 ( .A(n_1374), .B(n_1424), .Y(n_1428) );
NOR2xp33_ASAP7_75t_L g1451 ( .A(n_1374), .B(n_1415), .Y(n_1451) );
INVx2_ASAP7_75t_L g1374 ( .A(n_1375), .Y(n_1374) );
AND2x2_ASAP7_75t_L g1446 ( .A(n_1375), .B(n_1390), .Y(n_1446) );
NAND2xp5_ASAP7_75t_SL g1460 ( .A(n_1375), .B(n_1386), .Y(n_1460) );
INVx2_ASAP7_75t_L g1387 ( .A(n_1376), .Y(n_1387) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
OAI211xp5_ASAP7_75t_L g1395 ( .A1(n_1383), .A2(n_1396), .B(n_1400), .C(n_1407), .Y(n_1395) );
NOR2xp33_ASAP7_75t_L g1384 ( .A(n_1385), .B(n_1387), .Y(n_1384) );
INVx2_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
AOI21xp33_ASAP7_75t_L g1388 ( .A1(n_1389), .A2(n_1391), .B(n_1392), .Y(n_1388) );
NAND2xp5_ASAP7_75t_L g1422 ( .A(n_1389), .B(n_1423), .Y(n_1422) );
OAI221xp5_ASAP7_75t_L g1435 ( .A1(n_1389), .A2(n_1436), .B1(n_1437), .B2(n_1440), .C(n_1442), .Y(n_1435) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
OAI21xp5_ASAP7_75t_SL g1394 ( .A1(n_1395), .A2(n_1420), .B(n_1429), .Y(n_1394) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
NAND2xp5_ASAP7_75t_L g1403 ( .A(n_1398), .B(n_1404), .Y(n_1403) );
NAND2xp5_ASAP7_75t_L g1433 ( .A(n_1399), .B(n_1434), .Y(n_1433) );
OAI21xp5_ASAP7_75t_L g1400 ( .A1(n_1401), .A2(n_1402), .B(n_1405), .Y(n_1400) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1403), .Y(n_1402) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
O2A1O1Ixp33_ASAP7_75t_L g1407 ( .A1(n_1408), .A2(n_1409), .B(n_1410), .C(n_1411), .Y(n_1407) );
NOR2xp33_ASAP7_75t_L g1464 ( .A(n_1408), .B(n_1465), .Y(n_1464) );
CKINVDCx6p67_ASAP7_75t_R g1447 ( .A(n_1410), .Y(n_1447) );
NAND2xp5_ASAP7_75t_L g1411 ( .A(n_1412), .B(n_1416), .Y(n_1411) );
NAND2xp5_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1418), .Y(n_1416) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1417), .Y(n_1478) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1422), .Y(n_1421) );
OAI22xp33_ASAP7_75t_L g1448 ( .A1(n_1423), .A2(n_1449), .B1(n_1450), .B2(n_1452), .Y(n_1448) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
NAND3xp33_ASAP7_75t_L g1430 ( .A(n_1431), .B(n_1445), .C(n_1456), .Y(n_1430) );
CKINVDCx5p33_ASAP7_75t_R g1432 ( .A(n_1433), .Y(n_1432) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1434), .Y(n_1452) );
INVxp67_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
AOI221xp5_ASAP7_75t_L g1456 ( .A1(n_1457), .A2(n_1461), .B1(n_1463), .B2(n_1473), .C(n_1475), .Y(n_1456) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1472), .Y(n_1471) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
CKINVDCx20_ASAP7_75t_R g1483 ( .A(n_1484), .Y(n_1483) );
CKINVDCx20_ASAP7_75t_R g1484 ( .A(n_1485), .Y(n_1484) );
INVx4_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
INVx1_ASAP7_75t_L g1488 ( .A(n_1489), .Y(n_1488) );
NAND2xp5_ASAP7_75t_L g1489 ( .A(n_1490), .B(n_1509), .Y(n_1489) );
NAND3xp33_ASAP7_75t_L g1491 ( .A(n_1492), .B(n_1495), .C(n_1498), .Y(n_1491) );
AOI22xp33_ASAP7_75t_L g1517 ( .A1(n_1496), .A2(n_1497), .B1(n_1518), .B2(n_1520), .Y(n_1517) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1515), .Y(n_1514) );
INVx2_ASAP7_75t_L g1518 ( .A(n_1519), .Y(n_1518) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
INVx4_ASAP7_75t_L g1524 ( .A(n_1525), .Y(n_1524) );
INVx2_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
INVxp67_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
BUFx3_ASAP7_75t_L g1536 ( .A(n_1537), .Y(n_1536) );
INVx1_ASAP7_75t_SL g1541 ( .A(n_1542), .Y(n_1541) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1543), .Y(n_1542) );
NAND3x1_ASAP7_75t_L g1544 ( .A(n_1545), .B(n_1571), .C(n_1581), .Y(n_1544) );
NAND3xp33_ASAP7_75t_L g1561 ( .A(n_1562), .B(n_1567), .C(n_1570), .Y(n_1561) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
HB1xp67_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
BUFx6f_ASAP7_75t_L g1583 ( .A(n_1584), .Y(n_1583) );
INVx1_ASAP7_75t_SL g1586 ( .A(n_1587), .Y(n_1586) );
INVx2_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1592), .Y(n_1591) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
INVx1_ASAP7_75t_L g1595 ( .A(n_1596), .Y(n_1595) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1599), .Y(n_1598) );
endmodule