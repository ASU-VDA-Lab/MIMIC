module fake_jpeg_16979_n_70 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_70);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_70;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

INVx2_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_21),
.B(n_23),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_10),
.A2(n_15),
.B1(n_18),
.B2(n_11),
.Y(n_22)
);

OAI32xp33_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_24),
.A3(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_0),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_15),
.A2(n_1),
.B1(n_9),
.B2(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_16),
.B(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_14),
.B(n_4),
.Y(n_39)
);

MAJx2_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_17),
.C(n_11),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_20),
.C(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_17),
.Y(n_35)
);

XNOR2x2_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_41),
.Y(n_48)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_33),
.A2(n_13),
.B1(n_27),
.B2(n_26),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_20),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_41),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_28),
.B(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_29),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_39),
.B1(n_38),
.B2(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_49),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_34),
.B(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_48),
.B1(n_49),
.B2(n_47),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_58),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_55),
.B(n_34),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_57),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_36),
.C(n_32),
.Y(n_58)
);

OAI21x1_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_51),
.B(n_50),
.Y(n_62)
);

AOI31xp67_ASAP7_75t_SL g66 ( 
.A1(n_62),
.A2(n_2),
.A3(n_5),
.B(n_9),
.Y(n_66)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_5),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_59),
.B1(n_52),
.B2(n_8),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_67),
.C(n_63),
.Y(n_68)
);

AOI211xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_61),
.B(n_25),
.C(n_34),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_69),
.Y(n_70)
);


endmodule