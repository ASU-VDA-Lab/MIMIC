module real_jpeg_18930_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_613, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_613;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_611;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_323;
wire n_215;
wire n_596;
wire n_312;
wire n_325;
wire n_316;
wire n_594;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_572;
wire n_586;
wire n_155;
wire n_405;
wire n_412;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_358;
wire n_181;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_597;
wire n_42;
wire n_268;
wire n_313;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_0),
.A2(n_21),
.B(n_610),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_0),
.B(n_611),
.Y(n_610)
);

INVxp33_ASAP7_75t_L g611 ( 
.A(n_1),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_2),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_2),
.Y(n_136)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_2),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g539 ( 
.A(n_2),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_3),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_3),
.Y(n_103)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_3),
.Y(n_151)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_3),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_4),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_4),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_4),
.A2(n_234),
.B1(n_256),
.B2(n_259),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_4),
.A2(n_234),
.B1(n_310),
.B2(n_316),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_4),
.A2(n_234),
.B1(n_388),
.B2(n_390),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_5),
.A2(n_83),
.B1(n_162),
.B2(n_165),
.Y(n_161)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_5),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_5),
.A2(n_165),
.B1(n_270),
.B2(n_274),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_5),
.A2(n_165),
.B1(n_446),
.B2(n_451),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_SL g505 ( 
.A1(n_5),
.A2(n_165),
.B1(n_506),
.B2(n_511),
.Y(n_505)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_6),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_6),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_6),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g493 ( 
.A(n_6),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_7),
.A2(n_184),
.B1(n_185),
.B2(n_188),
.Y(n_183)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_7),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_7),
.A2(n_188),
.B1(n_223),
.B2(n_378),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_7),
.A2(n_188),
.B1(n_601),
.B2(n_604),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_8),
.A2(n_116),
.B1(n_173),
.B2(n_176),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_8),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_8),
.A2(n_176),
.B1(n_331),
.B2(n_336),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_8),
.A2(n_176),
.B1(n_577),
.B2(n_580),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_9),
.A2(n_139),
.B1(n_140),
.B2(n_143),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_9),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_9),
.A2(n_139),
.B1(n_302),
.B2(n_305),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_9),
.A2(n_139),
.B1(n_440),
.B2(n_444),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_9),
.A2(n_139),
.B1(n_524),
.B2(n_528),
.Y(n_527)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_10),
.A2(n_33),
.B1(n_38),
.B2(n_39),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_10),
.A2(n_38),
.B1(n_249),
.B2(n_252),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_10),
.A2(n_38),
.B1(n_378),
.B2(n_407),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_10),
.A2(n_38),
.B1(n_457),
.B2(n_458),
.Y(n_456)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_11),
.Y(n_112)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_11),
.Y(n_119)
);

BUFx4f_ASAP7_75t_L g187 ( 
.A(n_11),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_11),
.Y(n_510)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_12),
.A2(n_115),
.B1(n_120),
.B2(n_121),
.Y(n_114)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_12),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_12),
.A2(n_120),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_12),
.A2(n_120),
.B1(n_350),
.B2(n_352),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g569 ( 
.A1(n_12),
.A2(n_120),
.B1(n_570),
.B2(n_572),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_13),
.A2(n_126),
.B1(n_131),
.B2(n_133),
.Y(n_125)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_13),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_13),
.A2(n_133),
.B1(n_205),
.B2(n_208),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_13),
.A2(n_133),
.B1(n_367),
.B2(n_370),
.Y(n_366)
);

OAI22xp33_ASAP7_75t_SL g594 ( 
.A1(n_13),
.A2(n_133),
.B1(n_595),
.B2(n_597),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_15),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_68)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_15),
.A2(n_74),
.B1(n_286),
.B2(n_289),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_15),
.A2(n_74),
.B1(n_143),
.B2(n_346),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_15),
.A2(n_74),
.B1(n_426),
.B2(n_428),
.Y(n_425)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_16),
.B(n_166),
.Y(n_319)
);

OAI32xp33_ASAP7_75t_L g414 ( 
.A1(n_16),
.A2(n_54),
.A3(n_90),
.B1(n_415),
.B2(n_418),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_16),
.B(n_78),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_SL g472 ( 
.A1(n_16),
.A2(n_82),
.B1(n_473),
.B2(n_474),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_16),
.A2(n_105),
.B1(n_527),
.B2(n_534),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_17),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_17),
.Y(n_227)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_17),
.Y(n_239)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_17),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_17),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_19),
.Y(n_101)
);

BUFx8_ASAP7_75t_L g164 ( 
.A(n_19),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g573 ( 
.A(n_19),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_586),
.Y(n_21)
);

OAI21xp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_557),
.B(n_585),
.Y(n_22)
);

INVxp67_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_396),
.B(n_552),
.Y(n_24)
);

NAND3xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_323),
.C(n_358),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_261),
.B(n_293),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_27),
.B(n_261),
.C(n_554),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_167),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_28),
.B(n_168),
.C(n_228),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_79),
.C(n_137),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_30),
.B(n_137),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_45),
.B1(n_68),
.B2(n_77),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_32),
.A2(n_78),
.B1(n_269),
.B2(n_281),
.Y(n_268)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_36),
.Y(n_307)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_37),
.Y(n_273)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_41),
.Y(n_580)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_43),
.Y(n_304)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_44),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_45),
.A2(n_68),
.B1(n_77),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_45),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_45),
.A2(n_77),
.B1(n_255),
.B2(n_349),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_45),
.A2(n_77),
.B1(n_301),
.B2(n_472),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_45),
.A2(n_77),
.B1(n_366),
.B2(n_576),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_45),
.A2(n_77),
.B1(n_576),
.B2(n_600),
.Y(n_599)
);

AO21x1_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_54),
.B(n_60),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22x1_ASAP7_75t_SL g153 ( 
.A1(n_52),
.A2(n_154),
.B1(n_157),
.B2(n_159),
.Y(n_153)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_61),
.B1(n_63),
.B2(n_65),
.Y(n_60)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_57),
.Y(n_369)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_58),
.Y(n_351)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_59),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_61),
.Y(n_233)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_61),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g335 ( 
.A(n_62),
.Y(n_335)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_62),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_64),
.Y(n_207)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_64),
.Y(n_417)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_73),
.Y(n_579)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_78),
.A2(n_269),
.B1(n_281),
.B2(n_300),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_78),
.A2(n_281),
.B1(n_364),
.B2(n_365),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_79),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_104),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_80),
.B(n_104),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_87),
.B1(n_93),
.B2(n_97),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_SL g283 ( 
.A1(n_81),
.A2(n_82),
.B(n_252),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_82),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_82),
.B(n_487),
.Y(n_486)
);

OAI21xp33_ASAP7_75t_SL g497 ( 
.A1(n_82),
.A2(n_486),
.B(n_498),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_82),
.B(n_134),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_R g540 ( 
.A(n_82),
.B(n_192),
.Y(n_540)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx6_ASAP7_75t_L g604 ( 
.A(n_90),
.Y(n_604)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_92),
.Y(n_158)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_92),
.Y(n_258)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_92),
.Y(n_374)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_92),
.Y(n_476)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OA21x2_ASAP7_75t_L g147 ( 
.A1(n_98),
.A2(n_148),
.B(n_153),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_100),
.Y(n_251)
);

INVx6_ASAP7_75t_L g389 ( 
.A(n_100),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_113),
.B1(n_125),
.B2(n_134),
.Y(n_104)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_105),
.A2(n_125),
.B1(n_172),
.B2(n_241),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_105),
.A2(n_183),
.B(n_340),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_105),
.A2(n_456),
.B1(n_459),
.B2(n_463),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_105),
.A2(n_505),
.B1(n_527),
.B2(n_537),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_111),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_106),
.A2(n_170),
.B1(n_309),
.B2(n_425),
.Y(n_424)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_109),
.Y(n_244)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_112),
.Y(n_524)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_114),
.A2(n_170),
.B1(n_309),
.B2(n_317),
.Y(n_308)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_115),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_118),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_119),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_131),
.Y(n_184)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_135),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_136),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_147),
.B1(n_160),
.B2(n_166),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_138),
.A2(n_147),
.B1(n_166),
.B2(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_146),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_146),
.Y(n_391)
);

INVx5_ASAP7_75t_L g571 ( 
.A(n_146),
.Y(n_571)
);

INVx3_ASAP7_75t_SL g247 ( 
.A(n_147),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_147),
.A2(n_166),
.B1(n_593),
.B2(n_594),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_158),
.Y(n_260)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_161),
.A2(n_247),
.B1(n_248),
.B2(n_253),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g252 ( 
.A(n_164),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_166),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_228),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_189),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_169),
.A2(n_190),
.B(n_212),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_177),
.B2(n_182),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_170),
.A2(n_504),
.B1(n_513),
.B2(n_515),
.Y(n_503)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_181),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_186),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_212),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_203),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_191),
.A2(n_213),
.B1(n_285),
.B2(n_292),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_191),
.A2(n_213),
.B1(n_376),
.B2(n_377),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_191),
.A2(n_213),
.B1(n_439),
.B2(n_445),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_191),
.A2(n_213),
.B1(n_406),
.B2(n_445),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_191),
.A2(n_213),
.B1(n_439),
.B2(n_497),
.Y(n_496)
);

OA21x2_ASAP7_75t_L g581 ( 
.A1(n_191),
.A2(n_213),
.B(n_377),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_192),
.A2(n_222),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_192),
.A2(n_204),
.B1(n_231),
.B2(n_330),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_192),
.A2(n_231),
.B1(n_405),
.B2(n_411),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_197),
.B1(n_198),
.B2(n_200),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_199),
.Y(n_427)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_221),
.Y(n_212)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_216),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_216),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_219),
.Y(n_485)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_245),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_229),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_240),
.Y(n_229)
);

XOR2x2_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_240),
.Y(n_265)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_232),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_239),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_239),
.Y(n_291)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_239),
.Y(n_422)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_239),
.Y(n_489)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_243),
.Y(n_242)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_254),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_246),
.B(n_254),
.C(n_326),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_247),
.A2(n_248),
.B1(n_253),
.B2(n_345),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_247),
.A2(n_253),
.B1(n_345),
.B2(n_387),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_247),
.A2(n_253),
.B1(n_387),
.B2(n_569),
.Y(n_568)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_252),
.Y(n_597)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.C(n_266),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_262),
.A2(n_263),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_265),
.B(n_267),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_282),
.C(n_284),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_284),
.Y(n_296)
);

INVx8_ASAP7_75t_L g473 ( 
.A(n_270),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_273),
.Y(n_355)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_296),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_285),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_288),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_320),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_294),
.B(n_320),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_297),
.C(n_298),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_295),
.B(n_399),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_297),
.B(n_298),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_308),
.C(n_319),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_299),
.B(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx3_ASAP7_75t_SL g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_308),
.B(n_319),
.Y(n_403)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_314),
.Y(n_457)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_315),
.Y(n_458)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_317),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx6_ASAP7_75t_L g514 ( 
.A(n_318),
.Y(n_514)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_321),
.Y(n_322)
);

A2O1A1O1Ixp25_ASAP7_75t_L g552 ( 
.A1(n_323),
.A2(n_358),
.B(n_553),
.C(n_555),
.D(n_556),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_357),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_SL g555 ( 
.A(n_324),
.B(n_357),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_327),
.Y(n_324)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_325),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_342),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_328),
.B(n_394),
.C(n_395),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_329),
.A2(n_338),
.B1(n_339),
.B2(n_341),
.Y(n_328)
);

INVxp33_ASAP7_75t_SL g341 ( 
.A(n_329),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_329),
.B(n_339),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_330),
.Y(n_376)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_334),
.Y(n_484)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_335),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_338),
.A2(n_339),
.B1(n_385),
.B2(n_386),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_338),
.A2(n_392),
.B1(n_564),
.B2(n_613),
.Y(n_563)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_342),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_356),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_348),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_344),
.B(n_348),
.C(n_356),
.Y(n_360)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_346),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_349),
.Y(n_364)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_359),
.B(n_393),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_359),
.B(n_393),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_360),
.B(n_560),
.C(n_561),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_381),
.Y(n_361)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_362),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_363),
.A2(n_375),
.B(n_380),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_375),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_380),
.A2(n_566),
.B1(n_583),
.B2(n_584),
.Y(n_565)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_380),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g560 ( 
.A(n_381),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_382),
.A2(n_383),
.B1(n_384),
.B2(n_392),
.Y(n_381)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_382),
.Y(n_392)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_385),
.Y(n_564)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx3_ASAP7_75t_SL g390 ( 
.A(n_391),
.Y(n_390)
);

AOI21x1_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_433),
.B(n_551),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_398),
.B(n_400),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_404),
.C(n_412),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g546 ( 
.A(n_402),
.B(n_547),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_404),
.A2(n_412),
.B1(n_413),
.B2(n_548),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_404),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_423),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_414),
.A2(n_423),
.B1(n_424),
.B2(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_414),
.Y(n_468)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_425),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

OAI21x1_ASAP7_75t_L g433 ( 
.A1(n_434),
.A2(n_545),
.B(n_550),
.Y(n_433)
);

AOI21x1_ASAP7_75t_L g434 ( 
.A1(n_435),
.A2(n_479),
.B(n_544),
.Y(n_434)
);

NAND2xp33_ASAP7_75t_SL g435 ( 
.A(n_436),
.B(n_466),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_436),
.B(n_466),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_455),
.C(n_464),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_437),
.A2(n_438),
.B1(n_464),
.B2(n_465),
.Y(n_500)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_453),
.Y(n_498)
);

INVx5_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_455),
.B(n_500),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_456),
.Y(n_515)
);

OAI32xp33_ASAP7_75t_L g482 ( 
.A1(n_458),
.A2(n_483),
.A3(n_485),
.B1(n_486),
.B2(n_490),
.Y(n_482)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_458),
.Y(n_494)
);

BUFx5_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_469),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_467),
.B(n_470),
.C(n_478),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_470),
.A2(n_471),
.B1(n_477),
.B2(n_478),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

OAI21x1_ASAP7_75t_L g479 ( 
.A1(n_480),
.A2(n_501),
.B(n_543),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_499),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_481),
.B(n_499),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_495),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_482),
.A2(n_495),
.B1(n_496),
.B2(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_482),
.Y(n_517)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx5_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_494),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_502),
.A2(n_518),
.B(n_542),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_516),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_503),
.B(n_516),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_510),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_512),
.Y(n_511)
);

INVx6_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_519),
.A2(n_535),
.B(n_541),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_526),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_525),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_522),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_536),
.B(n_540),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_536),
.B(n_540),
.Y(n_541)
);

INVx6_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

BUFx12f_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

NOR2xp67_ASAP7_75t_SL g545 ( 
.A(n_546),
.B(n_549),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_546),
.B(n_549),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_559),
.B(n_562),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_559),
.B(n_562),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_565),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_563),
.B(n_583),
.C(n_607),
.Y(n_606)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_566),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_566),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_567),
.A2(n_568),
.B1(n_574),
.B2(n_582),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_567),
.B(n_575),
.C(n_581),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_567),
.A2(n_568),
.B1(n_591),
.B2(n_605),
.Y(n_590)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_569),
.Y(n_593)
);

INVx6_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_574),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_575),
.B(n_581),
.Y(n_574)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

XNOR2x1_ASAP7_75t_L g598 ( 
.A(n_581),
.B(n_599),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_SL g586 ( 
.A(n_587),
.B(n_608),
.Y(n_586)
);

NOR2x1_ASAP7_75t_L g587 ( 
.A(n_588),
.B(n_606),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_588),
.B(n_606),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_589),
.B(n_590),
.Y(n_588)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_591),
.Y(n_605)
);

XNOR2x1_ASAP7_75t_L g591 ( 
.A(n_592),
.B(n_598),
.Y(n_591)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_602),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

INVxp33_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);


endmodule