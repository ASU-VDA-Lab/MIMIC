module fake_jpeg_13632_n_267 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_267);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_267;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_155;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_51),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_27),
.Y(n_47)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_SL g89 ( 
.A(n_49),
.Y(n_89)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_33),
.Y(n_98)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_8),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_25),
.Y(n_75)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_62),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_44),
.B1(n_46),
.B2(n_54),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_65),
.A2(n_35),
.B1(n_29),
.B2(n_31),
.Y(n_116)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g134 ( 
.A(n_66),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_69),
.B(n_80),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_36),
.B1(n_16),
.B2(n_23),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_72),
.A2(n_86),
.B1(n_20),
.B2(n_1),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_78),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_19),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_19),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_25),
.C(n_34),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_96),
.C(n_30),
.Y(n_105)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_50),
.A2(n_37),
.B1(n_29),
.B2(n_16),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_41),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_98),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_39),
.A2(n_34),
.B(n_31),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_26),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_101),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_63),
.B(n_30),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_88),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_104),
.B(n_121),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_105),
.B(n_106),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_68),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_65),
.A2(n_36),
.B1(n_35),
.B2(n_37),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_107),
.A2(n_116),
.B1(n_125),
.B2(n_129),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_79),
.A2(n_57),
.B1(n_21),
.B2(n_26),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_135),
.B1(n_128),
.B2(n_121),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_35),
.Y(n_121)
);

FAx1_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_41),
.CI(n_9),
.CON(n_122),
.SN(n_122)
);

OAI32xp33_ASAP7_75t_L g165 ( 
.A1(n_122),
.A2(n_7),
.A3(n_12),
.B1(n_5),
.B2(n_6),
.Y(n_165)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_74),
.A2(n_20),
.B1(n_8),
.B2(n_10),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_126),
.Y(n_148)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_64),
.A2(n_8),
.B1(n_14),
.B2(n_12),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_7),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_130),
.B(n_132),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_74),
.A2(n_20),
.B1(n_7),
.B2(n_10),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_131),
.A2(n_71),
.B1(n_81),
.B2(n_84),
.Y(n_154)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_68),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_70),
.B(n_0),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_137),
.Y(n_138)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_135),
.A2(n_103),
.B1(n_100),
.B2(n_85),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_139),
.A2(n_141),
.B1(n_144),
.B2(n_131),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_109),
.B(n_99),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_140),
.B(n_151),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_105),
.A2(n_103),
.B1(n_85),
.B2(n_91),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_142),
.A2(n_2),
.B1(n_134),
.B2(n_168),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_136),
.B1(n_123),
.B2(n_122),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_90),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_149),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_93),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_93),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_122),
.B(n_134),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_152),
.B(n_167),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_1),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_165),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_154),
.A2(n_156),
.B1(n_115),
.B2(n_124),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_107),
.A2(n_71),
.B1(n_84),
.B2(n_66),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_125),
.A2(n_97),
.B1(n_66),
.B2(n_20),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_157),
.A2(n_154),
.B(n_158),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_118),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_161),
.B(n_114),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_110),
.A2(n_97),
.B(n_2),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_162),
.A2(n_106),
.B(n_115),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_110),
.B(n_11),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_118),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_170),
.B(n_175),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_139),
.A2(n_152),
.B1(n_143),
.B2(n_141),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_173),
.B(n_193),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_172),
.B(n_190),
.Y(n_215)
);

BUFx24_ASAP7_75t_L g174 ( 
.A(n_163),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_174),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_132),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_138),
.B(n_127),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_180),
.C(n_183),
.Y(n_198)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_166),
.B(n_140),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_186),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_119),
.B1(n_133),
.B2(n_114),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_182),
.A2(n_194),
.B1(n_145),
.B2(n_157),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_161),
.B(n_14),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_168),
.B(n_1),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_192),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_188),
.A2(n_163),
.B1(n_148),
.B2(n_164),
.Y(n_204)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_2),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_2),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_145),
.A2(n_165),
.B1(n_162),
.B2(n_149),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_174),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_205),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_204),
.B1(n_212),
.B2(n_186),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_146),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_203),
.B(n_210),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_174),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_174),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_189),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_148),
.C(n_159),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_211),
.C(n_188),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_178),
.A2(n_164),
.B(n_159),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_178),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_155),
.C(n_169),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_155),
.B1(n_169),
.B2(n_194),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_220),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_219),
.C(n_221),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_218),
.A2(n_201),
.B1(n_223),
.B2(n_228),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_175),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_176),
.C(n_183),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_181),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_223),
.C(n_225),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_191),
.C(n_182),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_170),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_198),
.B(n_214),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_226),
.B(n_224),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_197),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_229),
.Y(n_233)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_231),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_238),
.Y(n_246)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_234),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_211),
.C(n_209),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_237),
.C(n_225),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_202),
.C(n_206),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_228),
.A2(n_196),
.B1(n_213),
.B2(n_204),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_230),
.A2(n_184),
.B(n_199),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_219),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_245),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_221),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_242),
.C(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_248),
.B(n_249),
.Y(n_256)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_R g250 ( 
.A(n_240),
.B(n_213),
.C(n_173),
.Y(n_250)
);

AOI21x1_ASAP7_75t_L g252 ( 
.A1(n_250),
.A2(n_246),
.B(n_193),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_254),
.C(n_218),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_252),
.A2(n_253),
.B(n_250),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_242),
.B(n_239),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_247),
.A2(n_213),
.B1(n_177),
.B2(n_227),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_256),
.A2(n_246),
.B1(n_205),
.B2(n_195),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_259),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_200),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_SL g263 ( 
.A1(n_258),
.A2(n_200),
.B(n_179),
.C(n_185),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_260),
.B(n_251),
.Y(n_262)
);

OAI21x1_ASAP7_75t_L g265 ( 
.A1(n_262),
.A2(n_263),
.B(n_202),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_190),
.B(n_192),
.Y(n_264)
);

NAND2xp33_ASAP7_75t_SL g266 ( 
.A(n_264),
.B(n_265),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_155),
.Y(n_267)
);


endmodule