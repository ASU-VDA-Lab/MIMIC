module real_jpeg_19770_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_206;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_0),
.A2(n_37),
.B1(n_38),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_0),
.A2(n_56),
.B1(n_60),
.B2(n_70),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_0),
.A2(n_56),
.B1(n_66),
.B2(n_67),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_0),
.A2(n_26),
.B1(n_28),
.B2(n_56),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_1),
.A2(n_66),
.B1(n_67),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_1),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_1),
.A2(n_26),
.B1(n_28),
.B2(n_87),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_1),
.A2(n_37),
.B1(n_38),
.B2(n_87),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_2),
.A2(n_26),
.B1(n_28),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_4),
.A2(n_60),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_4),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_4),
.A2(n_65),
.B(n_67),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_4),
.B(n_73),
.Y(n_116)
);

A2O1A1O1Ixp25_ASAP7_75t_L g128 ( 
.A1(n_4),
.A2(n_37),
.B(n_42),
.C(n_129),
.D(n_130),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_4),
.B(n_37),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_4),
.B(n_81),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_4),
.A2(n_24),
.B(n_144),
.Y(n_164)
);

A2O1A1O1Ixp25_ASAP7_75t_L g177 ( 
.A1(n_4),
.A2(n_66),
.B(n_78),
.C(n_96),
.D(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_4),
.B(n_66),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_5),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_5),
.A2(n_26),
.B1(n_28),
.B2(n_40),
.Y(n_119)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_7),
.B(n_145),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_9),
.A2(n_66),
.B1(n_67),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_9),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_9),
.A2(n_60),
.B1(n_70),
.B2(n_84),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_9),
.A2(n_37),
.B1(n_38),
.B2(n_84),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_9),
.A2(n_26),
.B1(n_28),
.B2(n_84),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_10),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_11),
.A2(n_37),
.B1(n_38),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_11),
.A2(n_26),
.B1(n_28),
.B2(n_48),
.Y(n_104)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_12),
.Y(n_79)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_15),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_122),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_120),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_20),
.B(n_105),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_88),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_50),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_35),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.B1(n_30),
.B2(n_33),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_24),
.A2(n_27),
.B1(n_32),
.B2(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_24),
.A2(n_25),
.B1(n_104),
.B2(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_24),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_24),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_24),
.B(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_25),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_25),
.A2(n_151),
.B(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_25),
.B(n_69),
.Y(n_166)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_26),
.A2(n_28),
.B1(n_43),
.B2(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_26),
.A2(n_44),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_28),
.B(n_43),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_28),
.B(n_166),
.Y(n_165)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_31),
.A2(n_162),
.B(n_186),
.Y(n_185)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_49),
.B(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_37),
.A2(n_38),
.B1(n_79),
.B2(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_37),
.A2(n_178),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_43),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_38),
.B(n_82),
.Y(n_183)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_41),
.A2(n_49),
.B1(n_141),
.B2(n_176),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_41),
.A2(n_176),
.B(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_54),
.Y(n_53)
);

CKINVDCx9p33_ASAP7_75t_R g46 ( 
.A(n_43),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_49),
.B(n_55),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_49),
.A2(n_53),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_49),
.B(n_69),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.C(n_75),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_51),
.A2(n_52),
.B1(n_75),
.B2(n_76),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_68),
.B(n_71),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B(n_63),
.C(n_64),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_62),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_60),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_60),
.A2(n_62),
.B(n_69),
.C(n_102),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_91),
.B(n_92),
.Y(n_90)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

O2A1O1Ixp33_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_79),
.B(n_80),
.C(n_81),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_79),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_77),
.A2(n_86),
.B(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_115),
.Y(n_114)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_80),
.Y(n_184)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_83),
.A2(n_85),
.B(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_99),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_93),
.B1(n_94),
.B2(n_98),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_90),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

AOI22x1_ASAP7_75t_SL g108 ( 
.A1(n_100),
.A2(n_101),
.B1(n_103),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_103),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.C(n_110),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_106),
.B(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_108),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.C(n_117),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_112),
.A2(n_113),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_116),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_201),
.B(n_206),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_189),
.B(n_200),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_170),
.B(n_188),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_147),
.B(n_169),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_135),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_127),
.B(n_135),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_128),
.A2(n_131),
.B1(n_132),
.B2(n_156),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_142),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_140),
.C(n_142),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_143),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_157),
.B(n_168),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_155),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_149),
.B(n_155),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_163),
.B(n_167),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_159),
.B(n_160),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_171),
.B(n_172),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_181),
.B2(n_187),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_175),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_177),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_180),
.C(n_187),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_181),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_185),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_190),
.B(n_191),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_196),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_197),
.C(n_198),
.Y(n_202)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_193),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_202),
.B(n_203),
.Y(n_206)
);


endmodule