module fake_jpeg_9525_n_23 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_23);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_23;

wire n_13;
wire n_21;
wire n_10;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

OAI21xp33_ASAP7_75t_L g7 ( 
.A1(n_3),
.A2(n_5),
.B(n_0),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_2),
.B(n_6),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_4),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_6),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_16),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_0),
.C(n_11),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_8),
.A2(n_7),
.B(n_9),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_18),
.B1(n_13),
.B2(n_14),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_7),
.A2(n_9),
.B(n_12),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_20),
.B(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_19),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_19),
.C(n_15),
.Y(n_23)
);


endmodule