module fake_ariane_2394_n_1090 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1090);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1090;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_423;
wire n_347;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_908;
wire n_850;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_952;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_349;
wire n_391;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_1016;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_515;
wire n_445;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_945;
wire n_702;
wire n_958;
wire n_905;
wire n_207;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_926;
wire n_813;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_1018;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_840;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_795;
wire n_1053;
wire n_1084;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_821;
wire n_928;
wire n_218;
wire n_839;
wire n_770;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_644;
wire n_536;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_206;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_638;
wire n_334;
wire n_887;
wire n_729;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_490;
wire n_262;
wire n_209;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_772;
wire n_741;
wire n_939;
wire n_847;
wire n_747;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_1081;
wire n_696;
wire n_1040;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_933;
wire n_872;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_492;
wire n_234;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_1026;
wire n_213;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_931;
wire n_827;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_999;
wire n_998;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_204;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_767;
wire n_736;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_149),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_84),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_136),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_164),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_29),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_167),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_19),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_49),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_95),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_177),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_18),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_109),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_38),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_91),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_110),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_17),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_4),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_66),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_113),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_114),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_63),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_68),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_67),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_0),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_97),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_39),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_53),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_4),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_191),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_111),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_9),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_152),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_86),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_59),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_76),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_137),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_105),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_140),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_124),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_121),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_188),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_123),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_194),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_96),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_98),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_157),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_184),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_93),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_134),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_169),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_170),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_183),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_23),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_117),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_13),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_21),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_162),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_100),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_130),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_71),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_193),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_11),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_17),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_79),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_203),
.Y(n_265)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_200),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_203),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_203),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_228),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_203),
.B(n_0),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_203),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_203),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_219),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_203),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_222),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_219),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_205),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_261),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_222),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_227),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_205),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_264),
.Y(n_285)
);

INVxp33_ASAP7_75t_SL g286 ( 
.A(n_207),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_225),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_212),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_227),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_221),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_226),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_236),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_263),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_210),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_197),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_210),
.Y(n_296)
);

INVxp33_ASAP7_75t_SL g297 ( 
.A(n_213),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_210),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_225),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_229),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_236),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_264),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_220),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_208),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_217),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_224),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_230),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_231),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_231),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_253),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_232),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_233),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_255),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_235),
.Y(n_314)
);

AND2x6_ASAP7_75t_L g315 ( 
.A(n_268),
.B(n_265),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_268),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_279),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_269),
.A2(n_262),
.B1(n_256),
.B2(n_202),
.Y(n_318)
);

AND2x4_ASAP7_75t_L g319 ( 
.A(n_279),
.B(n_238),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_269),
.A2(n_216),
.B1(n_240),
.B2(n_258),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_265),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_271),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_271),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_267),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_310),
.Y(n_326)
);

AND2x4_ASAP7_75t_L g327 ( 
.A(n_295),
.B(n_239),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_272),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_295),
.B(n_248),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_272),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_274),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_274),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_286),
.A2(n_249),
.B1(n_250),
.B2(n_257),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_270),
.Y(n_334)
);

CKINVDCx11_ASAP7_75t_R g335 ( 
.A(n_303),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_292),
.A2(n_260),
.B1(n_259),
.B2(n_252),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_276),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_310),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_266),
.B(n_196),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_276),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_273),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_277),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_313),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_294),
.B(n_296),
.Y(n_344)
);

NAND2xp33_ASAP7_75t_L g345 ( 
.A(n_273),
.B(n_198),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_298),
.B(n_199),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_277),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_280),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_280),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_282),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_282),
.Y(n_351)
);

AND2x6_ASAP7_75t_L g352 ( 
.A(n_284),
.B(n_34),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_311),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_304),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_305),
.B(n_201),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_313),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_306),
.B(n_307),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_284),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_285),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_281),
.Y(n_360)
);

AND2x4_ASAP7_75t_L g361 ( 
.A(n_312),
.B(n_204),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_281),
.Y(n_362)
);

XNOR2x1_ASAP7_75t_L g363 ( 
.A(n_283),
.B(n_1),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_314),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_285),
.Y(n_365)
);

CKINVDCx6p67_ASAP7_75t_R g366 ( 
.A(n_275),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_308),
.A2(n_251),
.B1(n_247),
.B2(n_246),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_287),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_287),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_335),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_354),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_366),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_366),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_354),
.Y(n_374)
);

BUFx10_ASAP7_75t_L g375 ( 
.A(n_341),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_326),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_341),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_326),
.Y(n_378)
);

NAND2x1_ASAP7_75t_L g379 ( 
.A(n_352),
.B(n_299),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_R g380 ( 
.A(n_338),
.B(n_278),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_338),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_356),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_317),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_356),
.Y(n_384)
);

BUFx10_ASAP7_75t_L g385 ( 
.A(n_361),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_364),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_364),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_343),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_358),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_359),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_339),
.B(n_278),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_339),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_359),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_316),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_367),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_367),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_369),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_336),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_360),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_362),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_320),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_320),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_369),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_333),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_317),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_358),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_R g407 ( 
.A(n_345),
.B(n_283),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_317),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_365),
.Y(n_409)
);

CKINVDCx6p67_ASAP7_75t_R g410 ( 
.A(n_361),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g411 ( 
.A(n_323),
.B(n_300),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_365),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_346),
.B(n_297),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_344),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_R g415 ( 
.A(n_334),
.B(n_289),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_318),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_358),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_355),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_368),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_355),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_361),
.B(n_309),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_368),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_368),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_351),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_351),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_351),
.Y(n_426)
);

NAND2xp33_ASAP7_75t_R g427 ( 
.A(n_361),
.B(n_289),
.Y(n_427)
);

INVxp33_ASAP7_75t_SL g428 ( 
.A(n_357),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_351),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_357),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_316),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_351),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_319),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_334),
.Y(n_434)
);

NAND2xp33_ASAP7_75t_SL g435 ( 
.A(n_327),
.B(n_301),
.Y(n_435)
);

NAND2xp33_ASAP7_75t_SL g436 ( 
.A(n_327),
.B(n_301),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_340),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_340),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_316),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_319),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_349),
.Y(n_441)
);

BUFx8_ASAP7_75t_L g442 ( 
.A(n_319),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_316),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_381),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_373),
.Y(n_445)
);

INVx5_ASAP7_75t_L g446 ( 
.A(n_385),
.Y(n_446)
);

OR2x6_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_319),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_377),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_411),
.B(n_327),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_383),
.Y(n_450)
);

OR2x6_ASAP7_75t_L g451 ( 
.A(n_392),
.B(n_327),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_389),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_371),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_372),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_415),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_414),
.B(n_334),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_383),
.Y(n_457)
);

AO22x2_ASAP7_75t_L g458 ( 
.A1(n_401),
.A2(n_363),
.B1(n_329),
.B2(n_302),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_437),
.B(n_321),
.Y(n_459)
);

OR2x6_ASAP7_75t_L g460 ( 
.A(n_392),
.B(n_329),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_374),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_406),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_386),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_423),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_424),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_387),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_370),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_413),
.B(n_334),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_329),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_438),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_413),
.B(n_334),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_441),
.Y(n_472)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_439),
.B(n_329),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_409),
.B(n_321),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_428),
.B(n_322),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_398),
.B(n_352),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_394),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_382),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_426),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_412),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_391),
.B(n_322),
.Y(n_481)
);

NAND2x1_ASAP7_75t_L g482 ( 
.A(n_425),
.B(n_315),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_390),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_393),
.B(n_324),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_380),
.B(n_363),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_376),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_430),
.B(n_288),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_380),
.B(n_323),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_375),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_404),
.B(n_324),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_397),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_403),
.B(n_328),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_425),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_432),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_394),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_434),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_385),
.B(n_325),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_417),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_378),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_433),
.B(n_290),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_384),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_419),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_415),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_388),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_440),
.B(n_407),
.Y(n_505)
);

BUFx10_ASAP7_75t_L g506 ( 
.A(n_399),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_400),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_375),
.B(n_323),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_416),
.B(n_325),
.Y(n_509)
);

AND2x2_ASAP7_75t_SL g510 ( 
.A(n_395),
.B(n_396),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_422),
.B(n_325),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g512 ( 
.A(n_418),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_442),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_442),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_410),
.B(n_325),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_420),
.B(n_353),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_394),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_443),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_429),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_394),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_431),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_405),
.B(n_353),
.Y(n_522)
);

OR2x6_ASAP7_75t_L g523 ( 
.A(n_427),
.B(n_353),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_427),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_408),
.B(n_325),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_431),
.B(n_328),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_431),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_469),
.B(n_349),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_469),
.B(n_291),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_451),
.B(n_293),
.Y(n_530)
);

AO22x2_ASAP7_75t_L g531 ( 
.A1(n_458),
.A2(n_402),
.B1(n_435),
.B2(n_436),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_448),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_468),
.B(n_407),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_492),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_453),
.Y(n_535)
);

NAND2x1p5_ASAP7_75t_L g536 ( 
.A(n_446),
.B(n_337),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_461),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_451),
.B(n_337),
.Y(n_538)
);

AO22x1_ASAP7_75t_L g539 ( 
.A1(n_485),
.A2(n_352),
.B1(n_350),
.B2(n_348),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_463),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_507),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_452),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_492),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_466),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_470),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_504),
.Y(n_546)
);

AO22x2_ASAP7_75t_L g547 ( 
.A1(n_458),
.A2(n_299),
.B1(n_302),
.B2(n_342),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_472),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_471),
.B(n_475),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_462),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_481),
.B(n_330),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_486),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_464),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_490),
.B(n_431),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_480),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_467),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_484),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_477),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_474),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_474),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_477),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_483),
.Y(n_562)
);

OR2x2_ASAP7_75t_SL g563 ( 
.A(n_499),
.B(n_342),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_459),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_491),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_501),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_459),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_504),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_509),
.B(n_330),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_518),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_484),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_451),
.B(n_347),
.Y(n_572)
);

BUFx8_ASAP7_75t_L g573 ( 
.A(n_514),
.Y(n_573)
);

NAND2x1p5_ASAP7_75t_L g574 ( 
.A(n_446),
.B(n_347),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_524),
.A2(n_315),
.B1(n_348),
.B2(n_350),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_494),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_512),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_526),
.Y(n_578)
);

NAND2x1p5_ASAP7_75t_L g579 ( 
.A(n_446),
.B(n_513),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_526),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_460),
.B(n_379),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_493),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_512),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_477),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_460),
.B(n_331),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_495),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_449),
.B(n_488),
.Y(n_587)
);

AO22x2_ASAP7_75t_L g588 ( 
.A1(n_496),
.A2(n_331),
.B1(n_332),
.B2(n_3),
.Y(n_588)
);

A2O1A1Ixp33_ASAP7_75t_L g589 ( 
.A1(n_511),
.A2(n_449),
.B(n_456),
.C(n_515),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_516),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_487),
.B(n_332),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_523),
.A2(n_315),
.B1(n_316),
.B2(n_352),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_450),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_503),
.A2(n_315),
.B1(n_234),
.B2(n_245),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_549),
.A2(n_525),
.B(n_522),
.Y(n_595)
);

OAI21xp33_ASAP7_75t_L g596 ( 
.A1(n_559),
.A2(n_444),
.B(n_498),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_551),
.A2(n_503),
.B(n_497),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_560),
.B(n_487),
.Y(n_598)
);

NOR2xp67_ASAP7_75t_L g599 ( 
.A(n_532),
.B(n_455),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_557),
.A2(n_457),
.B(n_450),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_564),
.B(n_510),
.Y(n_601)
);

A2O1A1Ixp33_ASAP7_75t_L g602 ( 
.A1(n_567),
.A2(n_502),
.B(n_476),
.C(n_508),
.Y(n_602)
);

O2A1O1Ixp33_ASAP7_75t_L g603 ( 
.A1(n_557),
.A2(n_460),
.B(n_505),
.C(n_500),
.Y(n_603)
);

NOR3xp33_ASAP7_75t_L g604 ( 
.A(n_541),
.B(n_489),
.C(n_479),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_577),
.B(n_500),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_L g606 ( 
.A1(n_571),
.A2(n_521),
.B(n_520),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_558),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_528),
.B(n_523),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_571),
.A2(n_457),
.B(n_482),
.Y(n_609)
);

O2A1O1Ixp33_ASAP7_75t_L g610 ( 
.A1(n_590),
.A2(n_523),
.B(n_447),
.C(n_454),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_554),
.A2(n_479),
.B(n_465),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_L g612 ( 
.A1(n_534),
.A2(n_527),
.B(n_473),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_533),
.A2(n_569),
.B(n_543),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_529),
.B(n_506),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_568),
.B(n_506),
.Y(n_615)
);

O2A1O1Ixp33_ASAP7_75t_L g616 ( 
.A1(n_552),
.A2(n_447),
.B(n_476),
.C(n_445),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_528),
.A2(n_543),
.B1(n_534),
.B2(n_537),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_565),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_529),
.B(n_465),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_589),
.A2(n_519),
.B(n_517),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_556),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_558),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_535),
.A2(n_519),
.B1(n_447),
.B2(n_495),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_546),
.B(n_478),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_593),
.A2(n_517),
.B(n_495),
.Y(n_625)
);

AOI33xp33_ASAP7_75t_L g626 ( 
.A1(n_540),
.A2(n_478),
.A3(n_2),
.B1(n_3),
.B2(n_5),
.B3(n_6),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_583),
.B(n_517),
.Y(n_627)
);

AOI21x1_ASAP7_75t_L g628 ( 
.A1(n_539),
.A2(n_473),
.B(n_352),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_558),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_587),
.B(n_473),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_593),
.A2(n_209),
.B(n_206),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_530),
.B(n_211),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_585),
.B(n_473),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_530),
.B(n_315),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_578),
.A2(n_580),
.B(n_591),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_578),
.A2(n_215),
.B(n_214),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_538),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_544),
.A2(n_218),
.B1(n_223),
.B2(n_237),
.Y(n_638)
);

NOR3xp33_ASAP7_75t_L g639 ( 
.A(n_566),
.B(n_242),
.C(n_241),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_545),
.A2(n_243),
.B1(n_244),
.B2(n_5),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_538),
.B(n_572),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_572),
.B(n_548),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_561),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_563),
.B(n_1),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_576),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_555),
.Y(n_646)
);

AO21x1_ASAP7_75t_L g647 ( 
.A1(n_580),
.A2(n_352),
.B(n_315),
.Y(n_647)
);

AO21x1_ASAP7_75t_L g648 ( 
.A1(n_562),
.A2(n_352),
.B(n_315),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_585),
.B(n_2),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_582),
.A2(n_36),
.B(n_35),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_581),
.A2(n_40),
.B(n_37),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_579),
.B(n_6),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_573),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_547),
.B(n_7),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_547),
.B(n_7),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_542),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g657 ( 
.A1(n_595),
.A2(n_594),
.B(n_575),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_598),
.B(n_531),
.Y(n_658)
);

A2O1A1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_603),
.A2(n_581),
.B(n_592),
.C(n_553),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_646),
.Y(n_660)
);

NOR3xp33_ASAP7_75t_SL g661 ( 
.A(n_621),
.B(n_596),
.C(n_640),
.Y(n_661)
);

NAND2x1p5_ASAP7_75t_L g662 ( 
.A(n_608),
.B(n_561),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_613),
.A2(n_584),
.B(n_561),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_645),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_620),
.A2(n_586),
.B(n_584),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_601),
.B(n_531),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_619),
.B(n_573),
.Y(n_667)
);

OAI21xp33_ASAP7_75t_L g668 ( 
.A1(n_626),
.A2(n_644),
.B(n_588),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_605),
.B(n_550),
.Y(n_669)
);

A2O1A1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_630),
.A2(n_616),
.B(n_602),
.C(n_617),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_599),
.A2(n_574),
.B1(n_536),
.B2(n_588),
.Y(n_671)
);

OAI21xp33_ASAP7_75t_L g672 ( 
.A1(n_654),
.A2(n_570),
.B(n_584),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_614),
.B(n_8),
.Y(n_673)
);

A2O1A1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_597),
.A2(n_586),
.B(n_9),
.C(n_10),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_611),
.A2(n_586),
.B(n_42),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_618),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_609),
.A2(n_600),
.B(n_612),
.Y(n_677)
);

INVx8_ASAP7_75t_L g678 ( 
.A(n_608),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_642),
.B(n_637),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_656),
.Y(n_680)
);

OAI21xp33_ASAP7_75t_L g681 ( 
.A1(n_655),
.A2(n_604),
.B(n_615),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_641),
.B(n_8),
.Y(n_682)
);

O2A1O1Ixp33_ASAP7_75t_L g683 ( 
.A1(n_632),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_683)
);

NOR3xp33_ASAP7_75t_SL g684 ( 
.A(n_624),
.B(n_12),
.C(n_13),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_607),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_627),
.B(n_14),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_649),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_623),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_688)
);

O2A1O1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_638),
.A2(n_15),
.B(n_16),
.C(n_18),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_607),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_633),
.B(n_19),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_635),
.Y(n_692)
);

AND2x6_ASAP7_75t_L g693 ( 
.A(n_633),
.B(n_41),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_606),
.A2(n_44),
.B(n_43),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_652),
.B(n_20),
.Y(n_695)
);

OAI21x1_ASAP7_75t_L g696 ( 
.A1(n_625),
.A2(n_46),
.B(n_45),
.Y(n_696)
);

NOR2xp67_ASAP7_75t_L g697 ( 
.A(n_634),
.B(n_47),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_607),
.Y(n_698)
);

INVx5_ASAP7_75t_L g699 ( 
.A(n_622),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_610),
.B(n_20),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_653),
.Y(n_701)
);

A2O1A1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_636),
.A2(n_21),
.B(n_22),
.C(n_23),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_622),
.Y(n_703)
);

OA22x2_ASAP7_75t_L g704 ( 
.A1(n_639),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_622),
.B(n_24),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_629),
.Y(n_706)
);

OAI21x1_ASAP7_75t_L g707 ( 
.A1(n_628),
.A2(n_128),
.B(n_195),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_629),
.B(n_25),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_SL g709 ( 
.A(n_629),
.B(n_48),
.Y(n_709)
);

CKINVDCx20_ASAP7_75t_R g710 ( 
.A(n_643),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_631),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_651),
.A2(n_129),
.B(n_192),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_643),
.B(n_26),
.Y(n_713)
);

NAND2xp33_ASAP7_75t_L g714 ( 
.A(n_643),
.B(n_27),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_650),
.B(n_50),
.Y(n_715)
);

INVx6_ASAP7_75t_SL g716 ( 
.A(n_715),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_692),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_701),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_668),
.A2(n_647),
.B1(n_648),
.B2(n_30),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_676),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_660),
.Y(n_721)
);

BUFx5_ASAP7_75t_L g722 ( 
.A(n_693),
.Y(n_722)
);

BUFx2_ASAP7_75t_SL g723 ( 
.A(n_710),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_666),
.B(n_28),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_664),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_673),
.B(n_29),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_715),
.Y(n_727)
);

BUFx6f_ASAP7_75t_SL g728 ( 
.A(n_693),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_678),
.Y(n_729)
);

BUFx4f_ASAP7_75t_SL g730 ( 
.A(n_706),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_679),
.B(n_30),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_678),
.Y(n_732)
);

BUFx6f_ASAP7_75t_SL g733 ( 
.A(n_693),
.Y(n_733)
);

INVx3_ASAP7_75t_SL g734 ( 
.A(n_699),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_695),
.B(n_31),
.Y(n_735)
);

BUFx2_ASAP7_75t_SL g736 ( 
.A(n_699),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_680),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_678),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_669),
.Y(n_739)
);

INVx4_ASAP7_75t_L g740 ( 
.A(n_699),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_684),
.B(n_31),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_687),
.Y(n_742)
);

INVx1_ASAP7_75t_SL g743 ( 
.A(n_667),
.Y(n_743)
);

BUFx12f_ASAP7_75t_L g744 ( 
.A(n_693),
.Y(n_744)
);

INVx1_ASAP7_75t_SL g745 ( 
.A(n_662),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_700),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_685),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_668),
.B(n_32),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_690),
.Y(n_749)
);

OR2x2_ASAP7_75t_L g750 ( 
.A(n_658),
.B(n_686),
.Y(n_750)
);

BUFx4_ASAP7_75t_SL g751 ( 
.A(n_661),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_698),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_703),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_682),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_696),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_691),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_704),
.B(n_32),
.Y(n_757)
);

INVx5_ASAP7_75t_SL g758 ( 
.A(n_709),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_707),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_665),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_657),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_713),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_714),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_681),
.B(n_33),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_671),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_681),
.Y(n_766)
);

BUFx12f_ASAP7_75t_L g767 ( 
.A(n_683),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_705),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_672),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_708),
.Y(n_770)
);

INVxp67_ASAP7_75t_SL g771 ( 
.A(n_663),
.Y(n_771)
);

CKINVDCx16_ASAP7_75t_R g772 ( 
.A(n_711),
.Y(n_772)
);

INVx8_ASAP7_75t_L g773 ( 
.A(n_659),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_674),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_670),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_675),
.Y(n_776)
);

CKINVDCx6p67_ASAP7_75t_R g777 ( 
.A(n_689),
.Y(n_777)
);

OR2x6_ASAP7_75t_L g778 ( 
.A(n_744),
.B(n_677),
.Y(n_778)
);

OAI221xp5_ASAP7_75t_L g779 ( 
.A1(n_748),
.A2(n_702),
.B1(n_688),
.B2(n_694),
.C(n_712),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_746),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_L g781 ( 
.A1(n_775),
.A2(n_697),
.B(n_33),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_727),
.B(n_697),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_766),
.A2(n_746),
.B(n_774),
.Y(n_783)
);

OAI21x1_ASAP7_75t_L g784 ( 
.A1(n_776),
.A2(n_51),
.B(n_52),
.Y(n_784)
);

AOI21x1_ASAP7_75t_L g785 ( 
.A1(n_759),
.A2(n_54),
.B(n_55),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_718),
.Y(n_786)
);

OAI21x1_ASAP7_75t_L g787 ( 
.A1(n_776),
.A2(n_56),
.B(n_57),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_743),
.B(n_58),
.Y(n_788)
);

OA21x2_ASAP7_75t_L g789 ( 
.A1(n_759),
.A2(n_60),
.B(n_61),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_750),
.B(n_62),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_718),
.Y(n_791)
);

AOI221xp5_ASAP7_75t_L g792 ( 
.A1(n_757),
.A2(n_64),
.B1(n_65),
.B2(n_69),
.C(n_70),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_721),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_725),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_772),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_795)
);

AO21x2_ASAP7_75t_L g796 ( 
.A1(n_755),
.A2(n_75),
.B(n_77),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_SL g797 ( 
.A1(n_731),
.A2(n_78),
.B(n_80),
.C(n_81),
.Y(n_797)
);

AOI22x1_ASAP7_75t_L g798 ( 
.A1(n_767),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_798)
);

O2A1O1Ixp33_ASAP7_75t_SL g799 ( 
.A1(n_754),
.A2(n_87),
.B(n_88),
.C(n_89),
.Y(n_799)
);

AO31x2_ASAP7_75t_L g800 ( 
.A1(n_755),
.A2(n_90),
.A3(n_92),
.B(n_94),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_719),
.A2(n_99),
.B(n_101),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_723),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_742),
.B(n_102),
.Y(n_803)
);

OAI21x1_ASAP7_75t_L g804 ( 
.A1(n_776),
.A2(n_103),
.B(n_104),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_739),
.B(n_106),
.Y(n_805)
);

AO31x2_ASAP7_75t_L g806 ( 
.A1(n_761),
.A2(n_107),
.A3(n_108),
.B(n_112),
.Y(n_806)
);

NAND2x1p5_ASAP7_75t_L g807 ( 
.A(n_763),
.B(n_115),
.Y(n_807)
);

CKINVDCx11_ASAP7_75t_R g808 ( 
.A(n_762),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_730),
.B(n_116),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_756),
.Y(n_810)
);

OAI21x1_ASAP7_75t_L g811 ( 
.A1(n_760),
.A2(n_118),
.B(n_119),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_737),
.Y(n_812)
);

NAND2x1p5_ASAP7_75t_L g813 ( 
.A(n_763),
.B(n_120),
.Y(n_813)
);

AOI21x1_ASAP7_75t_L g814 ( 
.A1(n_717),
.A2(n_122),
.B(n_125),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_719),
.A2(n_126),
.B(n_127),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_730),
.Y(n_816)
);

OA21x2_ASAP7_75t_L g817 ( 
.A1(n_771),
.A2(n_131),
.B(n_133),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_SL g818 ( 
.A1(n_728),
.A2(n_135),
.B(n_138),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_726),
.B(n_139),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_762),
.B(n_141),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_717),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_777),
.A2(n_763),
.B1(n_716),
.B2(n_764),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_720),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_752),
.Y(n_824)
);

CKINVDCx11_ASAP7_75t_R g825 ( 
.A(n_762),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_753),
.Y(n_826)
);

OAI21x1_ASAP7_75t_L g827 ( 
.A1(n_760),
.A2(n_142),
.B(n_143),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_777),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_769),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_765),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_727),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_762),
.B(n_147),
.Y(n_832)
);

OA21x2_ASAP7_75t_L g833 ( 
.A1(n_761),
.A2(n_148),
.B(n_150),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_808),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_786),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_780),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_794),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_831),
.B(n_793),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_812),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_829),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_821),
.Y(n_841)
);

CKINVDCx16_ASAP7_75t_R g842 ( 
.A(n_822),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_824),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_823),
.Y(n_844)
);

OAI21x1_ASAP7_75t_L g845 ( 
.A1(n_814),
.A2(n_760),
.B(n_727),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_826),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_830),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_783),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_801),
.A2(n_773),
.B1(n_767),
.B2(n_765),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_789),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_783),
.Y(n_851)
);

BUFx4_ASAP7_75t_SL g852 ( 
.A(n_791),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_801),
.A2(n_773),
.B1(n_728),
.B2(n_733),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_810),
.B(n_735),
.Y(n_854)
);

AOI21x1_ASAP7_75t_L g855 ( 
.A1(n_817),
.A2(n_724),
.B(n_741),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_778),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_778),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_778),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_822),
.B(n_773),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_800),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_789),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_825),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_802),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_800),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_800),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_806),
.Y(n_866)
);

INVx8_ASAP7_75t_L g867 ( 
.A(n_782),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_782),
.Y(n_868)
);

INVx6_ASAP7_75t_L g869 ( 
.A(n_832),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_807),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_815),
.A2(n_728),
.B1(n_733),
.B2(n_744),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_833),
.Y(n_872)
);

OAI21x1_ASAP7_75t_SL g873 ( 
.A1(n_781),
.A2(n_740),
.B(n_716),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_803),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_790),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_807),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_815),
.B(n_722),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_852),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_838),
.B(n_816),
.Y(n_879)
);

INVx8_ASAP7_75t_L g880 ( 
.A(n_867),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_835),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_840),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_849),
.A2(n_828),
.B1(n_781),
.B2(n_716),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_877),
.A2(n_779),
.B1(n_792),
.B2(n_733),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_836),
.B(n_838),
.Y(n_885)
);

NOR3xp33_ASAP7_75t_SL g886 ( 
.A(n_835),
.B(n_842),
.C(n_841),
.Y(n_886)
);

NAND2xp33_ASAP7_75t_R g887 ( 
.A(n_859),
.B(n_788),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_854),
.B(n_817),
.Y(n_888)
);

CKINVDCx16_ASAP7_75t_R g889 ( 
.A(n_834),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_877),
.A2(n_828),
.B1(n_798),
.B2(n_722),
.Y(n_890)
);

CKINVDCx16_ASAP7_75t_R g891 ( 
.A(n_834),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_862),
.Y(n_892)
);

CKINVDCx16_ASAP7_75t_R g893 ( 
.A(n_862),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_844),
.Y(n_894)
);

INVx4_ASAP7_75t_L g895 ( 
.A(n_870),
.Y(n_895)
);

O2A1O1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_874),
.A2(n_819),
.B(n_797),
.C(n_799),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_854),
.B(n_722),
.Y(n_897)
);

CKINVDCx16_ASAP7_75t_R g898 ( 
.A(n_842),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_837),
.Y(n_899)
);

NOR3xp33_ASAP7_75t_SL g900 ( 
.A(n_841),
.B(n_809),
.C(n_820),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_863),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_844),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_837),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_869),
.Y(n_904)
);

OAI21x1_ASAP7_75t_L g905 ( 
.A1(n_845),
.A2(n_785),
.B(n_787),
.Y(n_905)
);

NOR3xp33_ASAP7_75t_SL g906 ( 
.A(n_856),
.B(n_805),
.C(n_751),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_895),
.Y(n_907)
);

NOR2x1_ASAP7_75t_L g908 ( 
.A(n_888),
.B(n_859),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_888),
.B(n_856),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_898),
.B(n_857),
.Y(n_910)
);

NAND3xp33_ASAP7_75t_L g911 ( 
.A(n_900),
.B(n_848),
.C(n_851),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_879),
.B(n_857),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_899),
.Y(n_913)
);

OAI221xp5_ASAP7_75t_L g914 ( 
.A1(n_887),
.A2(n_853),
.B1(n_875),
.B2(n_871),
.C(n_855),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_882),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_895),
.B(n_897),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_904),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_899),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_903),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_903),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_878),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_879),
.B(n_858),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_883),
.A2(n_851),
.B1(n_848),
.B2(n_860),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_894),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_894),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_895),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_902),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_901),
.B(n_858),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_915),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_913),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_908),
.B(n_886),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_913),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_915),
.B(n_911),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_911),
.B(n_885),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_921),
.B(n_889),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_918),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_917),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_917),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_918),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_910),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_914),
.A2(n_896),
.B(n_890),
.C(n_906),
.Y(n_941)
);

O2A1O1Ixp5_ASAP7_75t_L g942 ( 
.A1(n_928),
.A2(n_897),
.B(n_855),
.C(n_839),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_908),
.B(n_904),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_929),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_934),
.B(n_923),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_931),
.B(n_916),
.Y(n_946)
);

NAND3xp33_ASAP7_75t_L g947 ( 
.A(n_933),
.B(n_941),
.C(n_942),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_940),
.A2(n_893),
.B1(n_891),
.B2(n_884),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_930),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_931),
.B(n_916),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_943),
.B(n_937),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_930),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_943),
.B(n_916),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_932),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_932),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_937),
.B(n_916),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_949),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_949),
.Y(n_958)
);

INVx1_ASAP7_75t_SL g959 ( 
.A(n_951),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_946),
.B(n_938),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_952),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_947),
.A2(n_938),
.B(n_940),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_946),
.B(n_928),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_956),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_959),
.B(n_944),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_960),
.B(n_951),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_964),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_964),
.B(n_945),
.Y(n_968)
);

OR2x6_ASAP7_75t_L g969 ( 
.A(n_962),
.B(n_935),
.Y(n_969)
);

NOR2x1p5_ASAP7_75t_L g970 ( 
.A(n_961),
.B(n_878),
.Y(n_970)
);

NAND3xp33_ASAP7_75t_L g971 ( 
.A(n_962),
.B(n_955),
.C(n_954),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_969),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_966),
.Y(n_973)
);

AOI221xp5_ASAP7_75t_L g974 ( 
.A1(n_968),
.A2(n_971),
.B1(n_957),
.B2(n_958),
.C(n_965),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_967),
.B(n_957),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_970),
.Y(n_976)
);

OAI21x1_ASAP7_75t_L g977 ( 
.A1(n_969),
.A2(n_958),
.B(n_956),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_966),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_965),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_965),
.B(n_963),
.Y(n_980)
);

OR2x2_ASAP7_75t_L g981 ( 
.A(n_965),
.B(n_953),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_966),
.B(n_950),
.Y(n_982)
);

XNOR2x1_ASAP7_75t_L g983 ( 
.A(n_979),
.B(n_948),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_973),
.B(n_978),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_982),
.B(n_953),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_980),
.B(n_936),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_972),
.A2(n_892),
.B1(n_936),
.B2(n_939),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_975),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_974),
.B(n_939),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_974),
.B(n_909),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_981),
.B(n_892),
.Y(n_991)
);

OAI32xp33_ASAP7_75t_L g992 ( 
.A1(n_990),
.A2(n_976),
.A3(n_975),
.B1(n_977),
.B2(n_907),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_985),
.B(n_881),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_984),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_986),
.B(n_919),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_989),
.A2(n_881),
.B(n_910),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_983),
.A2(n_919),
.B1(n_920),
.B2(n_922),
.Y(n_997)
);

OAI22xp33_ASAP7_75t_L g998 ( 
.A1(n_988),
.A2(n_870),
.B1(n_926),
.B2(n_907),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_991),
.B(n_912),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_987),
.A2(n_909),
.B1(n_870),
.B2(n_876),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_993),
.B(n_994),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_997),
.B(n_995),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_999),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_992),
.B(n_907),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_996),
.B(n_907),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_1000),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_998),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_993),
.B(n_912),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_1001),
.A2(n_818),
.B(n_920),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_1003),
.B(n_926),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_1002),
.Y(n_1011)
);

NAND2x1_ASAP7_75t_L g1012 ( 
.A(n_1004),
.B(n_926),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_1008),
.B(n_922),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1006),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1007),
.Y(n_1015)
);

OAI31xp33_ASAP7_75t_SL g1016 ( 
.A1(n_1005),
.A2(n_751),
.A3(n_905),
.B(n_758),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_1011),
.A2(n_926),
.B(n_813),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_1015),
.B(n_839),
.Y(n_1018)
);

NOR3xp33_ASAP7_75t_L g1019 ( 
.A(n_1014),
.B(n_827),
.C(n_811),
.Y(n_1019)
);

NOR2x1_ASAP7_75t_L g1020 ( 
.A(n_1012),
.B(n_736),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_SL g1021 ( 
.A1(n_1010),
.A2(n_813),
.B(n_833),
.Y(n_1021)
);

BUFx2_ASAP7_75t_R g1022 ( 
.A(n_1016),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_1013),
.A2(n_1009),
.B1(n_876),
.B2(n_758),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_1018),
.B(n_843),
.Y(n_1024)
);

OAI211xp5_ASAP7_75t_L g1025 ( 
.A1(n_1017),
.A2(n_795),
.B(n_880),
.C(n_740),
.Y(n_1025)
);

OAI321xp33_ASAP7_75t_L g1026 ( 
.A1(n_1023),
.A2(n_870),
.A3(n_846),
.B1(n_843),
.B2(n_770),
.C(n_768),
.Y(n_1026)
);

NAND4xp25_ASAP7_75t_L g1027 ( 
.A(n_1020),
.B(n_1022),
.C(n_1019),
.D(n_1021),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_1018),
.A2(n_880),
.B(n_873),
.Y(n_1028)
);

OAI21xp33_ASAP7_75t_L g1029 ( 
.A1(n_1027),
.A2(n_770),
.B(n_768),
.Y(n_1029)
);

AOI221xp5_ASAP7_75t_SL g1030 ( 
.A1(n_1028),
.A2(n_770),
.B1(n_768),
.B2(n_870),
.C(n_846),
.Y(n_1030)
);

NOR3x1_ASAP7_75t_L g1031 ( 
.A(n_1025),
.B(n_784),
.C(n_804),
.Y(n_1031)
);

NAND3xp33_ASAP7_75t_L g1032 ( 
.A(n_1024),
.B(n_740),
.C(n_770),
.Y(n_1032)
);

OAI22x1_ASAP7_75t_L g1033 ( 
.A1(n_1026),
.A2(n_734),
.B1(n_876),
.B2(n_868),
.Y(n_1033)
);

OAI211xp5_ASAP7_75t_SL g1034 ( 
.A1(n_1025),
.A2(n_868),
.B(n_758),
.C(n_927),
.Y(n_1034)
);

AOI222xp33_ASAP7_75t_L g1035 ( 
.A1(n_1026),
.A2(n_866),
.B1(n_864),
.B2(n_865),
.C1(n_860),
.C2(n_872),
.Y(n_1035)
);

AOI221xp5_ASAP7_75t_L g1036 ( 
.A1(n_1027),
.A2(n_768),
.B1(n_866),
.B2(n_924),
.C(n_925),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_1027),
.A2(n_880),
.B(n_873),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_1029),
.B(n_1034),
.Y(n_1038)
);

AOI221xp5_ASAP7_75t_L g1039 ( 
.A1(n_1036),
.A2(n_925),
.B1(n_924),
.B2(n_927),
.C(n_864),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1037),
.B(n_1030),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1032),
.Y(n_1041)
);

OAI21xp33_ASAP7_75t_SL g1042 ( 
.A1(n_1031),
.A2(n_905),
.B(n_845),
.Y(n_1042)
);

NOR2x1_ASAP7_75t_L g1043 ( 
.A(n_1033),
.B(n_796),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_1035),
.A2(n_734),
.B(n_796),
.C(n_729),
.Y(n_1044)
);

AOI222xp33_ASAP7_75t_L g1045 ( 
.A1(n_1036),
.A2(n_865),
.B1(n_925),
.B2(n_924),
.C1(n_872),
.C2(n_850),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_1037),
.B(n_880),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_1040),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1041),
.A2(n_869),
.B1(n_745),
.B2(n_729),
.Y(n_1048)
);

OR2x2_ASAP7_75t_L g1049 ( 
.A(n_1038),
.B(n_868),
.Y(n_1049)
);

NAND4xp25_ASAP7_75t_SL g1050 ( 
.A(n_1046),
.B(n_749),
.C(n_861),
.D(n_850),
.Y(n_1050)
);

NAND3xp33_ASAP7_75t_SL g1051 ( 
.A(n_1044),
.B(n_1039),
.C(n_1045),
.Y(n_1051)
);

OAI221xp5_ASAP7_75t_SL g1052 ( 
.A1(n_1042),
.A2(n_732),
.B1(n_861),
.B2(n_847),
.C(n_902),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1043),
.B(n_806),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_1041),
.A2(n_732),
.B(n_806),
.C(n_847),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1041),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_1038),
.A2(n_869),
.B1(n_867),
.B2(n_722),
.Y(n_1056)
);

NOR2xp67_ASAP7_75t_L g1057 ( 
.A(n_1040),
.B(n_151),
.Y(n_1057)
);

NOR3x1_ASAP7_75t_L g1058 ( 
.A(n_1041),
.B(n_153),
.C(n_154),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1041),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_R g1060 ( 
.A(n_1047),
.B(n_1059),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1055),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1057),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_1049),
.Y(n_1063)
);

INVxp67_ASAP7_75t_L g1064 ( 
.A(n_1051),
.Y(n_1064)
);

OA21x2_ASAP7_75t_L g1065 ( 
.A1(n_1053),
.A2(n_155),
.B(n_156),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_1048),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_1058),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1054),
.B(n_1056),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_1060),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1061),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_SL g1071 ( 
.A(n_1064),
.B(n_1052),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1063),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_SL g1073 ( 
.A1(n_1067),
.A2(n_1062),
.B1(n_1066),
.B2(n_1068),
.Y(n_1073)
);

CKINVDCx16_ASAP7_75t_R g1074 ( 
.A(n_1065),
.Y(n_1074)
);

AOI221x1_ASAP7_75t_L g1075 ( 
.A1(n_1072),
.A2(n_1065),
.B1(n_1050),
.B2(n_738),
.C(n_161),
.Y(n_1075)
);

OAI22x1_ASAP7_75t_SL g1076 ( 
.A1(n_1070),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_1069),
.A2(n_867),
.B(n_165),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1075),
.Y(n_1078)
);

OA22x2_ASAP7_75t_L g1079 ( 
.A1(n_1078),
.A2(n_1073),
.B1(n_1077),
.B2(n_1071),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1079),
.B(n_1074),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1080),
.A2(n_1076),
.B1(n_869),
.B2(n_738),
.Y(n_1081)
);

AOI221xp5_ASAP7_75t_SL g1082 ( 
.A1(n_1080),
.A2(n_163),
.B1(n_166),
.B2(n_168),
.C(n_171),
.Y(n_1082)
);

AOI222xp33_ASAP7_75t_L g1083 ( 
.A1(n_1082),
.A2(n_1081),
.B1(n_738),
.B2(n_174),
.C1(n_175),
.C2(n_176),
.Y(n_1083)
);

XOR2xp5_ASAP7_75t_L g1084 ( 
.A(n_1081),
.B(n_172),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_1083),
.A2(n_738),
.B1(n_722),
.B2(n_867),
.Y(n_1085)
);

AOI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1084),
.A2(n_722),
.B1(n_867),
.B2(n_179),
.Y(n_1086)
);

OA21x2_ASAP7_75t_L g1087 ( 
.A1(n_1085),
.A2(n_173),
.B(n_178),
.Y(n_1087)
);

OR2x6_ASAP7_75t_L g1088 ( 
.A(n_1086),
.B(n_747),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1087),
.A2(n_181),
.B(n_182),
.Y(n_1089)
);

AOI211xp5_ASAP7_75t_L g1090 ( 
.A1(n_1089),
.A2(n_1088),
.B(n_185),
.C(n_186),
.Y(n_1090)
);


endmodule