module fake_jpeg_24651_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_29),
.Y(n_50)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_26),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_50),
.B(n_0),
.Y(n_101)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_55),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_23),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_62),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_32),
.B1(n_26),
.B2(n_28),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_63),
.A2(n_26),
.B1(n_47),
.B2(n_28),
.Y(n_77)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_27),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_26),
.B1(n_32),
.B2(n_28),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_69),
.A2(n_83),
.B1(n_84),
.B2(n_100),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_55),
.B(n_37),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_73),
.B(n_85),
.Y(n_137)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_75),
.Y(n_110)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_77),
.A2(n_89),
.B1(n_93),
.B2(n_105),
.Y(n_112)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_80),
.Y(n_122)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_81),
.Y(n_121)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_44),
.B1(n_29),
.B2(n_45),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_32),
.B1(n_40),
.B2(n_23),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_53),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_87),
.Y(n_123)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

AO22x2_ASAP7_75t_L g91 ( 
.A1(n_63),
.A2(n_45),
.B1(n_38),
.B2(n_43),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_57),
.B1(n_40),
.B2(n_48),
.Y(n_111)
);

CKINVDCx12_ASAP7_75t_R g92 ( 
.A(n_52),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_20),
.Y(n_94)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_94),
.Y(n_135)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_51),
.A2(n_44),
.B1(n_45),
.B2(n_38),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_11),
.Y(n_133)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

CKINVDCx12_ASAP7_75t_R g106 ( 
.A(n_56),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_107),
.B(n_34),
.Y(n_127)
);

CKINVDCx12_ASAP7_75t_R g107 ( 
.A(n_64),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_50),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_116),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_51),
.B(n_62),
.Y(n_109)
);

AO21x1_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_97),
.B(n_20),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_118),
.B1(n_68),
.B2(n_60),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_65),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_60),
.B1(n_48),
.B2(n_38),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_70),
.B(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_43),
.Y(n_158)
);

O2A1O1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_88),
.A2(n_43),
.B(n_41),
.C(n_35),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_132),
.B1(n_16),
.B2(n_20),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_133),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_60),
.B1(n_48),
.B2(n_35),
.Y(n_132)
);

OAI22x1_ASAP7_75t_SL g138 ( 
.A1(n_119),
.A2(n_104),
.B1(n_83),
.B2(n_41),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_138),
.A2(n_133),
.B1(n_95),
.B2(n_21),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_139),
.A2(n_156),
.B(n_153),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_137),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_140),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_71),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_141),
.B(n_142),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_25),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_143),
.A2(n_156),
.B1(n_133),
.B2(n_123),
.Y(n_194)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_149),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_110),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_146),
.B(n_148),
.Y(n_184)
);

AO22x1_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_99),
.B1(n_43),
.B2(n_41),
.Y(n_147)
);

OA21x2_ASAP7_75t_L g189 ( 
.A1(n_147),
.A2(n_95),
.B(n_41),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_122),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_132),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_128),
.A2(n_78),
.B1(n_76),
.B2(n_93),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

AND2x6_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_104),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_158),
.C(n_126),
.Y(n_171)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_159),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_108),
.B(n_71),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_163),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_72),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_157),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_160),
.B(n_162),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_114),
.B(n_19),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_125),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_164),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_22),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_114),
.B(n_120),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_168),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_113),
.A2(n_43),
.B1(n_41),
.B2(n_16),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_167),
.A2(n_129),
.B1(n_130),
.B2(n_124),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_120),
.B(n_130),
.Y(n_168)
);

HAxp5_ASAP7_75t_SL g170 ( 
.A(n_138),
.B(n_126),
.CON(n_170),
.SN(n_170)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_170),
.A2(n_171),
.B(n_181),
.Y(n_212)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_176),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_179),
.A2(n_185),
.B1(n_194),
.B2(n_195),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_149),
.A2(n_129),
.B1(n_135),
.B2(n_115),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_180),
.A2(n_186),
.B1(n_139),
.B2(n_148),
.Y(n_217)
);

O2A1O1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_95),
.B(n_134),
.C(n_31),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_124),
.B1(n_136),
.B2(n_134),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_158),
.A2(n_27),
.B1(n_35),
.B2(n_16),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_189),
.A2(n_165),
.B1(n_145),
.B2(n_164),
.Y(n_213)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_191),
.Y(n_204)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_198),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_147),
.A2(n_27),
.B1(n_18),
.B2(n_25),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_197),
.B1(n_202),
.B2(n_142),
.Y(n_219)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_144),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_174),
.Y(n_218)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_201),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_139),
.A2(n_25),
.B1(n_18),
.B2(n_34),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_144),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_206),
.C(n_232),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_151),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_SL g235 ( 
.A(n_205),
.B(n_213),
.C(n_219),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_190),
.C(n_172),
.Y(n_206)
);

CKINVDCx12_ASAP7_75t_R g207 ( 
.A(n_169),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_217),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_187),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_209),
.Y(n_245)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_195),
.B(n_153),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_212),
.Y(n_236)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_222),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_192),
.B(n_162),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_221),
.B(n_228),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_140),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_183),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_224),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_184),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_193),
.A2(n_18),
.B(n_31),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_225),
.A2(n_196),
.B(n_24),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_200),
.A2(n_162),
.B1(n_160),
.B2(n_31),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_226),
.A2(n_181),
.B1(n_173),
.B2(n_182),
.Y(n_242)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_176),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_188),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_229),
.Y(n_255)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_177),
.B(n_160),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_173),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_30),
.C(n_24),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_249),
.Y(n_269)
);

NOR3xp33_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_177),
.C(n_180),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_237),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_244),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_175),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_241),
.C(n_250),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_187),
.C(n_188),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_182),
.B1(n_223),
.B2(n_232),
.Y(n_262)
);

NOR3xp33_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_202),
.C(n_189),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_205),
.A2(n_212),
.B1(n_214),
.B2(n_213),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_215),
.B1(n_217),
.B2(n_226),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_186),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_178),
.C(n_169),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_225),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_204),
.B(n_178),
.C(n_189),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_208),
.C(n_222),
.Y(n_264)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_228),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_256),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_235),
.A2(n_253),
.B1(n_205),
.B2(n_243),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_258),
.A2(n_260),
.B1(n_262),
.B2(n_277),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_235),
.A2(n_230),
.B1(n_218),
.B2(n_208),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_229),
.B(n_189),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_263),
.A2(n_0),
.B(n_1),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_270),
.C(n_272),
.Y(n_284)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_266),
.B(n_275),
.Y(n_294)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_271),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_227),
.C(n_220),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_227),
.C(n_211),
.Y(n_272)
);

INVxp33_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_211),
.C(n_30),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_252),
.C(n_251),
.Y(n_286)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

INVxp33_ASAP7_75t_SL g276 ( 
.A(n_245),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_255),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_248),
.A2(n_30),
.B1(n_19),
.B2(n_33),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_236),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_281),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_287),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_240),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g282 ( 
.A(n_264),
.B(n_249),
.CI(n_250),
.CON(n_282),
.SN(n_282)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_273),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_286),
.A2(n_288),
.B(n_277),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_268),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_246),
.C(n_233),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_258),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_291),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_257),
.B(n_242),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_260),
.B(n_238),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_263),
.C(n_265),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_8),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_280),
.A2(n_259),
.B1(n_272),
.B2(n_274),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_295),
.A2(n_297),
.B1(n_303),
.B2(n_308),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_296),
.A2(n_285),
.B(n_284),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_299),
.B(n_302),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_275),
.Y(n_302)
);

A2O1A1O1Ixp25_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_261),
.B(n_8),
.C(n_9),
.D(n_15),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_307),
.C(n_286),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_8),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_306),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_284),
.A2(n_7),
.B(n_15),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_294),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_290),
.A2(n_33),
.B1(n_1),
.B2(n_2),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_278),
.Y(n_309)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_309),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_289),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_318),
.Y(n_322)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_312),
.Y(n_320)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_314),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_288),
.C(n_282),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_315),
.A2(n_317),
.B(n_307),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_281),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_7),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_304),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_325),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_317),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_315),
.A2(n_297),
.B(n_312),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_318),
.Y(n_327)
);

AOI322xp5_ASAP7_75t_L g330 ( 
.A1(n_327),
.A2(n_323),
.A3(n_320),
.B1(n_319),
.B2(n_313),
.C1(n_309),
.C2(n_311),
.Y(n_330)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_322),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_328),
.A2(n_329),
.B1(n_9),
.B2(n_13),
.Y(n_331)
);

AO21x1_ASAP7_75t_L g332 ( 
.A1(n_330),
.A2(n_331),
.B(n_329),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_326),
.B(n_10),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_15),
.C(n_13),
.Y(n_334)
);

AOI322xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_10),
.A3(n_12),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_0),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_10),
.C(n_12),
.Y(n_336)
);

AOI321xp33_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_2),
.A3(n_3),
.B1(n_5),
.B2(n_300),
.C(n_237),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_2),
.Y(n_338)
);


endmodule