module fake_jpeg_25518_n_166 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_166);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_166;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx8_ASAP7_75t_SL g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_11),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_58),
.Y(n_65)
);

NAND2x1_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_67),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_0),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_70),
.B1(n_71),
.B2(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_1),
.Y(n_69)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_51),
.B(n_21),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_44),
.B(n_64),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_70),
.A2(n_52),
.B1(n_55),
.B2(n_46),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_45),
.Y(n_88)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_50),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_95),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_94),
.B1(n_102),
.B2(n_47),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_83),
.B1(n_79),
.B2(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_42),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_62),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_2),
.B(n_3),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_74),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_100),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_47),
.B1(n_59),
.B2(n_51),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_45),
.C(n_63),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_106),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_107),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_63),
.C(n_59),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_48),
.B1(n_47),
.B2(n_57),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_61),
.C(n_62),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_112),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_54),
.B(n_56),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_43),
.Y(n_119)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_117),
.B(n_98),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_94),
.B1(n_93),
.B2(n_86),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_122),
.B1(n_6),
.B2(n_7),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_48),
.B(n_3),
.Y(n_131)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_96),
.Y(n_126)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_121),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_109),
.A2(n_101),
.B1(n_89),
.B2(n_91),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_126),
.B(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_26),
.B(n_30),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_128),
.A2(n_131),
.B(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_92),
.Y(n_129)
);

FAx1_ASAP7_75t_SL g130 ( 
.A(n_116),
.B(n_54),
.CI(n_53),
.CON(n_130),
.SN(n_130)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_140),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_123),
.A2(n_20),
.B(n_41),
.Y(n_132)
);

OAI32xp33_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_2),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_136),
.B1(n_9),
.B2(n_10),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_4),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_135),
.B(n_138),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_25),
.C(n_40),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_11),
.B(n_12),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_124),
.B(n_8),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_139),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_141),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_147),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_149),
.C(n_137),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_140),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_142),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_155),
.Y(n_156)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_144),
.C(n_153),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_143),
.Y(n_158)
);

OAI221xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_146),
.B1(n_150),
.B2(n_145),
.C(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_134),
.B(n_19),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_18),
.C(n_24),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_27),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_164),
.Y(n_165)
);

FAx1_ASAP7_75t_SL g166 ( 
.A(n_165),
.B(n_130),
.CI(n_29),
.CON(n_166),
.SN(n_166)
);


endmodule