module fake_jpeg_18950_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx24_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_34),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_27),
.Y(n_53)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_33),
.A2(n_24),
.B1(n_17),
.B2(n_28),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_49),
.A2(n_34),
.B1(n_28),
.B2(n_29),
.Y(n_59)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_35),
.A2(n_23),
.B1(n_30),
.B2(n_16),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_51),
.B1(n_58),
.B2(n_24),
.Y(n_88)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NOR2x1_ASAP7_75t_R g92 ( 
.A(n_59),
.B(n_40),
.Y(n_92)
);

INVx5_ASAP7_75t_SL g61 ( 
.A(n_43),
.Y(n_61)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_30),
.B1(n_23),
.B2(n_36),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_88),
.B1(n_54),
.B2(n_50),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_65),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_32),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_32),
.Y(n_69)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_19),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_40),
.C(n_45),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_80),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_73),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_19),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_81),
.Y(n_100)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_43),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_18),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_19),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_19),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_94),
.Y(n_119)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_92),
.A2(n_67),
.B(n_57),
.Y(n_135)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_99),
.B(n_107),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_103),
.B(n_66),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_64),
.A2(n_72),
.B1(n_70),
.B2(n_73),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_106),
.A2(n_77),
.B1(n_23),
.B2(n_78),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_66),
.Y(n_107)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_22),
.C(n_18),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_106),
.C(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_111),
.B(n_117),
.Y(n_132)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_118),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_25),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_125),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_108),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_124),
.A2(n_135),
.B(n_138),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_76),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_128),
.Y(n_155)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_22),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_134),
.Y(n_159)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_96),
.A2(n_89),
.B1(n_91),
.B2(n_79),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_136),
.A2(n_27),
.B1(n_26),
.B2(n_18),
.Y(n_167)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_95),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_74),
.B(n_61),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_18),
.B(n_27),
.Y(n_170)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_102),
.A2(n_25),
.B(n_29),
.C(n_80),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_146),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_101),
.B1(n_113),
.B2(n_112),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_86),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_144),
.B(n_116),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_98),
.B(n_86),
.C(n_82),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_101),
.C(n_116),
.Y(n_150)
);

AO22x1_ASAP7_75t_L g146 ( 
.A1(n_98),
.A2(n_45),
.B1(n_68),
.B2(n_22),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_148),
.A2(n_165),
.B1(n_155),
.B2(n_179),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_153),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_22),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_166),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_157),
.B(n_162),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_128),
.B1(n_142),
.B2(n_124),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_158),
.A2(n_139),
.B1(n_145),
.B2(n_146),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_127),
.Y(n_162)
);

XOR2x1_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_22),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_174),
.B(n_179),
.Y(n_183)
);

OR2x6_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_18),
.Y(n_165)
);

AO22x1_ASAP7_75t_SL g182 ( 
.A1(n_165),
.A2(n_146),
.B1(n_135),
.B2(n_141),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_113),
.C(n_105),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_120),
.B1(n_138),
.B2(n_140),
.Y(n_194)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_122),
.B(n_27),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_178),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_170),
.A2(n_173),
.B(n_0),
.Y(n_209)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_136),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_119),
.A2(n_115),
.B(n_1),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_121),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_126),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_27),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_119),
.A2(n_27),
.B(n_115),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_185),
.Y(n_217)
);

OA21x2_ASAP7_75t_L g184 ( 
.A1(n_165),
.A2(n_135),
.B(n_120),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_184),
.A2(n_197),
.B(n_209),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_164),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_149),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_190),
.B(n_196),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_192),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_132),
.Y(n_193)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_194),
.A2(n_151),
.B1(n_173),
.B2(n_147),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_154),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_151),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_205),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_158),
.B1(n_161),
.B2(n_148),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_202),
.A2(n_203),
.B1(n_207),
.B2(n_211),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_140),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_204),
.B(n_206),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_152),
.B(n_31),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_161),
.B(n_10),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_152),
.B(n_31),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_212),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_21),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_210),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_165),
.A2(n_174),
.B1(n_170),
.B2(n_163),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_31),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_198),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_226),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_180),
.B(n_153),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_220),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_216),
.A2(n_202),
.B1(n_184),
.B2(n_182),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_180),
.B(n_156),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_173),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_223),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_167),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_183),
.B(n_203),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_229),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_187),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_147),
.B(n_10),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_227),
.A2(n_206),
.B1(n_195),
.B2(n_189),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_10),
.Y(n_228)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_200),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_21),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_233),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_21),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_208),
.C(n_205),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_244),
.C(n_245),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_224),
.Y(n_239)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_242),
.A2(n_248),
.B1(n_257),
.B2(n_218),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_186),
.C(n_184),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_209),
.C(n_212),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_237),
.A2(n_194),
.B1(n_188),
.B2(n_195),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_223),
.B1(n_229),
.B2(n_237),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_216),
.A2(n_182),
.B1(n_185),
.B2(n_188),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_236),
.Y(n_249)
);

AOI21xp33_ASAP7_75t_L g259 ( 
.A1(n_249),
.A2(n_221),
.B(n_227),
.Y(n_259)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_215),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_256),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_255),
.B(n_8),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_231),
.A2(n_199),
.B(n_191),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_225),
.A2(n_189),
.B1(n_191),
.B2(n_11),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_219),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_238),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_259),
.A2(n_0),
.B(n_1),
.Y(n_288)
);

INVxp33_ASAP7_75t_SL g260 ( 
.A(n_253),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_260),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_274),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_231),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_269),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_265),
.A2(n_14),
.B1(n_11),
.B2(n_8),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_240),
.A2(n_218),
.B1(n_235),
.B2(n_222),
.Y(n_266)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_248),
.B1(n_232),
.B2(n_257),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_276),
.B1(n_245),
.B2(n_247),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_268),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_26),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_20),
.C(n_26),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_0),
.C(n_2),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_7),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_269),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g276 ( 
.A(n_254),
.B(n_7),
.CI(n_13),
.CON(n_276),
.SN(n_276)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_284),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_281),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_254),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_262),
.A2(n_247),
.B1(n_14),
.B2(n_12),
.Y(n_283)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_288),
.B1(n_276),
.B2(n_4),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_272),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_5),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_273),
.Y(n_296)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_281),
.B(n_263),
.CI(n_275),
.CON(n_293),
.SN(n_293)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_264),
.C(n_271),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_299),
.C(n_278),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_302),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_297),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_3),
.C(n_4),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_3),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_300),
.A2(n_284),
.B(n_290),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_287),
.A2(n_5),
.B(n_3),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_291),
.Y(n_308)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_289),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_292),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_308),
.B(n_309),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_286),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_312),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_289),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_294),
.C(n_307),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_314),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_293),
.Y(n_320)
);

AOI31xp33_ASAP7_75t_L g318 ( 
.A1(n_304),
.A2(n_301),
.A3(n_298),
.B(n_293),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_305),
.B(n_311),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_319),
.B(n_320),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_321),
.B(n_315),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_313),
.C(n_317),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_316),
.B(n_299),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_4),
.C(n_5),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_326),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_4),
.Y(n_328)
);


endmodule